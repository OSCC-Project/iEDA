module gcd (
clk,
req_rdy,
req_val,
reset,
resp_rdy,
resp_val,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
req_msg,
resp_msg,
resp_msg,
resp_msg,
resp_msg,
resp_msg,
resp_msg,
resp_msg,
resp_msg,
resp_msg,
resp_msg,
resp_msg,
resp_msg,
resp_msg,
resp_msg,
resp_msg,
resp_msg
);

input clk ;
output req_rdy ;
input req_val ;
input reset ;
input resp_rdy ;
output resp_val ;
input [31:0] req_msg[0] ;
input [31:0] req_msg[1] ;
input [31:0] req_msg[2] ;
input [31:0] req_msg[3] ;
input [31:0] req_msg[4] ;
input [31:0] req_msg[5] ;
input [31:0] req_msg[6] ;
input [31:0] req_msg[7] ;
input [31:0] req_msg[8] ;
input [31:0] req_msg[9] ;
input [31:0] req_msg[10] ;
input [31:0] req_msg[11] ;
input [31:0] req_msg[12] ;
input [31:0] req_msg[13] ;
input [31:0] req_msg[14] ;
input [31:0] req_msg[15] ;
input [31:0] req_msg[16] ;
input [31:0] req_msg[17] ;
input [31:0] req_msg[18] ;
input [31:0] req_msg[19] ;
input [31:0] req_msg[20] ;
input [31:0] req_msg[21] ;
input [31:0] req_msg[22] ;
input [31:0] req_msg[23] ;
input [31:0] req_msg[24] ;
input [31:0] req_msg[25] ;
input [31:0] req_msg[26] ;
input [31:0] req_msg[27] ;
input [31:0] req_msg[28] ;
input [31:0] req_msg[29] ;
input [31:0] req_msg[30] ;
input [31:0] req_msg[31] ;
output [15:0] resp_msg[0] ;
output [15:0] resp_msg[1] ;
output [15:0] resp_msg[2] ;
output [15:0] resp_msg[3] ;
output [15:0] resp_msg[4] ;
output [15:0] resp_msg[5] ;
output [15:0] resp_msg[6] ;
output [15:0] resp_msg[7] ;
output [15:0] resp_msg[8] ;
output [15:0] resp_msg[9] ;
output [15:0] resp_msg[10] ;
output [15:0] resp_msg[11] ;
output [15:0] resp_msg[12] ;
output [15:0] resp_msg[13] ;
output [15:0] resp_msg[14] ;
output [15:0] resp_msg[15] ;

wire ctrl$a_reg_en ;
wire ctrl$b_mux_sel ;
wire ctrl$b_reg_en ;
wire ctrl$is_a_lt_b ;
wire ctrl$is_b_zero ;
wire \ctrl/_00_ ;
wire \ctrl/_01_ ;
wire \ctrl/_02_ ;
wire \ctrl/_03_ ;
wire \ctrl/_04_ ;
wire \ctrl/_05_ ;
wire \ctrl/_06_ ;
wire \ctrl/_07_ ;
wire \ctrl/_08_ ;
wire \ctrl/_09_ ;
wire \ctrl/_10_ ;
wire \ctrl/_11_ ;
wire \ctrl/_12_ ;
wire \ctrl/_13_ ;
wire \ctrl/_14_ ;
wire \ctrl/_15_ ;
wire \ctrl/_16_ ;
wire \ctrl/state/_00_ ;
wire \ctrl/state/_01_ ;
wire \ctrl/state/_02_ ;
wire \ctrl/state/_03_ ;
wire \ctrl/state/_04_ ;
wire \ctrl/state/_05_ ;
wire \ctrl/state/_06_ ;
wire \dpath/a_lt_b/_000_ ;
wire \dpath/a_lt_b/_001_ ;
wire \dpath/a_lt_b/_002_ ;
wire \dpath/a_lt_b/_003_ ;
wire \dpath/a_lt_b/_004_ ;
wire \dpath/a_lt_b/_005_ ;
wire \dpath/a_lt_b/_006_ ;
wire \dpath/a_lt_b/_007_ ;
wire \dpath/a_lt_b/_008_ ;
wire \dpath/a_lt_b/_009_ ;
wire \dpath/a_lt_b/_010_ ;
wire \dpath/a_lt_b/_011_ ;
wire \dpath/a_lt_b/_012_ ;
wire \dpath/a_lt_b/_013_ ;
wire \dpath/a_lt_b/_014_ ;
wire \dpath/a_lt_b/_015_ ;
wire \dpath/a_lt_b/_016_ ;
wire \dpath/a_lt_b/_017_ ;
wire \dpath/a_lt_b/_018_ ;
wire \dpath/a_lt_b/_019_ ;
wire \dpath/a_lt_b/_020_ ;
wire \dpath/a_lt_b/_021_ ;
wire \dpath/a_lt_b/_022_ ;
wire \dpath/a_lt_b/_023_ ;
wire \dpath/a_lt_b/_024_ ;
wire \dpath/a_lt_b/_025_ ;
wire \dpath/a_lt_b/_026_ ;
wire \dpath/a_lt_b/_027_ ;
wire \dpath/a_lt_b/_028_ ;
wire \dpath/a_lt_b/_029_ ;
wire \dpath/a_lt_b/_030_ ;
wire \dpath/a_lt_b/_031_ ;
wire \dpath/a_lt_b/_032_ ;
wire \dpath/a_lt_b/_033_ ;
wire \dpath/a_lt_b/_034_ ;
wire \dpath/a_lt_b/_035_ ;
wire \dpath/a_lt_b/_036_ ;
wire \dpath/a_lt_b/_037_ ;
wire \dpath/a_lt_b/_038_ ;
wire \dpath/a_lt_b/_039_ ;
wire \dpath/a_lt_b/_040_ ;
wire \dpath/a_lt_b/_041_ ;
wire \dpath/a_lt_b/_042_ ;
wire \dpath/a_lt_b/_043_ ;
wire \dpath/a_lt_b/_044_ ;
wire \dpath/a_lt_b/_045_ ;
wire \dpath/a_lt_b/_046_ ;
wire \dpath/a_lt_b/_047_ ;
wire \dpath/a_lt_b/_048_ ;
wire \dpath/a_lt_b/_049_ ;
wire \dpath/a_lt_b/_050_ ;
wire \dpath/a_lt_b/_051_ ;
wire \dpath/a_lt_b/_052_ ;
wire \dpath/a_lt_b/_053_ ;
wire \dpath/a_lt_b/_054_ ;
wire \dpath/a_lt_b/_055_ ;
wire \dpath/a_lt_b/_056_ ;
wire \dpath/a_lt_b/_057_ ;
wire \dpath/a_lt_b/_058_ ;
wire \dpath/a_lt_b/_059_ ;
wire \dpath/a_lt_b/_060_ ;
wire \dpath/a_lt_b/_061_ ;
wire \dpath/a_lt_b/_062_ ;
wire \dpath/a_lt_b/_063_ ;
wire \dpath/a_lt_b/_064_ ;
wire \dpath/a_lt_b/_065_ ;
wire \dpath/a_lt_b/_066_ ;
wire \dpath/a_lt_b/_067_ ;
wire \dpath/a_lt_b/_068_ ;
wire \dpath/a_lt_b/_069_ ;
wire \dpath/a_lt_b/_070_ ;
wire \dpath/a_lt_b/_071_ ;
wire \dpath/a_lt_b/_072_ ;
wire \dpath/a_lt_b/_073_ ;
wire \dpath/a_lt_b/_074_ ;
wire \dpath/a_lt_b/_075_ ;
wire \dpath/a_lt_b/_076_ ;
wire \dpath/a_lt_b/_077_ ;
wire \dpath/a_lt_b/_078_ ;
wire \dpath/a_lt_b/_079_ ;
wire \dpath/a_lt_b/_080_ ;
wire \dpath/a_lt_b/_081_ ;
wire \dpath/a_lt_b/_082_ ;
wire \dpath/a_lt_b/_083_ ;
wire \dpath/a_lt_b/_084_ ;
wire \dpath/a_lt_b/_085_ ;
wire \dpath/a_lt_b/_086_ ;
wire \dpath/a_lt_b/_087_ ;
wire \dpath/a_lt_b/_088_ ;
wire \dpath/a_lt_b/_089_ ;
wire \dpath/a_mux/_000_ ;
wire \dpath/a_mux/_001_ ;
wire \dpath/a_mux/_002_ ;
wire \dpath/a_mux/_003_ ;
wire \dpath/a_mux/_004_ ;
wire \dpath/a_mux/_005_ ;
wire \dpath/a_mux/_006_ ;
wire \dpath/a_mux/_007_ ;
wire \dpath/a_mux/_008_ ;
wire \dpath/a_mux/_009_ ;
wire \dpath/a_mux/_010_ ;
wire \dpath/a_mux/_011_ ;
wire \dpath/a_mux/_012_ ;
wire \dpath/a_mux/_013_ ;
wire \dpath/a_mux/_014_ ;
wire \dpath/a_mux/_015_ ;
wire \dpath/a_mux/_016_ ;
wire \dpath/a_mux/_017_ ;
wire \dpath/a_mux/_018_ ;
wire \dpath/a_mux/_019_ ;
wire \dpath/a_mux/_020_ ;
wire \dpath/a_mux/_021_ ;
wire \dpath/a_mux/_022_ ;
wire \dpath/a_mux/_023_ ;
wire \dpath/a_mux/_024_ ;
wire \dpath/a_mux/_025_ ;
wire \dpath/a_mux/_026_ ;
wire \dpath/a_mux/_027_ ;
wire \dpath/a_mux/_028_ ;
wire \dpath/a_mux/_029_ ;
wire \dpath/a_mux/_030_ ;
wire \dpath/a_mux/_031_ ;
wire \dpath/a_mux/_032_ ;
wire \dpath/a_mux/_033_ ;
wire \dpath/a_mux/_034_ ;
wire \dpath/a_mux/_035_ ;
wire \dpath/a_mux/_036_ ;
wire \dpath/a_mux/_037_ ;
wire \dpath/a_mux/_038_ ;
wire \dpath/a_mux/_039_ ;
wire \dpath/a_mux/_040_ ;
wire \dpath/a_mux/_041_ ;
wire \dpath/a_mux/_042_ ;
wire \dpath/a_mux/_043_ ;
wire \dpath/a_mux/_044_ ;
wire \dpath/a_mux/_045_ ;
wire \dpath/a_mux/_046_ ;
wire \dpath/a_mux/_047_ ;
wire \dpath/a_mux/_048_ ;
wire \dpath/a_mux/_049_ ;
wire \dpath/a_mux/_050_ ;
wire \dpath/a_mux/_051_ ;
wire \dpath/a_mux/_052_ ;
wire \dpath/a_mux/_053_ ;
wire \dpath/a_mux/_054_ ;
wire \dpath/a_mux/_055_ ;
wire \dpath/a_mux/_056_ ;
wire \dpath/a_mux/_057_ ;
wire \dpath/a_mux/_058_ ;
wire \dpath/a_mux/_059_ ;
wire \dpath/a_mux/_060_ ;
wire \dpath/a_mux/_061_ ;
wire \dpath/a_mux/_062_ ;
wire \dpath/a_mux/_063_ ;
wire \dpath/a_mux/_064_ ;
wire \dpath/a_mux/_065_ ;
wire \dpath/a_mux/_066_ ;
wire \dpath/a_mux/_067_ ;
wire \dpath/a_mux/_068_ ;
wire \dpath/a_mux/_069_ ;
wire \dpath/a_mux/_070_ ;
wire \dpath/a_mux/_071_ ;
wire \dpath/a_mux/_072_ ;
wire \dpath/a_mux/_073_ ;
wire \dpath/a_mux/_074_ ;
wire \dpath/a_mux/_075_ ;
wire \dpath/a_mux/_076_ ;
wire \dpath/a_mux/_077_ ;
wire \dpath/a_mux/_078_ ;
wire \dpath/a_mux/_079_ ;
wire \dpath/a_mux/_080_ ;
wire \dpath/a_mux/_081_ ;
wire \dpath/a_mux/_082_ ;
wire \dpath/a_mux/_083_ ;
wire \dpath/a_mux/_084_ ;
wire \dpath/a_mux/_085_ ;
wire \dpath/a_mux/_086_ ;
wire \dpath/a_mux/_087_ ;
wire \dpath/a_mux/_088_ ;
wire \dpath/a_mux/_089_ ;
wire \dpath/a_mux/_090_ ;
wire \dpath/a_mux/_091_ ;
wire \dpath/a_mux/_092_ ;
wire \dpath/a_mux/_093_ ;
wire \dpath/a_mux/_094_ ;
wire \dpath/a_mux/_095_ ;
wire \dpath/a_mux/_096_ ;
wire \dpath/a_mux/_097_ ;
wire \dpath/a_mux/_098_ ;
wire \dpath/a_mux/_099_ ;
wire \dpath/a_mux/_100_ ;
wire \dpath/a_mux/_101_ ;
wire \dpath/a_mux/_102_ ;
wire \dpath/a_mux/_103_ ;
wire \dpath/a_reg/_000_ ;
wire \dpath/a_reg/_001_ ;
wire \dpath/a_reg/_002_ ;
wire \dpath/a_reg/_003_ ;
wire \dpath/a_reg/_004_ ;
wire \dpath/a_reg/_005_ ;
wire \dpath/a_reg/_006_ ;
wire \dpath/a_reg/_007_ ;
wire \dpath/a_reg/_008_ ;
wire \dpath/a_reg/_009_ ;
wire \dpath/a_reg/_010_ ;
wire \dpath/a_reg/_011_ ;
wire \dpath/a_reg/_012_ ;
wire \dpath/a_reg/_013_ ;
wire \dpath/a_reg/_014_ ;
wire \dpath/a_reg/_015_ ;
wire \dpath/a_reg/_016_ ;
wire \dpath/a_reg/_017_ ;
wire \dpath/a_reg/_018_ ;
wire \dpath/a_reg/_019_ ;
wire \dpath/a_reg/_020_ ;
wire \dpath/a_reg/_021_ ;
wire \dpath/a_reg/_022_ ;
wire \dpath/a_reg/_023_ ;
wire \dpath/a_reg/_024_ ;
wire \dpath/a_reg/_025_ ;
wire \dpath/a_reg/_026_ ;
wire \dpath/a_reg/_027_ ;
wire \dpath/a_reg/_028_ ;
wire \dpath/a_reg/_029_ ;
wire \dpath/a_reg/_030_ ;
wire \dpath/a_reg/_031_ ;
wire \dpath/a_reg/_032_ ;
wire \dpath/a_reg/_033_ ;
wire \dpath/a_reg/_034_ ;
wire \dpath/a_reg/_035_ ;
wire \dpath/a_reg/_036_ ;
wire \dpath/a_reg/_037_ ;
wire \dpath/a_reg/_038_ ;
wire \dpath/a_reg/_039_ ;
wire \dpath/a_reg/_040_ ;
wire \dpath/a_reg/_041_ ;
wire \dpath/a_reg/_042_ ;
wire \dpath/a_reg/_043_ ;
wire \dpath/a_reg/_044_ ;
wire \dpath/a_reg/_045_ ;
wire \dpath/a_reg/_046_ ;
wire \dpath/a_reg/_047_ ;
wire \dpath/a_reg/_048_ ;
wire \dpath/a_reg/_049_ ;
wire \dpath/a_reg/_050_ ;
wire \dpath/a_reg/_051_ ;
wire \dpath/a_reg/_052_ ;
wire \dpath/a_reg/_053_ ;
wire \dpath/a_reg/_054_ ;
wire \dpath/a_reg/_055_ ;
wire \dpath/a_reg/_056_ ;
wire \dpath/a_reg/_057_ ;
wire \dpath/a_reg/_058_ ;
wire \dpath/a_reg/_059_ ;
wire \dpath/a_reg/_060_ ;
wire \dpath/a_reg/_061_ ;
wire \dpath/a_reg/_062_ ;
wire \dpath/a_reg/_063_ ;
wire \dpath/a_reg/_064_ ;
wire \dpath/a_reg/_065_ ;
wire \dpath/b_mux/_000_ ;
wire \dpath/b_mux/_001_ ;
wire \dpath/b_mux/_002_ ;
wire \dpath/b_mux/_003_ ;
wire \dpath/b_mux/_004_ ;
wire \dpath/b_mux/_005_ ;
wire \dpath/b_mux/_006_ ;
wire \dpath/b_mux/_007_ ;
wire \dpath/b_mux/_008_ ;
wire \dpath/b_mux/_009_ ;
wire \dpath/b_mux/_010_ ;
wire \dpath/b_mux/_011_ ;
wire \dpath/b_mux/_012_ ;
wire \dpath/b_mux/_013_ ;
wire \dpath/b_mux/_014_ ;
wire \dpath/b_mux/_015_ ;
wire \dpath/b_mux/_016_ ;
wire \dpath/b_mux/_017_ ;
wire \dpath/b_mux/_018_ ;
wire \dpath/b_mux/_019_ ;
wire \dpath/b_mux/_020_ ;
wire \dpath/b_mux/_021_ ;
wire \dpath/b_mux/_022_ ;
wire \dpath/b_mux/_023_ ;
wire \dpath/b_mux/_024_ ;
wire \dpath/b_mux/_025_ ;
wire \dpath/b_mux/_026_ ;
wire \dpath/b_mux/_027_ ;
wire \dpath/b_mux/_028_ ;
wire \dpath/b_mux/_029_ ;
wire \dpath/b_mux/_030_ ;
wire \dpath/b_mux/_031_ ;
wire \dpath/b_mux/_032_ ;
wire \dpath/b_mux/_033_ ;
wire \dpath/b_mux/_034_ ;
wire \dpath/b_mux/_035_ ;
wire \dpath/b_mux/_036_ ;
wire \dpath/b_mux/_037_ ;
wire \dpath/b_mux/_038_ ;
wire \dpath/b_mux/_039_ ;
wire \dpath/b_mux/_040_ ;
wire \dpath/b_mux/_041_ ;
wire \dpath/b_mux/_042_ ;
wire \dpath/b_mux/_043_ ;
wire \dpath/b_mux/_044_ ;
wire \dpath/b_mux/_045_ ;
wire \dpath/b_mux/_046_ ;
wire \dpath/b_mux/_047_ ;
wire \dpath/b_mux/_048_ ;
wire \dpath/b_mux/_049_ ;
wire \dpath/b_reg/_000_ ;
wire \dpath/b_reg/_001_ ;
wire \dpath/b_reg/_002_ ;
wire \dpath/b_reg/_003_ ;
wire \dpath/b_reg/_004_ ;
wire \dpath/b_reg/_005_ ;
wire \dpath/b_reg/_006_ ;
wire \dpath/b_reg/_007_ ;
wire \dpath/b_reg/_008_ ;
wire \dpath/b_reg/_009_ ;
wire \dpath/b_reg/_010_ ;
wire \dpath/b_reg/_011_ ;
wire \dpath/b_reg/_012_ ;
wire \dpath/b_reg/_013_ ;
wire \dpath/b_reg/_014_ ;
wire \dpath/b_reg/_015_ ;
wire \dpath/b_reg/_016_ ;
wire \dpath/b_reg/_017_ ;
wire \dpath/b_reg/_018_ ;
wire \dpath/b_reg/_019_ ;
wire \dpath/b_reg/_020_ ;
wire \dpath/b_reg/_021_ ;
wire \dpath/b_reg/_022_ ;
wire \dpath/b_reg/_023_ ;
wire \dpath/b_reg/_024_ ;
wire \dpath/b_reg/_025_ ;
wire \dpath/b_reg/_026_ ;
wire \dpath/b_reg/_027_ ;
wire \dpath/b_reg/_028_ ;
wire \dpath/b_reg/_029_ ;
wire \dpath/b_reg/_030_ ;
wire \dpath/b_reg/_031_ ;
wire \dpath/b_reg/_032_ ;
wire \dpath/b_reg/_033_ ;
wire \dpath/b_reg/_034_ ;
wire \dpath/b_reg/_035_ ;
wire \dpath/b_reg/_036_ ;
wire \dpath/b_reg/_037_ ;
wire \dpath/b_reg/_038_ ;
wire \dpath/b_reg/_039_ ;
wire \dpath/b_reg/_040_ ;
wire \dpath/b_reg/_041_ ;
wire \dpath/b_reg/_042_ ;
wire \dpath/b_reg/_043_ ;
wire \dpath/b_reg/_044_ ;
wire \dpath/b_reg/_045_ ;
wire \dpath/b_reg/_046_ ;
wire \dpath/b_reg/_047_ ;
wire \dpath/b_reg/_048_ ;
wire \dpath/b_reg/_049_ ;
wire \dpath/b_reg/_050_ ;
wire \dpath/b_reg/_051_ ;
wire \dpath/b_reg/_052_ ;
wire \dpath/b_reg/_053_ ;
wire \dpath/b_reg/_054_ ;
wire \dpath/b_reg/_055_ ;
wire \dpath/b_reg/_056_ ;
wire \dpath/b_reg/_057_ ;
wire \dpath/b_reg/_058_ ;
wire \dpath/b_reg/_059_ ;
wire \dpath/b_reg/_060_ ;
wire \dpath/b_reg/_061_ ;
wire \dpath/b_reg/_062_ ;
wire \dpath/b_reg/_063_ ;
wire \dpath/b_reg/_064_ ;
wire \dpath/b_reg/_065_ ;
wire \dpath/b_zero/_00_ ;
wire \dpath/b_zero/_01_ ;
wire \dpath/b_zero/_02_ ;
wire \dpath/b_zero/_03_ ;
wire \dpath/b_zero/_04_ ;
wire \dpath/b_zero/_05_ ;
wire \dpath/b_zero/_06_ ;
wire \dpath/b_zero/_07_ ;
wire \dpath/b_zero/_08_ ;
wire \dpath/b_zero/_09_ ;
wire \dpath/b_zero/_10_ ;
wire \dpath/b_zero/_11_ ;
wire \dpath/b_zero/_12_ ;
wire \dpath/b_zero/_13_ ;
wire \dpath/b_zero/_14_ ;
wire \dpath/b_zero/_15_ ;
wire \dpath/b_zero/_16_ ;
wire \dpath/b_zero/_17_ ;
wire \dpath/b_zero/_18_ ;
wire \dpath/b_zero/_19_ ;
wire \dpath/b_zero/_20_ ;
wire \dpath/b_zero/_21_ ;
wire \dpath/b_zero/_22_ ;
wire \dpath/b_zero/_23_ ;
wire \dpath/b_zero/_24_ ;
wire \dpath/sub/_000_ ;
wire \dpath/sub/_001_ ;
wire \dpath/sub/_002_ ;
wire \dpath/sub/_003_ ;
wire \dpath/sub/_004_ ;
wire \dpath/sub/_005_ ;
wire \dpath/sub/_006_ ;
wire \dpath/sub/_007_ ;
wire \dpath/sub/_008_ ;
wire \dpath/sub/_009_ ;
wire \dpath/sub/_010_ ;
wire \dpath/sub/_011_ ;
wire \dpath/sub/_012_ ;
wire \dpath/sub/_013_ ;
wire \dpath/sub/_014_ ;
wire \dpath/sub/_015_ ;
wire \dpath/sub/_016_ ;
wire \dpath/sub/_017_ ;
wire \dpath/sub/_018_ ;
wire \dpath/sub/_019_ ;
wire \dpath/sub/_020_ ;
wire \dpath/sub/_021_ ;
wire \dpath/sub/_022_ ;
wire \dpath/sub/_023_ ;
wire \dpath/sub/_024_ ;
wire \dpath/sub/_025_ ;
wire \dpath/sub/_026_ ;
wire \dpath/sub/_027_ ;
wire \dpath/sub/_028_ ;
wire \dpath/sub/_029_ ;
wire \dpath/sub/_030_ ;
wire \dpath/sub/_031_ ;
wire \dpath/sub/_032_ ;
wire \dpath/sub/_033_ ;
wire \dpath/sub/_034_ ;
wire \dpath/sub/_035_ ;
wire \dpath/sub/_036_ ;
wire \dpath/sub/_037_ ;
wire \dpath/sub/_038_ ;
wire \dpath/sub/_039_ ;
wire \dpath/sub/_040_ ;
wire \dpath/sub/_041_ ;
wire \dpath/sub/_042_ ;
wire \dpath/sub/_043_ ;
wire \dpath/sub/_044_ ;
wire \dpath/sub/_045_ ;
wire \dpath/sub/_046_ ;
wire \dpath/sub/_047_ ;
wire \dpath/sub/_048_ ;
wire \dpath/sub/_049_ ;
wire \dpath/sub/_050_ ;
wire \dpath/sub/_051_ ;
wire \dpath/sub/_052_ ;
wire \dpath/sub/_053_ ;
wire \dpath/sub/_054_ ;
wire \dpath/sub/_055_ ;
wire \dpath/sub/_056_ ;
wire \dpath/sub/_057_ ;
wire \dpath/sub/_058_ ;
wire \dpath/sub/_059_ ;
wire \dpath/sub/_060_ ;
wire \dpath/sub/_061_ ;
wire \dpath/sub/_062_ ;
wire \dpath/sub/_063_ ;
wire \dpath/sub/_064_ ;
wire \dpath/sub/_065_ ;
wire \dpath/sub/_066_ ;
wire \dpath/sub/_067_ ;
wire \dpath/sub/_068_ ;
wire \dpath/sub/_069_ ;
wire \dpath/sub/_070_ ;
wire \dpath/sub/_071_ ;
wire \dpath/sub/_072_ ;
wire \dpath/sub/_073_ ;
wire \dpath/sub/_074_ ;
wire \dpath/sub/_075_ ;
wire \dpath/sub/_076_ ;
wire \dpath/sub/_077_ ;
wire \dpath/sub/_078_ ;
wire \dpath/sub/_079_ ;
wire \dpath/sub/_080_ ;
wire \dpath/sub/_081_ ;
wire \dpath/sub/_082_ ;
wire \dpath/sub/_083_ ;
wire \dpath/sub/_084_ ;
wire \dpath/sub/_085_ ;
wire \dpath/sub/_086_ ;
wire \dpath/sub/_087_ ;
wire \dpath/sub/_088_ ;
wire \dpath/sub/_089_ ;
wire \dpath/sub/_090_ ;
wire \dpath/sub/_091_ ;
wire \dpath/sub/_092_ ;
wire \dpath/sub/_093_ ;
wire \dpath/sub/_094_ ;
wire \dpath/sub/_095_ ;
wire \dpath/sub/_096_ ;
wire \dpath/sub/_097_ ;
wire \dpath/sub/_098_ ;
wire \dpath/sub/_099_ ;
wire \dpath/sub/_100_ ;
wire \dpath/sub/_101_ ;
wire \dpath/sub/_102_ ;
wire \dpath/sub/_103_ ;
wire \dpath/sub/_104_ ;
wire \dpath/sub/_105_ ;
wire \dpath/sub/_106_ ;
wire \dpath/sub/_107_ ;
wire \dpath/sub/_108_ ;
wire \dpath/sub/_109_ ;
wire \dpath/sub/_110_ ;
wire \dpath/sub/_111_ ;
wire \dpath/sub/_112_ ;
wire \dpath/sub/_113_ ;
wire \dpath/sub/_114_ ;
wire \dpath/sub/_115_ ;
wire \dpath/sub/_116_ ;
wire \dpath/sub/_117_ ;
wire \dpath/sub/_118_ ;
wire \dpath/sub/_119_ ;
wire \dpath/sub/_120_ ;
wire req_rdy ;
wire resp_val ;
wire req_val ;
wire resp_rdy ;
wire reset ;
wire clk ;
wire clk_86 ;
wire clk_85 ;
wire clk_84 ;
wire clk_83 ;
wire clk_82 ;
wire clk_81 ;
wire clk_80 ;
wire clk_79 ;
wire clk_78 ;
wire clk_77 ;
wire clk_76 ;
wire clk_75 ;
wire clk_74 ;
wire clk_73 ;
wire clk_72 ;
wire clk_71 ;
wire clk_70 ;
wire clk_69 ;
wire clk_68 ;
wire clk_67 ;
wire clk_66 ;
wire clk_65 ;
wire clk_64 ;
wire clk_63 ;
wire clk_62 ;
wire clk_61 ;
wire clk_60 ;
wire clk_59 ;
wire clk_58 ;
wire clk_57 ;
wire clk_56 ;
wire clk_55 ;
wire clk_54 ;
wire clk_53 ;
wire clk_52 ;
wire clk_51 ;
wire clk_50 ;
wire clk_49 ;
wire clk_48 ;
wire clk_47 ;
wire clk_46 ;
wire clk_45 ;
wire clk_44 ;
wire clk_43 ;
wire clk_42 ;
wire clk_41 ;
wire clk_40 ;
wire clk_39 ;
wire clk_38 ;
wire clk_37 ;
wire clk_36 ;
wire clk_35 ;
wire clk_34 ;
wire clk_33 ;
wire clk_32 ;
wire clk_31 ;
wire clk_30 ;
wire clk_29 ;
wire clk_28 ;
wire clk_27 ;
wire clk_26 ;
wire clk_25 ;
wire clk_24 ;
wire clk_23 ;
wire clk_22 ;
wire clk_21 ;
wire clk_20 ;
wire clk_19 ;
wire clk_18 ;
wire clk_17 ;
wire clk_16 ;
wire clk_15 ;
wire clk_14 ;
wire clk_13 ;
wire clk_12 ;
wire clk_11 ;
wire clk_10 ;
wire clk_9 ;
wire clk_8 ;
wire clk_7 ;
wire clk_6 ;
wire clk_5 ;
wire clk_4 ;
wire clk_3 ;
wire clk_2 ;
wire clk_1 ;
wire clk_0 ;
wire [1:0] ctrl$a_mux_sel ;
wire [1:0] \ctrl/curr_state__0 ;
wire [1:0] \ctrl/next_state__0 ;
wire [15:0] \dpath/a_lt_b$in0 ;
wire [15:0] \dpath/a_lt_b$in1 ;
wire [15:0] \dpath/a_mux$out ;
wire [15:0] \dpath/b_mux$out ;
wire [15:0] resp_msg ;
wire [31:0] req_msg ;

sky130_fd_sc_hs__nor2_1 \ctrl/_17_ ( .A(\ctrl/_05_ ), .B(\ctrl/_06_ ), .Y(\ctrl/_03_ ) );
sky130_fd_sc_hs__and2b_1 \ctrl/_18_ ( .A_N(\ctrl/_05_ ), .B(\ctrl/_06_ ), .X(\ctrl/_16_ ) );
sky130_fd_sc_hs__nor3b_1 \ctrl/_19_ ( .A(\ctrl/_06_ ), .B(\ctrl/_07_ ), .C_N(\ctrl/_05_ ), .Y(\ctrl/_00_ ) );
sky130_fd_sc_hs__and3b_1 \ctrl/_20_ ( .A_N(\ctrl/_06_ ), .B(\ctrl/_05_ ), .C(\ctrl/_07_ ), .X(\ctrl/_01_ ) );
sky130_fd_sc_hs__nor3b_1 \ctrl/_21_ ( .A(\ctrl/_05_ ), .B(\ctrl/_06_ ), .C_N(\ctrl/_14_ ), .Y(\ctrl/_09_ ) );
sky130_fd_sc_hs__nor2b_4 \ctrl/_22_ ( .A(\ctrl/_07_ ), .B_N(\ctrl/_08_ ), .Y(\ctrl/_10_ ) );
sky130_fd_sc_hs__inv_1 \ctrl/_23_ ( .A(\ctrl/_06_ ), .Y(\ctrl/_02_ ) );
sky130_fd_sc_hs__nand3_2 \ctrl/_24_ ( .A(\ctrl/_10_ ), .B(\ctrl/_05_ ), .C(\ctrl/_02_ ), .Y(\ctrl/_11_ ) );
sky130_fd_sc_hs__o21a_1 \ctrl/_25_ ( .A1(\ctrl/_05_ ), .A2(\ctrl/_09_ ), .B1(\ctrl/_11_ ), .X(\ctrl/_12_ ) );
sky130_fd_sc_hs__a22oi_1 \ctrl/_26_ ( .A1(\ctrl/_15_ ), .A2(\ctrl/_16_ ), .B1(\ctrl/_11_ ), .B2(\ctrl/_02_ ), .Y(\ctrl/_13_ ) );
sky130_fd_sc_hs__o21bai_1 \ctrl/_27_ ( .A1(\ctrl/_05_ ), .A2(\ctrl/_06_ ), .B1_N(\ctrl/_01_ ), .Y(\ctrl/_04_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/_28_ ( .A(ctrl$b_mux_sel ), .X(req_rdy ) );
sky130_fd_sc_hs__buf_1 \ctrl/_29_ ( .A(\ctrl/curr_state__0[0] ), .X(\ctrl/_05_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/_30_ ( .A(\ctrl/curr_state__0[1] ), .X(\ctrl/_06_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/_31_ ( .A(\ctrl/_03_ ), .X(ctrl$b_mux_sel ) );
sky130_fd_sc_hs__buf_1 \ctrl/_32_ ( .A(\ctrl/_16_ ), .X(resp_val ) );
sky130_fd_sc_hs__buf_1 \ctrl/_33_ ( .A(ctrl$is_a_lt_b ), .X(\ctrl/_07_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/_34_ ( .A(\ctrl/_00_ ), .X(\ctrl$a_mux_sel[0] ) );
sky130_fd_sc_hs__buf_1 \ctrl/_35_ ( .A(\ctrl/_01_ ), .X(\ctrl$a_mux_sel[1] ) );
sky130_fd_sc_hs__buf_1 \ctrl/_36_ ( .A(req_val ), .X(\ctrl/_14_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/_37_ ( .A(ctrl$is_b_zero ), .X(\ctrl/_08_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/_38_ ( .A(resp_rdy ), .X(\ctrl/_15_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/_39_ ( .A(\ctrl/_12_ ), .X(\ctrl/next_state__0[0] ) );
sky130_fd_sc_hs__buf_1 \ctrl/_40_ ( .A(\ctrl/_13_ ), .X(\ctrl/next_state__0[1] ) );
sky130_fd_sc_hs__buf_1 \ctrl/_41_ ( .A(\ctrl/_04_ ), .X(ctrl$b_reg_en ) );
sky130_fd_sc_hs__buf_1 \ctrl/_42_ ( .A(\ctrl/_02_ ), .X(ctrl$a_reg_en ) );
sky130_fd_sc_hs__nor2b_2 \ctrl/state/_07_ ( .A(\ctrl/state/_06_ ), .B_N(\ctrl/state/_04_ ), .Y(\ctrl/state/_02_ ) );
sky130_fd_sc_hs__nor2b_2 \ctrl/state/_08_ ( .A(\ctrl/state/_06_ ), .B_N(\ctrl/state/_05_ ), .Y(\ctrl/state/_03_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/state/_09_ ( .A(\ctrl/next_state__0[0] ), .X(\ctrl/state/_04_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/state/_10_ ( .A(reset ), .X(\ctrl/state/_06_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/state/_11_ ( .A(\ctrl/state/_02_ ), .X(\ctrl/state/_00_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/state/_12_ ( .A(\ctrl/next_state__0[1] ), .X(\ctrl/state/_05_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/state/_13_ ( .A(\ctrl/state/_03_ ), .X(\ctrl/state/_01_ ) );
sky130_fd_sc_hs__dfxtp_1 \ctrl/state/_14_ ( .D(\ctrl/state/_00_ ), .Q(\ctrl/curr_state__0[0] ), .CLK(clk_85 ) );
sky130_fd_sc_hs__dfxtp_1 \ctrl/state/_15_ ( .D(\ctrl/state/_01_ ), .Q(\ctrl/curr_state__0[1] ), .CLK(clk_85 ) );
sky130_fd_sc_hs__nor2b_2 \dpath/a_lt_b/_090_ ( .A(\dpath/a_lt_b/_025_ ), .B_N(\dpath/a_lt_b/_009_ ), .Y(\dpath/a_lt_b/_032_ ) );
sky130_fd_sc_hs__nand2b_2 \dpath/a_lt_b/_091_ ( .A_N(\dpath/a_lt_b/_009_ ), .B(\dpath/a_lt_b/_025_ ), .Y(\dpath/a_lt_b/_033_ ) );
sky130_fd_sc_hs__and3b_1 \dpath/a_lt_b/_092_ ( .A_N(\dpath/a_lt_b/_024_ ), .B(\dpath/a_lt_b/_033_ ), .C(\dpath/a_lt_b/_008_ ), .X(\dpath/a_lt_b/_034_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/a_lt_b/_093_ ( .A(\dpath/a_lt_b/_024_ ), .B(\dpath/a_lt_b/_008_ ), .Y(\dpath/a_lt_b/_035_ ) );
sky130_fd_sc_hs__and3b_1 \dpath/a_lt_b/_094_ ( .A_N(\dpath/a_lt_b/_032_ ), .B(\dpath/a_lt_b/_035_ ), .C(\dpath/a_lt_b/_033_ ), .X(\dpath/a_lt_b/_036_ ) );
sky130_fd_sc_hs__inv_8 \dpath/a_lt_b/_095_ ( .A(\dpath/a_lt_b/_023_ ), .Y(\dpath/a_lt_b/_037_ ) );
sky130_fd_sc_hs__nand2b_4 \dpath/a_lt_b/_096_ ( .A_N(\dpath/a_lt_b/_000_ ), .B(\dpath/a_lt_b/_016_ ), .Y(\dpath/a_lt_b/_038_ ) );
sky130_fd_sc_hs__maj3_1 \dpath/a_lt_b/_097_ ( .A(\dpath/a_lt_b/_037_ ), .B(\dpath/a_lt_b/_038_ ), .C(\dpath/a_lt_b/_007_ ), .X(\dpath/a_lt_b/_039_ ) );
sky130_fd_sc_hs__and2_1 \dpath/a_lt_b/_098_ ( .A(\dpath/a_lt_b/_036_ ), .B(\dpath/a_lt_b/_039_ ), .X(\dpath/a_lt_b/_040_ ) );
sky130_fd_sc_hs__inv_1 \dpath/a_lt_b/_099_ ( .A(\dpath/a_lt_b/_026_ ), .Y(\dpath/a_lt_b/_041_ ) );
sky130_fd_sc_hs__nor2b_1 \dpath/a_lt_b/_100_ ( .A(\dpath/a_lt_b/_027_ ), .B_N(\dpath/a_lt_b/_011_ ), .Y(\dpath/a_lt_b/_042_ ) );
sky130_fd_sc_hs__a21o_1 \dpath/a_lt_b/_101_ ( .A1(\dpath/a_lt_b/_010_ ), .A2(\dpath/a_lt_b/_041_ ), .B1(\dpath/a_lt_b/_042_ ), .X(\dpath/a_lt_b/_043_ ) );
sky130_fd_sc_hs__nor2b_4 \dpath/a_lt_b/_102_ ( .A(\dpath/a_lt_b/_013_ ), .B_N(\dpath/a_lt_b/_029_ ), .Y(\dpath/a_lt_b/_044_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/a_lt_b/_103_ ( .A(\dpath/a_lt_b/_028_ ), .B(\dpath/a_lt_b/_012_ ), .Y(\dpath/a_lt_b/_045_ ) );
sky130_fd_sc_hs__nand2b_1 \dpath/a_lt_b/_104_ ( .A_N(\dpath/a_lt_b/_029_ ), .B(\dpath/a_lt_b/_013_ ), .Y(\dpath/a_lt_b/_046_ ) );
sky130_fd_sc_hs__and3b_1 \dpath/a_lt_b/_105_ ( .A_N(\dpath/a_lt_b/_044_ ), .B(\dpath/a_lt_b/_045_ ), .C(\dpath/a_lt_b/_046_ ), .X(\dpath/a_lt_b/_047_ ) );
sky130_fd_sc_hs__nor2b_4 \dpath/a_lt_b/_106_ ( .A(\dpath/a_lt_b/_011_ ), .B_N(\dpath/a_lt_b/_027_ ), .Y(\dpath/a_lt_b/_048_ ) );
sky130_fd_sc_hs__o21ba_1 \dpath/a_lt_b/_107_ ( .A1(\dpath/a_lt_b/_010_ ), .A2(\dpath/a_lt_b/_041_ ), .B1_N(\dpath/a_lt_b/_048_ ), .X(\dpath/a_lt_b/_049_ ) );
sky130_fd_sc_hs__and3b_1 \dpath/a_lt_b/_108_ ( .A_N(\dpath/a_lt_b/_043_ ), .B(\dpath/a_lt_b/_047_ ), .C(\dpath/a_lt_b/_049_ ), .X(\dpath/a_lt_b/_050_ ) );
sky130_fd_sc_hs__o31ai_1 \dpath/a_lt_b/_109_ ( .A1(\dpath/a_lt_b/_032_ ), .A2(\dpath/a_lt_b/_034_ ), .A3(\dpath/a_lt_b/_040_ ), .B1(\dpath/a_lt_b/_050_ ), .Y(\dpath/a_lt_b/_051_ ) );
sky130_fd_sc_hs__nor2b_2 \dpath/a_lt_b/_110_ ( .A(\dpath/a_lt_b/_028_ ), .B_N(\dpath/a_lt_b/_012_ ), .Y(\dpath/a_lt_b/_052_ ) );
sky130_fd_sc_hs__nor2b_1 \dpath/a_lt_b/_111_ ( .A(\dpath/a_lt_b/_052_ ), .B_N(\dpath/a_lt_b/_046_ ), .Y(\dpath/a_lt_b/_053_ ) );
sky130_fd_sc_hs__or2_1 \dpath/a_lt_b/_112_ ( .A(\dpath/a_lt_b/_044_ ), .B(\dpath/a_lt_b/_053_ ), .X(\dpath/a_lt_b/_054_ ) );
sky130_fd_sc_hs__nand3b_1 \dpath/a_lt_b/_113_ ( .A_N(\dpath/a_lt_b/_048_ ), .B(\dpath/a_lt_b/_047_ ), .C(\dpath/a_lt_b/_043_ ), .Y(\dpath/a_lt_b/_055_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/a_lt_b/_114_ ( .A(\dpath/a_lt_b/_020_ ), .B_N(\dpath/a_lt_b/_004_ ), .X(\dpath/a_lt_b/_056_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/a_lt_b/_115_ ( .A(\dpath/a_lt_b/_019_ ), .B_N(\dpath/a_lt_b/_003_ ), .X(\dpath/a_lt_b/_057_ ) );
sky130_fd_sc_hs__nand2_2 \dpath/a_lt_b/_116_ ( .A(\dpath/a_lt_b/_056_ ), .B(\dpath/a_lt_b/_057_ ), .Y(\dpath/a_lt_b/_058_ ) );
sky130_fd_sc_hs__and2b_2 \dpath/a_lt_b/_117_ ( .A_N(\dpath/a_lt_b/_005_ ), .B(\dpath/a_lt_b/_021_ ), .X(\dpath/a_lt_b/_059_ ) );
sky130_fd_sc_hs__nor2b_2 \dpath/a_lt_b/_118_ ( .A(\dpath/a_lt_b/_006_ ), .B_N(\dpath/a_lt_b/_022_ ), .Y(\dpath/a_lt_b/_060_ ) );
sky130_fd_sc_hs__nand2b_2 \dpath/a_lt_b/_119_ ( .A_N(\dpath/a_lt_b/_021_ ), .B(\dpath/a_lt_b/_005_ ), .Y(\dpath/a_lt_b/_061_ ) );
sky130_fd_sc_hs__nand2b_4 \dpath/a_lt_b/_120_ ( .A_N(\dpath/a_lt_b/_022_ ), .B(\dpath/a_lt_b/_006_ ), .Y(\dpath/a_lt_b/_062_ ) );
sky130_fd_sc_hs__nand3b_1 \dpath/a_lt_b/_121_ ( .A_N(\dpath/a_lt_b/_060_ ), .B(\dpath/a_lt_b/_061_ ), .C(\dpath/a_lt_b/_062_ ), .Y(\dpath/a_lt_b/_063_ ) );
sky130_fd_sc_hs__nor2_2 \dpath/a_lt_b/_122_ ( .A(\dpath/a_lt_b/_059_ ), .B(\dpath/a_lt_b/_063_ ), .Y(\dpath/a_lt_b/_064_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/a_lt_b/_123_ ( .A(\dpath/a_lt_b/_004_ ), .B_N(\dpath/a_lt_b/_020_ ), .X(\dpath/a_lt_b/_065_ ) );
sky130_fd_sc_hs__or2b_4 \dpath/a_lt_b/_124_ ( .A(\dpath/a_lt_b/_003_ ), .B_N(\dpath/a_lt_b/_019_ ), .X(\dpath/a_lt_b/_066_ ) );
sky130_fd_sc_hs__nand3_2 \dpath/a_lt_b/_125_ ( .A(\dpath/a_lt_b/_064_ ), .B(\dpath/a_lt_b/_065_ ), .C(\dpath/a_lt_b/_066_ ), .Y(\dpath/a_lt_b/_067_ ) );
sky130_fd_sc_hs__or2_1 \dpath/a_lt_b/_126_ ( .A(\dpath/a_lt_b/_058_ ), .B(\dpath/a_lt_b/_067_ ), .X(\dpath/a_lt_b/_068_ ) );
sky130_fd_sc_hs__inv_1 \dpath/a_lt_b/_127_ ( .A(\dpath/a_lt_b/_001_ ), .Y(\dpath/a_lt_b/_069_ ) );
sky130_fd_sc_hs__nor2b_4 \dpath/a_lt_b/_128_ ( .A(\dpath/a_lt_b/_018_ ), .B_N(\dpath/a_lt_b/_002_ ), .Y(\dpath/a_lt_b/_070_ ) );
sky130_fd_sc_hs__nor2b_4 \dpath/a_lt_b/_129_ ( .A(\dpath/a_lt_b/_017_ ), .B_N(\dpath/a_lt_b/_001_ ), .Y(\dpath/a_lt_b/_071_ ) );
sky130_fd_sc_hs__nor2b_2 \dpath/a_lt_b/_130_ ( .A(\dpath/a_lt_b/_002_ ), .B_N(\dpath/a_lt_b/_018_ ), .Y(\dpath/a_lt_b/_072_ ) );
sky130_fd_sc_hs__or3_1 \dpath/a_lt_b/_131_ ( .A(\dpath/a_lt_b/_070_ ), .B(\dpath/a_lt_b/_071_ ), .C(\dpath/a_lt_b/_072_ ), .X(\dpath/a_lt_b/_073_ ) );
sky130_fd_sc_hs__a21oi_4 \dpath/a_lt_b/_132_ ( .A1(\dpath/a_lt_b/_017_ ), .A2(\dpath/a_lt_b/_069_ ), .B1(\dpath/a_lt_b/_073_ ), .Y(\dpath/a_lt_b/_074_ ) );
sky130_fd_sc_hs__and2b_2 \dpath/a_lt_b/_133_ ( .A_N(\dpath/a_lt_b/_015_ ), .B(\dpath/a_lt_b/_031_ ), .X(\dpath/a_lt_b/_075_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/a_lt_b/_134_ ( .A(\dpath/a_lt_b/_014_ ), .B(\dpath/a_lt_b/_030_ ), .Y(\dpath/a_lt_b/_076_ ) );
sky130_fd_sc_hs__or2b_2 \dpath/a_lt_b/_135_ ( .A(\dpath/a_lt_b/_031_ ), .B_N(\dpath/a_lt_b/_015_ ), .X(\dpath/a_lt_b/_077_ ) );
sky130_fd_sc_hs__and3b_1 \dpath/a_lt_b/_136_ ( .A_N(\dpath/a_lt_b/_075_ ), .B(\dpath/a_lt_b/_076_ ), .C(\dpath/a_lt_b/_077_ ), .X(\dpath/a_lt_b/_078_ ) );
sky130_fd_sc_hs__nand3b_1 \dpath/a_lt_b/_137_ ( .A_N(\dpath/a_lt_b/_068_ ), .B(\dpath/a_lt_b/_074_ ), .C(\dpath/a_lt_b/_078_ ), .Y(\dpath/a_lt_b/_079_ ) );
sky130_fd_sc_hs__a31o_1 \dpath/a_lt_b/_138_ ( .A1(\dpath/a_lt_b/_051_ ), .A2(\dpath/a_lt_b/_054_ ), .A3(\dpath/a_lt_b/_055_ ), .B1(\dpath/a_lt_b/_079_ ), .X(\dpath/a_lt_b/_080_ ) );
sky130_fd_sc_hs__nor3b_1 \dpath/a_lt_b/_139_ ( .A(\dpath/a_lt_b/_070_ ), .B(\dpath/a_lt_b/_072_ ), .C_N(\dpath/a_lt_b/_071_ ), .Y(\dpath/a_lt_b/_081_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/a_lt_b/_140_ ( .A(\dpath/a_lt_b/_030_ ), .B_N(\dpath/a_lt_b/_014_ ), .X(\dpath/a_lt_b/_082_ ) );
sky130_fd_sc_hs__a21oi_1 \dpath/a_lt_b/_141_ ( .A1(\dpath/a_lt_b/_077_ ), .A2(\dpath/a_lt_b/_082_ ), .B1(\dpath/a_lt_b/_075_ ), .Y(\dpath/a_lt_b/_083_ ) );
sky130_fd_sc_hs__and2_1 \dpath/a_lt_b/_142_ ( .A(\dpath/a_lt_b/_074_ ), .B(\dpath/a_lt_b/_083_ ), .X(\dpath/a_lt_b/_084_ ) );
sky130_fd_sc_hs__nor2_1 \dpath/a_lt_b/_143_ ( .A(\dpath/a_lt_b/_058_ ), .B(\dpath/a_lt_b/_067_ ), .Y(\dpath/a_lt_b/_085_ ) );
sky130_fd_sc_hs__o31ai_1 \dpath/a_lt_b/_144_ ( .A1(\dpath/a_lt_b/_070_ ), .A2(\dpath/a_lt_b/_081_ ), .A3(\dpath/a_lt_b/_084_ ), .B1(\dpath/a_lt_b/_085_ ), .Y(\dpath/a_lt_b/_086_ ) );
sky130_fd_sc_hs__a21o_1 \dpath/a_lt_b/_145_ ( .A1(\dpath/a_lt_b/_061_ ), .A2(\dpath/a_lt_b/_062_ ), .B1(\dpath/a_lt_b/_060_ ), .X(\dpath/a_lt_b/_087_ ) );
sky130_fd_sc_hs__nand3_1 \dpath/a_lt_b/_146_ ( .A(\dpath/a_lt_b/_064_ ), .B(\dpath/a_lt_b/_058_ ), .C(\dpath/a_lt_b/_065_ ), .Y(\dpath/a_lt_b/_088_ ) );
sky130_fd_sc_hs__and4_1 \dpath/a_lt_b/_147_ ( .A(\dpath/a_lt_b/_080_ ), .B(\dpath/a_lt_b/_086_ ), .C(\dpath/a_lt_b/_087_ ), .D(\dpath/a_lt_b/_088_ ), .X(\dpath/a_lt_b/_089_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_148_ ( .A(\dpath/a_lt_b$in0[8] ), .X(\dpath/a_lt_b/_014_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_149_ ( .A(\dpath/a_lt_b$in1[8] ), .X(\dpath/a_lt_b/_030_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_150_ ( .A(\dpath/a_lt_b$in1[7] ), .X(\dpath/a_lt_b/_029_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_151_ ( .A(\dpath/a_lt_b$in0[7] ), .X(\dpath/a_lt_b/_013_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_152_ ( .A(\dpath/a_lt_b$in1[6] ), .X(\dpath/a_lt_b/_028_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_153_ ( .A(\dpath/a_lt_b$in0[6] ), .X(\dpath/a_lt_b/_012_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_154_ ( .A(\dpath/a_lt_b$in1[5] ), .X(\dpath/a_lt_b/_027_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_155_ ( .A(\dpath/a_lt_b$in0[5] ), .X(\dpath/a_lt_b/_011_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_156_ ( .A(\dpath/a_lt_b$in0[4] ), .X(\dpath/a_lt_b/_010_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_157_ ( .A(\dpath/a_lt_b$in1[4] ), .X(\dpath/a_lt_b/_026_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_158_ ( .A(\dpath/a_lt_b$in1[3] ), .X(\dpath/a_lt_b/_025_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_159_ ( .A(\dpath/a_lt_b$in0[3] ), .X(\dpath/a_lt_b/_009_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_160_ ( .A(\dpath/a_lt_b$in1[2] ), .X(\dpath/a_lt_b/_024_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_161_ ( .A(\dpath/a_lt_b$in0[2] ), .X(\dpath/a_lt_b/_008_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_162_ ( .A(\dpath/a_lt_b$in1[1] ), .X(\dpath/a_lt_b/_023_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_163_ ( .A(\dpath/a_lt_b$in0[1] ), .X(\dpath/a_lt_b/_007_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_164_ ( .A(\dpath/a_lt_b$in1[0] ), .X(\dpath/a_lt_b/_016_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_165_ ( .A(\dpath/a_lt_b$in0[0] ), .X(\dpath/a_lt_b/_000_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_166_ ( .A(\dpath/a_lt_b/_089_ ), .X(ctrl$is_a_lt_b ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_167_ ( .A(\dpath/a_lt_b$in1[15] ), .X(\dpath/a_lt_b/_022_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_168_ ( .A(\dpath/a_lt_b$in0[15] ), .X(\dpath/a_lt_b/_006_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_169_ ( .A(\dpath/a_lt_b$in1[14] ), .X(\dpath/a_lt_b/_021_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_170_ ( .A(\dpath/a_lt_b$in0[14] ), .X(\dpath/a_lt_b/_005_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_171_ ( .A(\dpath/a_lt_b$in1[13] ), .X(\dpath/a_lt_b/_020_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_172_ ( .A(\dpath/a_lt_b$in0[13] ), .X(\dpath/a_lt_b/_004_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_173_ ( .A(\dpath/a_lt_b$in0[12] ), .X(\dpath/a_lt_b/_003_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_174_ ( .A(\dpath/a_lt_b$in1[12] ), .X(\dpath/a_lt_b/_019_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_175_ ( .A(\dpath/a_lt_b$in1[11] ), .X(\dpath/a_lt_b/_018_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_176_ ( .A(\dpath/a_lt_b$in0[11] ), .X(\dpath/a_lt_b/_002_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_177_ ( .A(\dpath/a_lt_b$in1[10] ), .X(\dpath/a_lt_b/_017_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_178_ ( .A(\dpath/a_lt_b$in0[10] ), .X(\dpath/a_lt_b/_001_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_179_ ( .A(\dpath/a_lt_b$in1[9] ), .X(\dpath/a_lt_b/_031_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_180_ ( .A(\dpath/a_lt_b$in0[9] ), .X(\dpath/a_lt_b/_015_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_104_ ( .A(\dpath/a_mux/_000_ ), .Y(\dpath/a_mux/_062_ ) );
sky130_fd_sc_hs__xor2_4 \dpath/a_mux/_105_ ( .A(\dpath/a_mux/_102_ ), .B(\dpath/a_mux/_103_ ), .X(\dpath/a_mux/_063_ ) );
sky130_fd_sc_hs__buf_4 \dpath/a_mux/_106_ ( .A(\dpath/a_mux/_063_ ), .X(\dpath/a_mux/_064_ ) );
sky130_fd_sc_hs__and2b_4 \dpath/a_mux/_107_ ( .A_N(\dpath/a_mux/_103_ ), .B(\dpath/a_mux/_102_ ), .X(\dpath/a_mux/_065_ ) );
sky130_fd_sc_hs__buf_16 \dpath/a_mux/_108_ ( .A(\dpath/a_mux/_065_ ), .X(\dpath/a_mux/_066_ ) );
sky130_fd_sc_hs__and2b_4 \dpath/a_mux/_109_ ( .A_N(\dpath/a_mux/_102_ ), .B(\dpath/a_mux/_103_ ), .X(\dpath/a_mux/_067_ ) );
sky130_fd_sc_hs__buf_8 \dpath/a_mux/_110_ ( .A(\dpath/a_mux/_067_ ), .X(\dpath/a_mux/_068_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_111_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_016_ ), .B1(\dpath/a_mux/_032_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_069_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_112_ ( .A1(\dpath/a_mux/_062_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_069_ ), .Y(\dpath/a_mux/_086_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_113_ ( .A(\dpath/a_mux/_007_ ), .Y(\dpath/a_mux/_070_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_114_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_023_ ), .B1(\dpath/a_mux/_039_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_071_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_115_ ( .A1(\dpath/a_mux/_070_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_071_ ), .Y(\dpath/a_mux/_093_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_116_ ( .A(\dpath/a_mux/_008_ ), .Y(\dpath/a_mux/_072_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_117_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_024_ ), .B1(\dpath/a_mux/_040_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_073_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_118_ ( .A1(\dpath/a_mux/_072_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_073_ ), .Y(\dpath/a_mux/_094_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_119_ ( .A(\dpath/a_mux/_009_ ), .Y(\dpath/a_mux/_074_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_120_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_025_ ), .B1(\dpath/a_mux/_041_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_075_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_121_ ( .A1(\dpath/a_mux/_074_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_075_ ), .Y(\dpath/a_mux/_095_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_122_ ( .A(\dpath/a_mux/_010_ ), .Y(\dpath/a_mux/_076_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_123_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_026_ ), .B1(\dpath/a_mux/_042_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_077_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_124_ ( .A1(\dpath/a_mux/_076_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_077_ ), .Y(\dpath/a_mux/_096_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_125_ ( .A(\dpath/a_mux/_011_ ), .Y(\dpath/a_mux/_078_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_126_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_027_ ), .B1(\dpath/a_mux/_043_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_079_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_127_ ( .A1(\dpath/a_mux/_078_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_079_ ), .Y(\dpath/a_mux/_097_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_128_ ( .A(\dpath/a_mux/_012_ ), .Y(\dpath/a_mux/_080_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_129_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_028_ ), .B1(\dpath/a_mux/_044_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_081_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_130_ ( .A1(\dpath/a_mux/_080_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_081_ ), .Y(\dpath/a_mux/_098_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_131_ ( .A(\dpath/a_mux/_013_ ), .Y(\dpath/a_mux/_082_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_132_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_029_ ), .B1(\dpath/a_mux/_045_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_083_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_133_ ( .A1(\dpath/a_mux/_082_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_083_ ), .Y(\dpath/a_mux/_099_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_134_ ( .A(\dpath/a_mux/_014_ ), .Y(\dpath/a_mux/_084_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_135_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_030_ ), .B1(\dpath/a_mux/_046_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_085_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_136_ ( .A1(\dpath/a_mux/_084_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_085_ ), .Y(\dpath/a_mux/_100_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_137_ ( .A(\dpath/a_mux/_015_ ), .Y(\dpath/a_mux/_048_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_138_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_031_ ), .B1(\dpath/a_mux/_047_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_049_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_139_ ( .A1(\dpath/a_mux/_048_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_049_ ), .Y(\dpath/a_mux/_101_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_140_ ( .A(\dpath/a_mux/_001_ ), .Y(\dpath/a_mux/_050_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_141_ ( .A1(\dpath/a_mux/_065_ ), .A2(\dpath/a_mux/_017_ ), .B1(\dpath/a_mux/_033_ ), .B2(\dpath/a_mux/_067_ ), .Y(\dpath/a_mux/_051_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_142_ ( .A1(\dpath/a_mux/_050_ ), .A2(\dpath/a_mux/_063_ ), .B1(\dpath/a_mux/_051_ ), .Y(\dpath/a_mux/_087_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_143_ ( .A(\dpath/a_mux/_002_ ), .Y(\dpath/a_mux/_052_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_144_ ( .A1(\dpath/a_mux/_065_ ), .A2(\dpath/a_mux/_018_ ), .B1(\dpath/a_mux/_034_ ), .B2(\dpath/a_mux/_067_ ), .Y(\dpath/a_mux/_053_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_145_ ( .A1(\dpath/a_mux/_052_ ), .A2(\dpath/a_mux/_063_ ), .B1(\dpath/a_mux/_053_ ), .Y(\dpath/a_mux/_088_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_146_ ( .A(\dpath/a_mux/_003_ ), .Y(\dpath/a_mux/_054_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_147_ ( .A1(\dpath/a_mux/_065_ ), .A2(\dpath/a_mux/_019_ ), .B1(\dpath/a_mux/_035_ ), .B2(\dpath/a_mux/_067_ ), .Y(\dpath/a_mux/_055_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_148_ ( .A1(\dpath/a_mux/_054_ ), .A2(\dpath/a_mux/_063_ ), .B1(\dpath/a_mux/_055_ ), .Y(\dpath/a_mux/_089_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_149_ ( .A(\dpath/a_mux/_004_ ), .Y(\dpath/a_mux/_056_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_150_ ( .A1(\dpath/a_mux/_065_ ), .A2(\dpath/a_mux/_020_ ), .B1(\dpath/a_mux/_036_ ), .B2(\dpath/a_mux/_067_ ), .Y(\dpath/a_mux/_057_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_151_ ( .A1(\dpath/a_mux/_056_ ), .A2(\dpath/a_mux/_063_ ), .B1(\dpath/a_mux/_057_ ), .Y(\dpath/a_mux/_090_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_152_ ( .A(\dpath/a_mux/_005_ ), .Y(\dpath/a_mux/_058_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_153_ ( .A1(\dpath/a_mux/_065_ ), .A2(\dpath/a_mux/_021_ ), .B1(\dpath/a_mux/_037_ ), .B2(\dpath/a_mux/_067_ ), .Y(\dpath/a_mux/_059_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_154_ ( .A1(\dpath/a_mux/_058_ ), .A2(\dpath/a_mux/_063_ ), .B1(\dpath/a_mux/_059_ ), .Y(\dpath/a_mux/_091_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_155_ ( .A(\dpath/a_mux/_006_ ), .Y(\dpath/a_mux/_060_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_156_ ( .A1(\dpath/a_mux/_065_ ), .A2(\dpath/a_mux/_022_ ), .B1(\dpath/a_mux/_038_ ), .B2(\dpath/a_mux/_067_ ), .Y(\dpath/a_mux/_061_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_157_ ( .A1(\dpath/a_mux/_060_ ), .A2(\dpath/a_mux/_063_ ), .B1(\dpath/a_mux/_061_ ), .Y(\dpath/a_mux/_092_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_158_ ( .A(\ctrl$a_mux_sel[0] ), .X(\dpath/a_mux/_102_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_159_ ( .A(\ctrl$a_mux_sel[1] ), .X(\dpath/a_mux/_103_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_160_ ( .A(\dpath/a_lt_b$in1[0] ), .X(\dpath/a_mux/_032_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_161_ ( .A(\resp_msg[0] ), .X(\dpath/a_mux/_016_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_162_ ( .A(\req_msg[16] ), .X(\dpath/a_mux/_000_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_163_ ( .A(\dpath/a_mux/_086_ ), .X(\dpath/a_mux$out[0] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_164_ ( .A(\dpath/a_lt_b$in1[1] ), .X(\dpath/a_mux/_039_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_165_ ( .A(\resp_msg[1] ), .X(\dpath/a_mux/_023_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_166_ ( .A(\req_msg[17] ), .X(\dpath/a_mux/_007_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_167_ ( .A(\dpath/a_mux/_093_ ), .X(\dpath/a_mux$out[1] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_168_ ( .A(\dpath/a_lt_b$in1[2] ), .X(\dpath/a_mux/_040_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_169_ ( .A(\resp_msg[2] ), .X(\dpath/a_mux/_024_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_170_ ( .A(\req_msg[18] ), .X(\dpath/a_mux/_008_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_171_ ( .A(\dpath/a_mux/_094_ ), .X(\dpath/a_mux$out[2] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_172_ ( .A(\dpath/a_lt_b$in1[3] ), .X(\dpath/a_mux/_041_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_173_ ( .A(\resp_msg[3] ), .X(\dpath/a_mux/_025_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_174_ ( .A(\req_msg[19] ), .X(\dpath/a_mux/_009_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_175_ ( .A(\dpath/a_mux/_095_ ), .X(\dpath/a_mux$out[3] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_176_ ( .A(\dpath/a_lt_b$in1[4] ), .X(\dpath/a_mux/_042_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_177_ ( .A(\resp_msg[4] ), .X(\dpath/a_mux/_026_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_178_ ( .A(\req_msg[20] ), .X(\dpath/a_mux/_010_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_179_ ( .A(\dpath/a_mux/_096_ ), .X(\dpath/a_mux$out[4] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_180_ ( .A(\dpath/a_lt_b$in1[5] ), .X(\dpath/a_mux/_043_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_181_ ( .A(\resp_msg[5] ), .X(\dpath/a_mux/_027_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_182_ ( .A(\req_msg[21] ), .X(\dpath/a_mux/_011_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_183_ ( .A(\dpath/a_mux/_097_ ), .X(\dpath/a_mux$out[5] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_184_ ( .A(\dpath/a_lt_b$in1[6] ), .X(\dpath/a_mux/_044_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_185_ ( .A(\resp_msg[6] ), .X(\dpath/a_mux/_028_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_186_ ( .A(\req_msg[22] ), .X(\dpath/a_mux/_012_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_187_ ( .A(\dpath/a_mux/_098_ ), .X(\dpath/a_mux$out[6] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_188_ ( .A(\dpath/a_lt_b$in1[7] ), .X(\dpath/a_mux/_045_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_189_ ( .A(\resp_msg[7] ), .X(\dpath/a_mux/_029_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_190_ ( .A(\req_msg[23] ), .X(\dpath/a_mux/_013_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_191_ ( .A(\dpath/a_mux/_099_ ), .X(\dpath/a_mux$out[7] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_192_ ( .A(\dpath/a_lt_b$in1[8] ), .X(\dpath/a_mux/_046_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_193_ ( .A(\resp_msg[8] ), .X(\dpath/a_mux/_030_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_194_ ( .A(\req_msg[24] ), .X(\dpath/a_mux/_014_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_195_ ( .A(\dpath/a_mux/_100_ ), .X(\dpath/a_mux$out[8] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_196_ ( .A(\dpath/a_lt_b$in1[9] ), .X(\dpath/a_mux/_047_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_197_ ( .A(\resp_msg[9] ), .X(\dpath/a_mux/_031_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_198_ ( .A(\req_msg[25] ), .X(\dpath/a_mux/_015_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_199_ ( .A(\dpath/a_mux/_101_ ), .X(\dpath/a_mux$out[9] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_200_ ( .A(\dpath/a_lt_b$in1[10] ), .X(\dpath/a_mux/_033_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_201_ ( .A(\resp_msg[10] ), .X(\dpath/a_mux/_017_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_202_ ( .A(\req_msg[26] ), .X(\dpath/a_mux/_001_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_203_ ( .A(\dpath/a_mux/_087_ ), .X(\dpath/a_mux$out[10] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_204_ ( .A(\dpath/a_lt_b$in1[11] ), .X(\dpath/a_mux/_034_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_205_ ( .A(\resp_msg[11] ), .X(\dpath/a_mux/_018_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_206_ ( .A(\req_msg[27] ), .X(\dpath/a_mux/_002_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_207_ ( .A(\dpath/a_mux/_088_ ), .X(\dpath/a_mux$out[11] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_208_ ( .A(\dpath/a_lt_b$in1[12] ), .X(\dpath/a_mux/_035_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_209_ ( .A(\resp_msg[12] ), .X(\dpath/a_mux/_019_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_210_ ( .A(\req_msg[28] ), .X(\dpath/a_mux/_003_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_211_ ( .A(\dpath/a_mux/_089_ ), .X(\dpath/a_mux$out[12] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_212_ ( .A(\dpath/a_lt_b$in1[13] ), .X(\dpath/a_mux/_036_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_213_ ( .A(\resp_msg[13] ), .X(\dpath/a_mux/_020_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_214_ ( .A(\req_msg[29] ), .X(\dpath/a_mux/_004_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_215_ ( .A(\dpath/a_mux/_090_ ), .X(\dpath/a_mux$out[13] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_216_ ( .A(\dpath/a_lt_b$in1[14] ), .X(\dpath/a_mux/_037_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_217_ ( .A(\resp_msg[14] ), .X(\dpath/a_mux/_021_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_218_ ( .A(\req_msg[30] ), .X(\dpath/a_mux/_005_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_219_ ( .A(\dpath/a_mux/_091_ ), .X(\dpath/a_mux$out[14] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_220_ ( .A(\dpath/a_lt_b$in1[15] ), .X(\dpath/a_mux/_038_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_221_ ( .A(\resp_msg[15] ), .X(\dpath/a_mux/_022_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_222_ ( .A(\req_msg[31] ), .X(\dpath/a_mux/_006_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_223_ ( .A(\dpath/a_mux/_092_ ), .X(\dpath/a_mux$out[15] ) );
sky130_fd_sc_hs__buf_16 \dpath/a_reg/_066_ ( .A(\dpath/a_reg/_032_ ), .X(\dpath/a_reg/_049_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_067_ ( .A0(\dpath/a_reg/_050_ ), .A1(\dpath/a_reg/_033_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_016_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_068_ ( .A0(\dpath/a_reg/_057_ ), .A1(\dpath/a_reg/_040_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_023_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_069_ ( .A0(\dpath/a_reg/_058_ ), .A1(\dpath/a_reg/_041_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_024_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_070_ ( .A0(\dpath/a_reg/_059_ ), .A1(\dpath/a_reg/_042_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_025_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_071_ ( .A0(\dpath/a_reg/_060_ ), .A1(\dpath/a_reg/_043_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_026_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_072_ ( .A0(\dpath/a_reg/_061_ ), .A1(\dpath/a_reg/_044_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_027_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_073_ ( .A0(\dpath/a_reg/_062_ ), .A1(\dpath/a_reg/_045_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_028_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_074_ ( .A0(\dpath/a_reg/_063_ ), .A1(\dpath/a_reg/_046_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_029_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_075_ ( .A0(\dpath/a_reg/_064_ ), .A1(\dpath/a_reg/_047_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_030_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_076_ ( .A0(\dpath/a_reg/_065_ ), .A1(\dpath/a_reg/_048_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_031_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_077_ ( .A0(\dpath/a_reg/_051_ ), .A1(\dpath/a_reg/_034_ ), .S(\dpath/a_reg/_032_ ), .X(\dpath/a_reg/_017_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_078_ ( .A0(\dpath/a_reg/_052_ ), .A1(\dpath/a_reg/_035_ ), .S(\dpath/a_reg/_032_ ), .X(\dpath/a_reg/_018_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_079_ ( .A0(\dpath/a_reg/_053_ ), .A1(\dpath/a_reg/_036_ ), .S(\dpath/a_reg/_032_ ), .X(\dpath/a_reg/_019_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_080_ ( .A0(\dpath/a_reg/_054_ ), .A1(\dpath/a_reg/_037_ ), .S(\dpath/a_reg/_032_ ), .X(\dpath/a_reg/_020_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_081_ ( .A0(\dpath/a_reg/_055_ ), .A1(\dpath/a_reg/_038_ ), .S(\dpath/a_reg/_032_ ), .X(\dpath/a_reg/_021_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_082_ ( .A0(\dpath/a_reg/_056_ ), .A1(\dpath/a_reg/_039_ ), .S(\dpath/a_reg/_032_ ), .X(\dpath/a_reg/_022_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_083_ ( .A(\dpath/a_lt_b$in0[0] ), .X(\dpath/a_reg/_050_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_084_ ( .A(\dpath/a_mux$out[0] ), .X(\dpath/a_reg/_033_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_085_ ( .A(ctrl$a_reg_en ), .X(\dpath/a_reg/_032_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_086_ ( .A(\dpath/a_reg/_016_ ), .X(\dpath/a_reg/_000_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_087_ ( .A(\dpath/a_lt_b$in0[1] ), .X(\dpath/a_reg/_057_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_088_ ( .A(\dpath/a_mux$out[1] ), .X(\dpath/a_reg/_040_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_089_ ( .A(\dpath/a_reg/_023_ ), .X(\dpath/a_reg/_007_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_090_ ( .A(\dpath/a_lt_b$in0[2] ), .X(\dpath/a_reg/_058_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_091_ ( .A(\dpath/a_mux$out[2] ), .X(\dpath/a_reg/_041_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_092_ ( .A(\dpath/a_reg/_024_ ), .X(\dpath/a_reg/_008_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_093_ ( .A(\dpath/a_lt_b$in0[3] ), .X(\dpath/a_reg/_059_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_094_ ( .A(\dpath/a_mux$out[3] ), .X(\dpath/a_reg/_042_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_095_ ( .A(\dpath/a_reg/_025_ ), .X(\dpath/a_reg/_009_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_096_ ( .A(\dpath/a_lt_b$in0[4] ), .X(\dpath/a_reg/_060_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_097_ ( .A(\dpath/a_mux$out[4] ), .X(\dpath/a_reg/_043_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_098_ ( .A(\dpath/a_reg/_026_ ), .X(\dpath/a_reg/_010_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_099_ ( .A(\dpath/a_lt_b$in0[5] ), .X(\dpath/a_reg/_061_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_100_ ( .A(\dpath/a_mux$out[5] ), .X(\dpath/a_reg/_044_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_101_ ( .A(\dpath/a_reg/_027_ ), .X(\dpath/a_reg/_011_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_102_ ( .A(\dpath/a_lt_b$in0[6] ), .X(\dpath/a_reg/_062_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_103_ ( .A(\dpath/a_mux$out[6] ), .X(\dpath/a_reg/_045_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_104_ ( .A(\dpath/a_reg/_028_ ), .X(\dpath/a_reg/_012_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_105_ ( .A(\dpath/a_lt_b$in0[7] ), .X(\dpath/a_reg/_063_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_106_ ( .A(\dpath/a_mux$out[7] ), .X(\dpath/a_reg/_046_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_107_ ( .A(\dpath/a_reg/_029_ ), .X(\dpath/a_reg/_013_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_108_ ( .A(\dpath/a_lt_b$in0[8] ), .X(\dpath/a_reg/_064_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_109_ ( .A(\dpath/a_mux$out[8] ), .X(\dpath/a_reg/_047_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_110_ ( .A(\dpath/a_reg/_030_ ), .X(\dpath/a_reg/_014_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_111_ ( .A(\dpath/a_lt_b$in0[9] ), .X(\dpath/a_reg/_065_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_112_ ( .A(\dpath/a_mux$out[9] ), .X(\dpath/a_reg/_048_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_113_ ( .A(\dpath/a_reg/_031_ ), .X(\dpath/a_reg/_015_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_114_ ( .A(\dpath/a_lt_b$in0[10] ), .X(\dpath/a_reg/_051_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_115_ ( .A(\dpath/a_mux$out[10] ), .X(\dpath/a_reg/_034_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_116_ ( .A(\dpath/a_reg/_017_ ), .X(\dpath/a_reg/_001_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_117_ ( .A(\dpath/a_lt_b$in0[11] ), .X(\dpath/a_reg/_052_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_118_ ( .A(\dpath/a_mux$out[11] ), .X(\dpath/a_reg/_035_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_119_ ( .A(\dpath/a_reg/_018_ ), .X(\dpath/a_reg/_002_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_120_ ( .A(\dpath/a_lt_b$in0[12] ), .X(\dpath/a_reg/_053_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_121_ ( .A(\dpath/a_mux$out[12] ), .X(\dpath/a_reg/_036_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_122_ ( .A(\dpath/a_reg/_019_ ), .X(\dpath/a_reg/_003_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_123_ ( .A(\dpath/a_lt_b$in0[13] ), .X(\dpath/a_reg/_054_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_124_ ( .A(\dpath/a_mux$out[13] ), .X(\dpath/a_reg/_037_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_125_ ( .A(\dpath/a_reg/_020_ ), .X(\dpath/a_reg/_004_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_126_ ( .A(\dpath/a_lt_b$in0[14] ), .X(\dpath/a_reg/_055_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_127_ ( .A(\dpath/a_mux$out[14] ), .X(\dpath/a_reg/_038_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_128_ ( .A(\dpath/a_reg/_021_ ), .X(\dpath/a_reg/_005_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_129_ ( .A(\dpath/a_lt_b$in0[15] ), .X(\dpath/a_reg/_056_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_130_ ( .A(\dpath/a_mux$out[15] ), .X(\dpath/a_reg/_039_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_131_ ( .A(\dpath/a_reg/_022_ ), .X(\dpath/a_reg/_006_ ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_132_ ( .D(\dpath/a_reg/_000_ ), .Q(\dpath/a_lt_b$in0[0] ), .CLK(clk_66 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_133_ ( .D(\dpath/a_reg/_007_ ), .Q(\dpath/a_lt_b$in0[1] ), .CLK(clk_64 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_134_ ( .D(\dpath/a_reg/_008_ ), .Q(\dpath/a_lt_b$in0[2] ), .CLK(clk_63 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_135_ ( .D(\dpath/a_reg/_009_ ), .Q(\dpath/a_lt_b$in0[3] ), .CLK(clk_63 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_136_ ( .D(\dpath/a_reg/_010_ ), .Q(\dpath/a_lt_b$in0[4] ), .CLK(clk_86 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_137_ ( .D(\dpath/a_reg/_011_ ), .Q(\dpath/a_lt_b$in0[5] ), .CLK(clk_86 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_138_ ( .D(\dpath/a_reg/_012_ ), .Q(\dpath/a_lt_b$in0[6] ), .CLK(clk_70 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_139_ ( .D(\dpath/a_reg/_013_ ), .Q(\dpath/a_lt_b$in0[7] ), .CLK(clk_68 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_140_ ( .D(\dpath/a_reg/_014_ ), .Q(\dpath/a_lt_b$in0[8] ), .CLK(clk_69 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_141_ ( .D(\dpath/a_reg/_015_ ), .Q(\dpath/a_lt_b$in0[9] ), .CLK(clk_74 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_142_ ( .D(\dpath/a_reg/_001_ ), .Q(\dpath/a_lt_b$in0[10] ), .CLK(clk_76 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_143_ ( .D(\dpath/a_reg/_002_ ), .Q(\dpath/a_lt_b$in0[11] ), .CLK(clk_78 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_144_ ( .D(\dpath/a_reg/_003_ ), .Q(\dpath/a_lt_b$in0[12] ), .CLK(clk_80 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_145_ ( .D(\dpath/a_reg/_004_ ), .Q(\dpath/a_lt_b$in0[13] ), .CLK(clk_79 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_146_ ( .D(\dpath/a_reg/_005_ ), .Q(\dpath/a_lt_b$in0[14] ), .CLK(clk_58 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_147_ ( .D(\dpath/a_reg/_006_ ), .Q(\dpath/a_lt_b$in0[15] ), .CLK(clk_82 ) );
sky130_fd_sc_hs__buf_16 \dpath/b_mux/_050_ ( .A(\dpath/b_mux/_049_ ), .X(\dpath/b_mux/_032_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_051_ ( .A0(\dpath/b_mux/_000_ ), .A1(\dpath/b_mux/_016_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_033_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_052_ ( .A0(\dpath/b_mux/_007_ ), .A1(\dpath/b_mux/_023_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_040_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_053_ ( .A0(\dpath/b_mux/_008_ ), .A1(\dpath/b_mux/_024_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_041_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_054_ ( .A0(\dpath/b_mux/_009_ ), .A1(\dpath/b_mux/_025_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_042_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_055_ ( .A0(\dpath/b_mux/_010_ ), .A1(\dpath/b_mux/_026_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_043_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_056_ ( .A0(\dpath/b_mux/_011_ ), .A1(\dpath/b_mux/_027_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_044_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_057_ ( .A0(\dpath/b_mux/_012_ ), .A1(\dpath/b_mux/_028_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_045_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_058_ ( .A0(\dpath/b_mux/_013_ ), .A1(\dpath/b_mux/_029_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_046_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_059_ ( .A0(\dpath/b_mux/_014_ ), .A1(\dpath/b_mux/_030_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_047_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_060_ ( .A0(\dpath/b_mux/_015_ ), .A1(\dpath/b_mux/_031_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_048_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_061_ ( .A0(\dpath/b_mux/_001_ ), .A1(\dpath/b_mux/_017_ ), .S(\dpath/b_mux/_049_ ), .X(\dpath/b_mux/_034_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_062_ ( .A0(\dpath/b_mux/_002_ ), .A1(\dpath/b_mux/_018_ ), .S(\dpath/b_mux/_049_ ), .X(\dpath/b_mux/_035_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_063_ ( .A0(\dpath/b_mux/_003_ ), .A1(\dpath/b_mux/_019_ ), .S(\dpath/b_mux/_049_ ), .X(\dpath/b_mux/_036_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_064_ ( .A0(\dpath/b_mux/_004_ ), .A1(\dpath/b_mux/_020_ ), .S(\dpath/b_mux/_049_ ), .X(\dpath/b_mux/_037_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_065_ ( .A0(\dpath/b_mux/_005_ ), .A1(\dpath/b_mux/_021_ ), .S(\dpath/b_mux/_049_ ), .X(\dpath/b_mux/_038_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_066_ ( .A0(\dpath/b_mux/_006_ ), .A1(\dpath/b_mux/_022_ ), .S(\dpath/b_mux/_049_ ), .X(\dpath/b_mux/_039_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_067_ ( .A(\dpath/a_lt_b$in0[0] ), .X(\dpath/b_mux/_000_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_068_ ( .A(\req_msg[0] ), .X(\dpath/b_mux/_016_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_069_ ( .A(ctrl$b_mux_sel ), .X(\dpath/b_mux/_049_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_070_ ( .A(\dpath/b_mux/_033_ ), .X(\dpath/b_mux$out[0] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_071_ ( .A(\dpath/a_lt_b$in0[1] ), .X(\dpath/b_mux/_007_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_072_ ( .A(\req_msg[1] ), .X(\dpath/b_mux/_023_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_073_ ( .A(\dpath/b_mux/_040_ ), .X(\dpath/b_mux$out[1] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_074_ ( .A(\dpath/a_lt_b$in0[2] ), .X(\dpath/b_mux/_008_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_075_ ( .A(\req_msg[2] ), .X(\dpath/b_mux/_024_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_076_ ( .A(\dpath/b_mux/_041_ ), .X(\dpath/b_mux$out[2] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_077_ ( .A(\dpath/a_lt_b$in0[3] ), .X(\dpath/b_mux/_009_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_078_ ( .A(\req_msg[3] ), .X(\dpath/b_mux/_025_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_079_ ( .A(\dpath/b_mux/_042_ ), .X(\dpath/b_mux$out[3] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_080_ ( .A(\dpath/a_lt_b$in0[4] ), .X(\dpath/b_mux/_010_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_081_ ( .A(\req_msg[4] ), .X(\dpath/b_mux/_026_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_082_ ( .A(\dpath/b_mux/_043_ ), .X(\dpath/b_mux$out[4] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_083_ ( .A(\dpath/a_lt_b$in0[5] ), .X(\dpath/b_mux/_011_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_084_ ( .A(\req_msg[5] ), .X(\dpath/b_mux/_027_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_085_ ( .A(\dpath/b_mux/_044_ ), .X(\dpath/b_mux$out[5] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_086_ ( .A(\dpath/a_lt_b$in0[6] ), .X(\dpath/b_mux/_012_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_087_ ( .A(\req_msg[6] ), .X(\dpath/b_mux/_028_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_088_ ( .A(\dpath/b_mux/_045_ ), .X(\dpath/b_mux$out[6] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_089_ ( .A(\dpath/a_lt_b$in0[7] ), .X(\dpath/b_mux/_013_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_090_ ( .A(\req_msg[7] ), .X(\dpath/b_mux/_029_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_091_ ( .A(\dpath/b_mux/_046_ ), .X(\dpath/b_mux$out[7] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_092_ ( .A(\dpath/a_lt_b$in0[8] ), .X(\dpath/b_mux/_014_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_093_ ( .A(\req_msg[8] ), .X(\dpath/b_mux/_030_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_094_ ( .A(\dpath/b_mux/_047_ ), .X(\dpath/b_mux$out[8] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_095_ ( .A(\dpath/a_lt_b$in0[9] ), .X(\dpath/b_mux/_015_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_096_ ( .A(\req_msg[9] ), .X(\dpath/b_mux/_031_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_097_ ( .A(\dpath/b_mux/_048_ ), .X(\dpath/b_mux$out[9] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_098_ ( .A(\dpath/a_lt_b$in0[10] ), .X(\dpath/b_mux/_001_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_099_ ( .A(\req_msg[10] ), .X(\dpath/b_mux/_017_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_100_ ( .A(\dpath/b_mux/_034_ ), .X(\dpath/b_mux$out[10] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_101_ ( .A(\dpath/a_lt_b$in0[11] ), .X(\dpath/b_mux/_002_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_102_ ( .A(\req_msg[11] ), .X(\dpath/b_mux/_018_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_103_ ( .A(\dpath/b_mux/_035_ ), .X(\dpath/b_mux$out[11] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_104_ ( .A(\dpath/a_lt_b$in0[12] ), .X(\dpath/b_mux/_003_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_105_ ( .A(\req_msg[12] ), .X(\dpath/b_mux/_019_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_106_ ( .A(\dpath/b_mux/_036_ ), .X(\dpath/b_mux$out[12] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_107_ ( .A(\dpath/a_lt_b$in0[13] ), .X(\dpath/b_mux/_004_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_108_ ( .A(\req_msg[13] ), .X(\dpath/b_mux/_020_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_109_ ( .A(\dpath/b_mux/_037_ ), .X(\dpath/b_mux$out[13] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_110_ ( .A(\dpath/a_lt_b$in0[14] ), .X(\dpath/b_mux/_005_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_111_ ( .A(\req_msg[14] ), .X(\dpath/b_mux/_021_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_112_ ( .A(\dpath/b_mux/_038_ ), .X(\dpath/b_mux$out[14] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_113_ ( .A(\dpath/a_lt_b$in0[15] ), .X(\dpath/b_mux/_006_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_114_ ( .A(\req_msg[15] ), .X(\dpath/b_mux/_022_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_115_ ( .A(\dpath/b_mux/_039_ ), .X(\dpath/b_mux$out[15] ) );
sky130_fd_sc_hs__buf_16 \dpath/b_reg/_066_ ( .A(\dpath/b_reg/_032_ ), .X(\dpath/b_reg/_049_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_067_ ( .A0(\dpath/b_reg/_050_ ), .A1(\dpath/b_reg/_033_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_016_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_068_ ( .A0(\dpath/b_reg/_057_ ), .A1(\dpath/b_reg/_040_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_023_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_069_ ( .A0(\dpath/b_reg/_058_ ), .A1(\dpath/b_reg/_041_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_024_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_070_ ( .A0(\dpath/b_reg/_059_ ), .A1(\dpath/b_reg/_042_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_025_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_071_ ( .A0(\dpath/b_reg/_060_ ), .A1(\dpath/b_reg/_043_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_026_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_072_ ( .A0(\dpath/b_reg/_061_ ), .A1(\dpath/b_reg/_044_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_027_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_073_ ( .A0(\dpath/b_reg/_062_ ), .A1(\dpath/b_reg/_045_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_028_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_074_ ( .A0(\dpath/b_reg/_063_ ), .A1(\dpath/b_reg/_046_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_029_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_075_ ( .A0(\dpath/b_reg/_064_ ), .A1(\dpath/b_reg/_047_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_030_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_076_ ( .A0(\dpath/b_reg/_065_ ), .A1(\dpath/b_reg/_048_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_031_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_077_ ( .A0(\dpath/b_reg/_051_ ), .A1(\dpath/b_reg/_034_ ), .S(\dpath/b_reg/_032_ ), .X(\dpath/b_reg/_017_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_078_ ( .A0(\dpath/b_reg/_052_ ), .A1(\dpath/b_reg/_035_ ), .S(\dpath/b_reg/_032_ ), .X(\dpath/b_reg/_018_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_079_ ( .A0(\dpath/b_reg/_053_ ), .A1(\dpath/b_reg/_036_ ), .S(\dpath/b_reg/_032_ ), .X(\dpath/b_reg/_019_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_080_ ( .A0(\dpath/b_reg/_054_ ), .A1(\dpath/b_reg/_037_ ), .S(\dpath/b_reg/_032_ ), .X(\dpath/b_reg/_020_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_081_ ( .A0(\dpath/b_reg/_055_ ), .A1(\dpath/b_reg/_038_ ), .S(\dpath/b_reg/_032_ ), .X(\dpath/b_reg/_021_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_082_ ( .A0(\dpath/b_reg/_056_ ), .A1(\dpath/b_reg/_039_ ), .S(\dpath/b_reg/_032_ ), .X(\dpath/b_reg/_022_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_083_ ( .A(\dpath/a_lt_b$in1[0] ), .X(\dpath/b_reg/_050_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_084_ ( .A(\dpath/b_mux$out[0] ), .X(\dpath/b_reg/_033_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_085_ ( .A(ctrl$b_reg_en ), .X(\dpath/b_reg/_032_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_086_ ( .A(\dpath/b_reg/_016_ ), .X(\dpath/b_reg/_000_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_087_ ( .A(\dpath/a_lt_b$in1[1] ), .X(\dpath/b_reg/_057_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_088_ ( .A(\dpath/b_mux$out[1] ), .X(\dpath/b_reg/_040_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_089_ ( .A(\dpath/b_reg/_023_ ), .X(\dpath/b_reg/_007_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_090_ ( .A(\dpath/a_lt_b$in1[2] ), .X(\dpath/b_reg/_058_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_091_ ( .A(\dpath/b_mux$out[2] ), .X(\dpath/b_reg/_041_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_092_ ( .A(\dpath/b_reg/_024_ ), .X(\dpath/b_reg/_008_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_093_ ( .A(\dpath/a_lt_b$in1[3] ), .X(\dpath/b_reg/_059_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_094_ ( .A(\dpath/b_mux$out[3] ), .X(\dpath/b_reg/_042_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_095_ ( .A(\dpath/b_reg/_025_ ), .X(\dpath/b_reg/_009_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_096_ ( .A(\dpath/a_lt_b$in1[4] ), .X(\dpath/b_reg/_060_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_097_ ( .A(\dpath/b_mux$out[4] ), .X(\dpath/b_reg/_043_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_098_ ( .A(\dpath/b_reg/_026_ ), .X(\dpath/b_reg/_010_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_099_ ( .A(\dpath/a_lt_b$in1[5] ), .X(\dpath/b_reg/_061_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_100_ ( .A(\dpath/b_mux$out[5] ), .X(\dpath/b_reg/_044_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_101_ ( .A(\dpath/b_reg/_027_ ), .X(\dpath/b_reg/_011_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_102_ ( .A(\dpath/a_lt_b$in1[6] ), .X(\dpath/b_reg/_062_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_103_ ( .A(\dpath/b_mux$out[6] ), .X(\dpath/b_reg/_045_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_104_ ( .A(\dpath/b_reg/_028_ ), .X(\dpath/b_reg/_012_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_105_ ( .A(\dpath/a_lt_b$in1[7] ), .X(\dpath/b_reg/_063_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_106_ ( .A(\dpath/b_mux$out[7] ), .X(\dpath/b_reg/_046_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_107_ ( .A(\dpath/b_reg/_029_ ), .X(\dpath/b_reg/_013_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_108_ ( .A(\dpath/a_lt_b$in1[8] ), .X(\dpath/b_reg/_064_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_109_ ( .A(\dpath/b_mux$out[8] ), .X(\dpath/b_reg/_047_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_110_ ( .A(\dpath/b_reg/_030_ ), .X(\dpath/b_reg/_014_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_111_ ( .A(\dpath/a_lt_b$in1[9] ), .X(\dpath/b_reg/_065_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_112_ ( .A(\dpath/b_mux$out[9] ), .X(\dpath/b_reg/_048_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_113_ ( .A(\dpath/b_reg/_031_ ), .X(\dpath/b_reg/_015_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_114_ ( .A(\dpath/a_lt_b$in1[10] ), .X(\dpath/b_reg/_051_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_115_ ( .A(\dpath/b_mux$out[10] ), .X(\dpath/b_reg/_034_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_116_ ( .A(\dpath/b_reg/_017_ ), .X(\dpath/b_reg/_001_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_117_ ( .A(\dpath/a_lt_b$in1[11] ), .X(\dpath/b_reg/_052_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_118_ ( .A(\dpath/b_mux$out[11] ), .X(\dpath/b_reg/_035_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_119_ ( .A(\dpath/b_reg/_018_ ), .X(\dpath/b_reg/_002_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_120_ ( .A(\dpath/a_lt_b$in1[12] ), .X(\dpath/b_reg/_053_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_121_ ( .A(\dpath/b_mux$out[12] ), .X(\dpath/b_reg/_036_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_122_ ( .A(\dpath/b_reg/_019_ ), .X(\dpath/b_reg/_003_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_123_ ( .A(\dpath/a_lt_b$in1[13] ), .X(\dpath/b_reg/_054_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_124_ ( .A(\dpath/b_mux$out[13] ), .X(\dpath/b_reg/_037_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_125_ ( .A(\dpath/b_reg/_020_ ), .X(\dpath/b_reg/_004_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_126_ ( .A(\dpath/a_lt_b$in1[14] ), .X(\dpath/b_reg/_055_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_127_ ( .A(\dpath/b_mux$out[14] ), .X(\dpath/b_reg/_038_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_128_ ( .A(\dpath/b_reg/_021_ ), .X(\dpath/b_reg/_005_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_129_ ( .A(\dpath/a_lt_b$in1[15] ), .X(\dpath/b_reg/_056_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_130_ ( .A(\dpath/b_mux$out[15] ), .X(\dpath/b_reg/_039_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_131_ ( .A(\dpath/b_reg/_022_ ), .X(\dpath/b_reg/_006_ ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_132_ ( .D(\dpath/b_reg/_000_ ), .Q(\dpath/a_lt_b$in1[0] ), .CLK(clk_67 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_133_ ( .D(\dpath/b_reg/_007_ ), .Q(\dpath/a_lt_b$in1[1] ), .CLK(clk_65 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_134_ ( .D(\dpath/b_reg/_008_ ), .Q(\dpath/a_lt_b$in1[2] ), .CLK(clk_62 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_135_ ( .D(\dpath/b_reg/_009_ ), .Q(\dpath/a_lt_b$in1[3] ), .CLK(clk_62 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_136_ ( .D(\dpath/b_reg/_010_ ), .Q(\dpath/a_lt_b$in1[4] ), .CLK(clk_72 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_137_ ( .D(\dpath/b_reg/_011_ ), .Q(\dpath/a_lt_b$in1[5] ), .CLK(clk_73 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_138_ ( .D(\dpath/b_reg/_012_ ), .Q(\dpath/a_lt_b$in1[6] ), .CLK(clk_75 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_139_ ( .D(\dpath/b_reg/_013_ ), .Q(\dpath/a_lt_b$in1[7] ), .CLK(clk_71 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_140_ ( .D(\dpath/b_reg/_014_ ), .Q(\dpath/a_lt_b$in1[8] ), .CLK(clk_77 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_141_ ( .D(\dpath/b_reg/_015_ ), .Q(\dpath/a_lt_b$in1[9] ), .CLK(clk_77 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_142_ ( .D(\dpath/b_reg/_001_ ), .Q(\dpath/a_lt_b$in1[10] ), .CLK(clk_76 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_143_ ( .D(\dpath/b_reg/_002_ ), .Q(\dpath/a_lt_b$in1[11] ), .CLK(clk_83 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_144_ ( .D(\dpath/b_reg/_003_ ), .Q(\dpath/a_lt_b$in1[12] ), .CLK(clk_84 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_145_ ( .D(\dpath/b_reg/_004_ ), .Q(\dpath/a_lt_b$in1[13] ), .CLK(clk_57 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_146_ ( .D(\dpath/b_reg/_005_ ), .Q(\dpath/a_lt_b$in1[14] ), .CLK(clk_81 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_147_ ( .D(\dpath/b_reg/_006_ ), .Q(\dpath/a_lt_b$in1[15] ), .CLK(clk_58 ) );
sky130_fd_sc_hs__nor2_2 \dpath/b_zero/_25_ ( .A(\dpath/b_zero/_10_ ), .B(\dpath/b_zero/_13_ ), .Y(\dpath/b_zero/_16_ ) );
sky130_fd_sc_hs__nor3b_1 \dpath/b_zero/_26_ ( .A(\dpath/b_zero/_07_ ), .B(\dpath/b_zero/_08_ ), .C_N(\dpath/b_zero/_16_ ), .Y(\dpath/b_zero/_17_ ) );
sky130_fd_sc_hs__nor2_4 \dpath/b_zero/_27_ ( .A(\dpath/b_zero/_04_ ), .B(\dpath/b_zero/_05_ ), .Y(\dpath/b_zero/_18_ ) );
sky130_fd_sc_hs__nor3b_1 \dpath/b_zero/_28_ ( .A(\dpath/b_zero/_14_ ), .B(\dpath/b_zero/_02_ ), .C_N(\dpath/b_zero/_18_ ), .Y(\dpath/b_zero/_19_ ) );
sky130_fd_sc_hs__nor2_1 \dpath/b_zero/_29_ ( .A(\dpath/b_zero/_00_ ), .B(\dpath/b_zero/_09_ ), .Y(\dpath/b_zero/_20_ ) );
sky130_fd_sc_hs__nor3b_2 \dpath/b_zero/_30_ ( .A(\dpath/b_zero/_11_ ), .B(\dpath/b_zero/_12_ ), .C_N(\dpath/b_zero/_20_ ), .Y(\dpath/b_zero/_21_ ) );
sky130_fd_sc_hs__nor2_1 \dpath/b_zero/_31_ ( .A(\dpath/b_zero/_03_ ), .B(\dpath/b_zero/_06_ ), .Y(\dpath/b_zero/_22_ ) );
sky130_fd_sc_hs__nor3b_2 \dpath/b_zero/_32_ ( .A(\dpath/b_zero/_15_ ), .B(\dpath/b_zero/_01_ ), .C_N(\dpath/b_zero/_22_ ), .Y(\dpath/b_zero/_23_ ) );
sky130_fd_sc_hs__and4_1 \dpath/b_zero/_33_ ( .A(\dpath/b_zero/_17_ ), .B(\dpath/b_zero/_19_ ), .C(\dpath/b_zero/_21_ ), .D(\dpath/b_zero/_23_ ), .X(\dpath/b_zero/_24_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_34_ ( .A(\dpath/a_lt_b$in1[1] ), .X(\dpath/b_zero/_07_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_35_ ( .A(\dpath/a_lt_b$in1[0] ), .X(\dpath/b_zero/_00_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_36_ ( .A(\dpath/a_lt_b$in1[3] ), .X(\dpath/b_zero/_09_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_37_ ( .A(\dpath/a_lt_b$in1[2] ), .X(\dpath/b_zero/_08_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_38_ ( .A(\dpath/a_lt_b$in1[5] ), .X(\dpath/b_zero/_11_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_39_ ( .A(\dpath/a_lt_b$in1[4] ), .X(\dpath/b_zero/_10_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_40_ ( .A(\dpath/a_lt_b$in1[7] ), .X(\dpath/b_zero/_13_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_41_ ( .A(\dpath/a_lt_b$in1[6] ), .X(\dpath/b_zero/_12_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_42_ ( .A(\dpath/a_lt_b$in1[9] ), .X(\dpath/b_zero/_15_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_43_ ( .A(\dpath/a_lt_b$in1[8] ), .X(\dpath/b_zero/_14_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_44_ ( .A(\dpath/a_lt_b$in1[11] ), .X(\dpath/b_zero/_02_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_45_ ( .A(\dpath/a_lt_b$in1[10] ), .X(\dpath/b_zero/_01_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_46_ ( .A(\dpath/a_lt_b$in1[13] ), .X(\dpath/b_zero/_04_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_47_ ( .A(\dpath/a_lt_b$in1[12] ), .X(\dpath/b_zero/_03_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_48_ ( .A(\dpath/a_lt_b$in1[15] ), .X(\dpath/b_zero/_06_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_49_ ( .A(\dpath/a_lt_b$in1[14] ), .X(\dpath/b_zero/_05_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_50_ ( .A(\dpath/b_zero/_24_ ), .X(ctrl$is_b_zero ) );
sky130_fd_sc_hs__xor2_1 \dpath/sub/_121_ ( .A(\dpath/sub/_000_ ), .B(\dpath/sub/_016_ ), .X(\dpath/sub/_105_ ) );
sky130_fd_sc_hs__nand2b_4 \dpath/sub/_122_ ( .A_N(\dpath/sub/_000_ ), .B(\dpath/sub/_016_ ), .Y(\dpath/sub/_063_ ) );
sky130_fd_sc_hs__xnor3_4 \dpath/sub/_123_ ( .A(\dpath/sub/_007_ ), .B(\dpath/sub/_023_ ), .C(\dpath/sub/_063_ ), .X(\dpath/sub/_112_ ) );
sky130_fd_sc_hs__nand2b_4 \dpath/sub/_124_ ( .A_N(\dpath/sub/_023_ ), .B(\dpath/sub/_007_ ), .Y(\dpath/sub/_064_ ) );
sky130_fd_sc_hs__nand2b_4 \dpath/sub/_125_ ( .A_N(\dpath/sub/_007_ ), .B(\dpath/sub/_023_ ), .Y(\dpath/sub/_065_ ) );
sky130_fd_sc_hs__nand3_2 \dpath/sub/_126_ ( .A(\dpath/sub/_063_ ), .B(\dpath/sub/_064_ ), .C(\dpath/sub/_065_ ), .Y(\dpath/sub/_066_ ) );
sky130_fd_sc_hs__nand2_2 \dpath/sub/_127_ ( .A(\dpath/sub/_066_ ), .B(\dpath/sub/_064_ ), .Y(\dpath/sub/_067_ ) );
sky130_fd_sc_hs__xnor3_4 \dpath/sub/_128_ ( .A(\dpath/sub/_008_ ), .B(\dpath/sub/_024_ ), .C(\dpath/sub/_067_ ), .X(\dpath/sub/_113_ ) );
sky130_fd_sc_hs__xnor2_4 \dpath/sub/_129_ ( .A(\dpath/sub/_009_ ), .B(\dpath/sub/_025_ ), .Y(\dpath/sub/_068_ ) );
sky130_fd_sc_hs__and2b_4 \dpath/sub/_130_ ( .A_N(\dpath/sub/_024_ ), .B(\dpath/sub/_008_ ), .X(\dpath/sub/_069_ ) );
sky130_fd_sc_hs__xnor2_4 \dpath/sub/_131_ ( .A(\dpath/sub/_008_ ), .B(\dpath/sub/_024_ ), .Y(\dpath/sub/_070_ ) );
sky130_fd_sc_hs__a21boi_1 \dpath/sub/_132_ ( .A1(\dpath/sub/_066_ ), .A2(\dpath/sub/_064_ ), .B1_N(\dpath/sub/_070_ ), .Y(\dpath/sub/_071_ ) );
sky130_fd_sc_hs__nor2_1 \dpath/sub/_133_ ( .A(\dpath/sub/_069_ ), .B(\dpath/sub/_071_ ), .Y(\dpath/sub/_072_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_134_ ( .A(\dpath/sub/_068_ ), .B(\dpath/sub/_072_ ), .Y(\dpath/sub/_114_ ) );
sky130_fd_sc_hs__nand3_4 \dpath/sub/_135_ ( .A(\dpath/sub/_067_ ), .B(\dpath/sub/_070_ ), .C(\dpath/sub/_068_ ), .Y(\dpath/sub/_073_ ) );
sky130_fd_sc_hs__nor2b_2 \dpath/sub/_136_ ( .A(\dpath/sub/_025_ ), .B_N(\dpath/sub/_009_ ), .Y(\dpath/sub/_074_ ) );
sky130_fd_sc_hs__a21oi_2 \dpath/sub/_137_ ( .A1(\dpath/sub/_068_ ), .A2(\dpath/sub/_069_ ), .B1(\dpath/sub/_074_ ), .Y(\dpath/sub/_075_ ) );
sky130_fd_sc_hs__xnor2_2 \dpath/sub/_138_ ( .A(\dpath/sub/_010_ ), .B(\dpath/sub/_026_ ), .Y(\dpath/sub/_076_ ) );
sky130_fd_sc_hs__a21bo_1 \dpath/sub/_139_ ( .A1(\dpath/sub/_073_ ), .A2(\dpath/sub/_075_ ), .B1_N(\dpath/sub/_076_ ), .X(\dpath/sub/_077_ ) );
sky130_fd_sc_hs__nand3b_1 \dpath/sub/_140_ ( .A_N(\dpath/sub/_076_ ), .B(\dpath/sub/_073_ ), .C(\dpath/sub/_075_ ), .Y(\dpath/sub/_078_ ) );
sky130_fd_sc_hs__and2_1 \dpath/sub/_141_ ( .A(\dpath/sub/_077_ ), .B(\dpath/sub/_078_ ), .X(\dpath/sub/_115_ ) );
sky130_fd_sc_hs__xnor2_4 \dpath/sub/_142_ ( .A(\dpath/sub/_011_ ), .B(\dpath/sub/_027_ ), .Y(\dpath/sub/_079_ ) );
sky130_fd_sc_hs__nor2b_4 \dpath/sub/_143_ ( .A(\dpath/sub/_026_ ), .B_N(\dpath/sub/_010_ ), .Y(\dpath/sub/_080_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_144_ ( .A_N(\dpath/sub/_080_ ), .B(\dpath/sub/_077_ ), .X(\dpath/sub/_081_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_145_ ( .A(\dpath/sub/_079_ ), .B(\dpath/sub/_081_ ), .Y(\dpath/sub/_116_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_146_ ( .A_N(\dpath/sub/_027_ ), .B(\dpath/sub/_011_ ), .X(\dpath/sub/_082_ ) );
sky130_fd_sc_hs__a21oi_2 \dpath/sub/_147_ ( .A1(\dpath/sub/_079_ ), .A2(\dpath/sub/_080_ ), .B1(\dpath/sub/_082_ ), .Y(\dpath/sub/_083_ ) );
sky130_fd_sc_hs__inv_2 \dpath/sub/_148_ ( .A(\dpath/sub/_083_ ), .Y(\dpath/sub/_084_ ) );
sky130_fd_sc_hs__xnor2_4 \dpath/sub/_149_ ( .A(\dpath/sub/_012_ ), .B(\dpath/sub/_028_ ), .Y(\dpath/sub/_085_ ) );
sky130_fd_sc_hs__and2_1 \dpath/sub/_150_ ( .A(\dpath/sub/_076_ ), .B(\dpath/sub/_079_ ), .X(\dpath/sub/_086_ ) );
sky130_fd_sc_hs__a21boi_1 \dpath/sub/_151_ ( .A1(\dpath/sub/_073_ ), .A2(\dpath/sub/_075_ ), .B1_N(\dpath/sub/_086_ ), .Y(\dpath/sub/_087_ ) );
sky130_fd_sc_hs__or3_1 \dpath/sub/_152_ ( .A(\dpath/sub/_084_ ), .B(\dpath/sub/_085_ ), .C(\dpath/sub/_087_ ), .X(\dpath/sub/_088_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/sub/_153_ ( .A1(\dpath/sub/_084_ ), .A2(\dpath/sub/_087_ ), .B1(\dpath/sub/_085_ ), .Y(\dpath/sub/_089_ ) );
sky130_fd_sc_hs__and2_1 \dpath/sub/_154_ ( .A(\dpath/sub/_088_ ), .B(\dpath/sub/_089_ ), .X(\dpath/sub/_117_ ) );
sky130_fd_sc_hs__xnor2_2 \dpath/sub/_155_ ( .A(\dpath/sub/_013_ ), .B(\dpath/sub/_029_ ), .Y(\dpath/sub/_090_ ) );
sky130_fd_sc_hs__inv_1 \dpath/sub/_156_ ( .A(\dpath/sub/_090_ ), .Y(\dpath/sub/_091_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/sub/_157_ ( .A(\dpath/sub/_028_ ), .B_N(\dpath/sub/_012_ ), .X(\dpath/sub/_092_ ) );
sky130_fd_sc_hs__nand2_1 \dpath/sub/_158_ ( .A(\dpath/sub/_089_ ), .B(\dpath/sub/_092_ ), .Y(\dpath/sub/_093_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_159_ ( .A(\dpath/sub/_091_ ), .B(\dpath/sub/_093_ ), .Y(\dpath/sub/_118_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_160_ ( .A(\dpath/sub/_014_ ), .B(\dpath/sub/_030_ ), .Y(\dpath/sub/_094_ ) );
sky130_fd_sc_hs__and4_1 \dpath/sub/_161_ ( .A(\dpath/sub/_076_ ), .B(\dpath/sub/_079_ ), .C(\dpath/sub/_085_ ), .D(\dpath/sub/_090_ ), .X(\dpath/sub/_095_ ) );
sky130_fd_sc_hs__a21boi_4 \dpath/sub/_162_ ( .A1(\dpath/sub/_073_ ), .A2(\dpath/sub/_075_ ), .B1_N(\dpath/sub/_095_ ), .Y(\dpath/sub/_096_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_163_ ( .A_N(\dpath/sub/_029_ ), .B(\dpath/sub/_013_ ), .X(\dpath/sub/_097_ ) );
sky130_fd_sc_hs__o21bai_1 \dpath/sub/_164_ ( .A1(\dpath/sub/_092_ ), .A2(\dpath/sub/_091_ ), .B1_N(\dpath/sub/_097_ ), .Y(\dpath/sub/_098_ ) );
sky130_fd_sc_hs__a31oi_1 \dpath/sub/_165_ ( .A1(\dpath/sub/_084_ ), .A2(\dpath/sub/_085_ ), .A3(\dpath/sub/_090_ ), .B1(\dpath/sub/_098_ ), .Y(\dpath/sub/_099_ ) );
sky130_fd_sc_hs__nor2b_2 \dpath/sub/_166_ ( .A(\dpath/sub/_096_ ), .B_N(\dpath/sub/_099_ ), .Y(\dpath/sub/_100_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_167_ ( .A(\dpath/sub/_094_ ), .B(\dpath/sub/_100_ ), .Y(\dpath/sub/_119_ ) );
sky130_fd_sc_hs__xnor2_4 \dpath/sub/_168_ ( .A(\dpath/sub/_015_ ), .B(\dpath/sub/_031_ ), .Y(\dpath/sub/_101_ ) );
sky130_fd_sc_hs__nor2b_4 \dpath/sub/_169_ ( .A(\dpath/sub/_030_ ), .B_N(\dpath/sub/_014_ ), .Y(\dpath/sub/_102_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/sub/_170_ ( .A(\dpath/sub/_100_ ), .B_N(\dpath/sub/_094_ ), .X(\dpath/sub/_103_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_171_ ( .A_N(\dpath/sub/_102_ ), .B(\dpath/sub/_103_ ), .X(\dpath/sub/_104_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_172_ ( .A(\dpath/sub/_101_ ), .B(\dpath/sub/_104_ ), .Y(\dpath/sub/_120_ ) );
sky130_fd_sc_hs__nand3b_1 \dpath/sub/_173_ ( .A_N(\dpath/sub/_100_ ), .B(\dpath/sub/_094_ ), .C(\dpath/sub/_101_ ), .Y(\dpath/sub/_032_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_174_ ( .A_N(\dpath/sub/_031_ ), .B(\dpath/sub/_015_ ), .X(\dpath/sub/_033_ ) );
sky130_fd_sc_hs__a21oi_4 \dpath/sub/_175_ ( .A1(\dpath/sub/_101_ ), .A2(\dpath/sub/_102_ ), .B1(\dpath/sub/_033_ ), .Y(\dpath/sub/_034_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_176_ ( .A(\dpath/sub/_001_ ), .B(\dpath/sub/_017_ ), .Y(\dpath/sub/_035_ ) );
sky130_fd_sc_hs__inv_1 \dpath/sub/_177_ ( .A(\dpath/sub/_035_ ), .Y(\dpath/sub/_036_ ) );
sky130_fd_sc_hs__a21o_1 \dpath/sub/_178_ ( .A1(\dpath/sub/_032_ ), .A2(\dpath/sub/_034_ ), .B1(\dpath/sub/_036_ ), .X(\dpath/sub/_037_ ) );
sky130_fd_sc_hs__nand3_1 \dpath/sub/_179_ ( .A(\dpath/sub/_032_ ), .B(\dpath/sub/_034_ ), .C(\dpath/sub/_036_ ), .Y(\dpath/sub/_038_ ) );
sky130_fd_sc_hs__and2_1 \dpath/sub/_180_ ( .A(\dpath/sub/_037_ ), .B(\dpath/sub/_038_ ), .X(\dpath/sub/_106_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_181_ ( .A(\dpath/sub/_002_ ), .B(\dpath/sub/_018_ ), .Y(\dpath/sub/_039_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_182_ ( .A_N(\dpath/sub/_017_ ), .B(\dpath/sub/_001_ ), .X(\dpath/sub/_040_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_183_ ( .A_N(\dpath/sub/_040_ ), .B(\dpath/sub/_037_ ), .X(\dpath/sub/_041_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_184_ ( .A(\dpath/sub/_039_ ), .B(\dpath/sub/_041_ ), .Y(\dpath/sub/_107_ ) );
sky130_fd_sc_hs__and4_1 \dpath/sub/_185_ ( .A(\dpath/sub/_094_ ), .B(\dpath/sub/_101_ ), .C(\dpath/sub/_035_ ), .D(\dpath/sub/_039_ ), .X(\dpath/sub/_042_ ) );
sky130_fd_sc_hs__nand2b_2 \dpath/sub/_186_ ( .A_N(\dpath/sub/_100_ ), .B(\dpath/sub/_042_ ), .Y(\dpath/sub/_043_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_187_ ( .A_N(\dpath/sub/_018_ ), .B(\dpath/sub/_002_ ), .X(\dpath/sub/_044_ ) );
sky130_fd_sc_hs__nor3b_1 \dpath/sub/_188_ ( .A(\dpath/sub/_036_ ), .B(\dpath/sub/_034_ ), .C_N(\dpath/sub/_039_ ), .Y(\dpath/sub/_045_ ) );
sky130_fd_sc_hs__a211oi_1 \dpath/sub/_189_ ( .A1(\dpath/sub/_040_ ), .A2(\dpath/sub/_039_ ), .B1(\dpath/sub/_044_ ), .C1(\dpath/sub/_045_ ), .Y(\dpath/sub/_046_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_190_ ( .A(\dpath/sub/_003_ ), .B(\dpath/sub/_019_ ), .Y(\dpath/sub/_047_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/sub/_191_ ( .A(\dpath/sub/_047_ ), .Y(\dpath/sub/_048_ ) );
sky130_fd_sc_hs__a21o_1 \dpath/sub/_192_ ( .A1(\dpath/sub/_043_ ), .A2(\dpath/sub/_046_ ), .B1(\dpath/sub/_048_ ), .X(\dpath/sub/_049_ ) );
sky130_fd_sc_hs__nand3_1 \dpath/sub/_193_ ( .A(\dpath/sub/_043_ ), .B(\dpath/sub/_046_ ), .C(\dpath/sub/_048_ ), .Y(\dpath/sub/_050_ ) );
sky130_fd_sc_hs__and2_1 \dpath/sub/_194_ ( .A(\dpath/sub/_049_ ), .B(\dpath/sub/_050_ ), .X(\dpath/sub/_108_ ) );
sky130_fd_sc_hs__xor2_1 \dpath/sub/_195_ ( .A(\dpath/sub/_004_ ), .B(\dpath/sub/_020_ ), .X(\dpath/sub/_051_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_196_ ( .A_N(\dpath/sub/_019_ ), .B(\dpath/sub/_003_ ), .X(\dpath/sub/_052_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/sub/_197_ ( .A(\dpath/sub/_052_ ), .Y(\dpath/sub/_053_ ) );
sky130_fd_sc_hs__nand2_1 \dpath/sub/_198_ ( .A(\dpath/sub/_049_ ), .B(\dpath/sub/_053_ ), .Y(\dpath/sub/_054_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_199_ ( .A(\dpath/sub/_051_ ), .B(\dpath/sub/_054_ ), .Y(\dpath/sub/_109_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/sub/_200_ ( .A(\dpath/sub/_020_ ), .B_N(\dpath/sub/_004_ ), .X(\dpath/sub/_055_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/sub/_201_ ( .A1(\dpath/sub/_053_ ), .A2(\dpath/sub/_051_ ), .B1(\dpath/sub/_055_ ), .Y(\dpath/sub/_056_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_202_ ( .A(\dpath/sub/_005_ ), .B(\dpath/sub/_021_ ), .Y(\dpath/sub/_057_ ) );
sky130_fd_sc_hs__a211oi_2 \dpath/sub/_203_ ( .A1(\dpath/sub/_043_ ), .A2(\dpath/sub/_046_ ), .B1(\dpath/sub/_048_ ), .C1(\dpath/sub/_051_ ), .Y(\dpath/sub/_058_ ) );
sky130_fd_sc_hs__or3_1 \dpath/sub/_204_ ( .A(\dpath/sub/_056_ ), .B(\dpath/sub/_057_ ), .C(\dpath/sub/_058_ ), .X(\dpath/sub/_059_ ) );
sky130_fd_sc_hs__o21ai_2 \dpath/sub/_205_ ( .A1(\dpath/sub/_056_ ), .A2(\dpath/sub/_058_ ), .B1(\dpath/sub/_057_ ), .Y(\dpath/sub/_060_ ) );
sky130_fd_sc_hs__and2_1 \dpath/sub/_206_ ( .A(\dpath/sub/_059_ ), .B(\dpath/sub/_060_ ), .X(\dpath/sub/_110_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/sub/_207_ ( .A(\dpath/sub/_021_ ), .B_N(\dpath/sub/_005_ ), .X(\dpath/sub/_061_ ) );
sky130_fd_sc_hs__nand2_1 \dpath/sub/_208_ ( .A(\dpath/sub/_060_ ), .B(\dpath/sub/_061_ ), .Y(\dpath/sub/_062_ ) );
sky130_fd_sc_hs__xnor3_1 \dpath/sub/_209_ ( .A(\dpath/sub/_006_ ), .B(\dpath/sub/_022_ ), .C(\dpath/sub/_062_ ), .X(\dpath/sub/_111_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_210_ ( .A(\dpath/a_lt_b$in0[0] ), .X(\dpath/sub/_000_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_211_ ( .A(\dpath/a_lt_b$in1[0] ), .X(\dpath/sub/_016_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_212_ ( .A(\dpath/sub/_105_ ), .X(\resp_msg[0] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_213_ ( .A(\dpath/a_lt_b$in0[1] ), .X(\dpath/sub/_007_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_214_ ( .A(\dpath/a_lt_b$in1[1] ), .X(\dpath/sub/_023_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_215_ ( .A(\dpath/sub/_112_ ), .X(\resp_msg[1] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_216_ ( .A(\dpath/a_lt_b$in0[2] ), .X(\dpath/sub/_008_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_217_ ( .A(\dpath/a_lt_b$in1[2] ), .X(\dpath/sub/_024_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_218_ ( .A(\dpath/sub/_113_ ), .X(\resp_msg[2] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_219_ ( .A(\dpath/a_lt_b$in0[3] ), .X(\dpath/sub/_009_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_220_ ( .A(\dpath/a_lt_b$in1[3] ), .X(\dpath/sub/_025_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_221_ ( .A(\dpath/sub/_114_ ), .X(\resp_msg[3] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_222_ ( .A(\dpath/a_lt_b$in0[4] ), .X(\dpath/sub/_010_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_223_ ( .A(\dpath/a_lt_b$in1[4] ), .X(\dpath/sub/_026_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_224_ ( .A(\dpath/sub/_115_ ), .X(\resp_msg[4] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_225_ ( .A(\dpath/a_lt_b$in0[5] ), .X(\dpath/sub/_011_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_226_ ( .A(\dpath/a_lt_b$in1[5] ), .X(\dpath/sub/_027_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_227_ ( .A(\dpath/sub/_116_ ), .X(\resp_msg[5] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_228_ ( .A(\dpath/a_lt_b$in0[6] ), .X(\dpath/sub/_012_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_229_ ( .A(\dpath/a_lt_b$in1[6] ), .X(\dpath/sub/_028_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_230_ ( .A(\dpath/sub/_117_ ), .X(\resp_msg[6] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_231_ ( .A(\dpath/a_lt_b$in0[7] ), .X(\dpath/sub/_013_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_232_ ( .A(\dpath/a_lt_b$in1[7] ), .X(\dpath/sub/_029_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_233_ ( .A(\dpath/sub/_118_ ), .X(\resp_msg[7] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_234_ ( .A(\dpath/a_lt_b$in0[8] ), .X(\dpath/sub/_014_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_235_ ( .A(\dpath/a_lt_b$in1[8] ), .X(\dpath/sub/_030_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_236_ ( .A(\dpath/sub/_119_ ), .X(\resp_msg[8] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_237_ ( .A(\dpath/a_lt_b$in0[9] ), .X(\dpath/sub/_015_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_238_ ( .A(\dpath/a_lt_b$in1[9] ), .X(\dpath/sub/_031_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_239_ ( .A(\dpath/sub/_120_ ), .X(\resp_msg[9] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_240_ ( .A(\dpath/a_lt_b$in0[10] ), .X(\dpath/sub/_001_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_241_ ( .A(\dpath/a_lt_b$in1[10] ), .X(\dpath/sub/_017_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_242_ ( .A(\dpath/sub/_106_ ), .X(\resp_msg[10] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_243_ ( .A(\dpath/a_lt_b$in0[11] ), .X(\dpath/sub/_002_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_244_ ( .A(\dpath/a_lt_b$in1[11] ), .X(\dpath/sub/_018_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_245_ ( .A(\dpath/sub/_107_ ), .X(\resp_msg[11] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_246_ ( .A(\dpath/a_lt_b$in0[12] ), .X(\dpath/sub/_003_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_247_ ( .A(\dpath/a_lt_b$in1[12] ), .X(\dpath/sub/_019_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_248_ ( .A(\dpath/sub/_108_ ), .X(\resp_msg[12] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_249_ ( .A(\dpath/a_lt_b$in0[13] ), .X(\dpath/sub/_004_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_250_ ( .A(\dpath/a_lt_b$in1[13] ), .X(\dpath/sub/_020_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_251_ ( .A(\dpath/sub/_109_ ), .X(\resp_msg[13] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_252_ ( .A(\dpath/a_lt_b$in0[14] ), .X(\dpath/sub/_005_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_253_ ( .A(\dpath/a_lt_b$in1[14] ), .X(\dpath/sub/_021_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_254_ ( .A(\dpath/sub/_110_ ), .X(\resp_msg[14] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_255_ ( .A(\dpath/a_lt_b$in0[15] ), .X(\dpath/sub/_006_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_256_ ( .A(\dpath/a_lt_b$in1[15] ), .X(\dpath/sub/_022_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_257_ ( .A(\dpath/sub/_111_ ), .X(\resp_msg[15] ) );
sky130_fd_sc_hs__tap_1 PHY_0 (  );
sky130_fd_sc_hs__tap_1 PHY_1 (  );
sky130_fd_sc_hs__tap_1 PHY_2 (  );
sky130_fd_sc_hs__tap_1 PHY_3 (  );
sky130_fd_sc_hs__tap_1 PHY_4 (  );
sky130_fd_sc_hs__tap_1 PHY_5 (  );
sky130_fd_sc_hs__tap_1 PHY_6 (  );
sky130_fd_sc_hs__tap_1 PHY_7 (  );
sky130_fd_sc_hs__tap_1 PHY_8 (  );
sky130_fd_sc_hs__tap_1 PHY_9 (  );
sky130_fd_sc_hs__tap_1 PHY_10 (  );
sky130_fd_sc_hs__tap_1 PHY_11 (  );
sky130_fd_sc_hs__tap_1 PHY_12 (  );
sky130_fd_sc_hs__tap_1 PHY_13 (  );
sky130_fd_sc_hs__tap_1 PHY_14 (  );
sky130_fd_sc_hs__tap_1 PHY_15 (  );
sky130_fd_sc_hs__tap_1 PHY_16 (  );
sky130_fd_sc_hs__tap_1 PHY_17 (  );
sky130_fd_sc_hs__tap_1 PHY_18 (  );
sky130_fd_sc_hs__tap_1 PHY_19 (  );
sky130_fd_sc_hs__tap_1 PHY_20 (  );
sky130_fd_sc_hs__tap_1 PHY_21 (  );
sky130_fd_sc_hs__tap_1 PHY_22 (  );
sky130_fd_sc_hs__tap_1 PHY_23 (  );
sky130_fd_sc_hs__tap_1 PHY_24 (  );
sky130_fd_sc_hs__tap_1 PHY_25 (  );
sky130_fd_sc_hs__tap_1 PHY_26 (  );
sky130_fd_sc_hs__tap_1 PHY_27 (  );
sky130_fd_sc_hs__tap_1 PHY_28 (  );
sky130_fd_sc_hs__tap_1 PHY_29 (  );
sky130_fd_sc_hs__tap_1 PHY_30 (  );
sky130_fd_sc_hs__tap_1 PHY_31 (  );
sky130_fd_sc_hs__tap_1 PHY_32 (  );
sky130_fd_sc_hs__tap_1 PHY_33 (  );
sky130_fd_sc_hs__tap_1 PHY_34 (  );
sky130_fd_sc_hs__tap_1 PHY_35 (  );
sky130_fd_sc_hs__tap_1 PHY_36 (  );
sky130_fd_sc_hs__tap_1 PHY_37 (  );
sky130_fd_sc_hs__tap_1 PHY_38 (  );
sky130_fd_sc_hs__tap_1 PHY_39 (  );
sky130_fd_sc_hs__tap_1 PHY_40 (  );
sky130_fd_sc_hs__tap_1 PHY_41 (  );
sky130_fd_sc_hs__tap_1 PHY_42 (  );
sky130_fd_sc_hs__tap_1 PHY_43 (  );
sky130_fd_sc_hs__tap_1 PHY_44 (  );
sky130_fd_sc_hs__tap_1 PHY_45 (  );
sky130_fd_sc_hs__tap_1 PHY_46 (  );
sky130_fd_sc_hs__tap_1 PHY_47 (  );
sky130_fd_sc_hs__tap_1 PHY_48 (  );
sky130_fd_sc_hs__tap_1 PHY_49 (  );
sky130_fd_sc_hs__tap_1 PHY_50 (  );
sky130_fd_sc_hs__tap_1 PHY_51 (  );
sky130_fd_sc_hs__tap_1 PHY_52 (  );
sky130_fd_sc_hs__tap_1 PHY_53 (  );
sky130_fd_sc_hs__tap_1 PHY_54 (  );
sky130_fd_sc_hs__tap_1 PHY_55 (  );
sky130_fd_sc_hs__tap_1 PHY_56 (  );
sky130_fd_sc_hs__tap_1 PHY_57 (  );
sky130_fd_sc_hs__tap_1 PHY_58 (  );
sky130_fd_sc_hs__tap_1 PHY_59 (  );
sky130_fd_sc_hs__tap_1 PHY_60 (  );
sky130_fd_sc_hs__tap_1 PHY_61 (  );
sky130_fd_sc_hs__tap_1 PHY_62 (  );
sky130_fd_sc_hs__tap_1 PHY_63 (  );
sky130_fd_sc_hs__tap_1 PHY_64 (  );
sky130_fd_sc_hs__tap_1 PHY_65 (  );
sky130_fd_sc_hs__tap_1 PHY_66 (  );
sky130_fd_sc_hs__tap_1 PHY_67 (  );
sky130_fd_sc_hs__tap_1 PHY_68 (  );
sky130_fd_sc_hs__tap_1 PHY_69 (  );
sky130_fd_sc_hs__tap_1 PHY_70 (  );
sky130_fd_sc_hs__tap_1 PHY_71 (  );
sky130_fd_sc_hs__tap_1 PHY_72 (  );
sky130_fd_sc_hs__tap_1 PHY_73 (  );
sky130_fd_sc_hs__tap_1 PHY_74 (  );
sky130_fd_sc_hs__tap_1 PHY_75 (  );
sky130_fd_sc_hs__tap_1 PHY_76 (  );
sky130_fd_sc_hs__tap_1 PHY_77 (  );
sky130_fd_sc_hs__tap_1 PHY_78 (  );
sky130_fd_sc_hs__tap_1 PHY_79 (  );
sky130_fd_sc_hs__tap_1 PHY_80 (  );
sky130_fd_sc_hs__tap_1 PHY_81 (  );
sky130_fd_sc_hs__tap_1 PHY_82 (  );
sky130_fd_sc_hs__tap_1 PHY_83 (  );
sky130_fd_sc_hs__tap_1 PHY_84 (  );
sky130_fd_sc_hs__tap_1 PHY_85 (  );
sky130_fd_sc_hs__tap_1 PHY_86 (  );
sky130_fd_sc_hs__tap_1 PHY_87 (  );
sky130_fd_sc_hs__tap_1 PHY_88 (  );
sky130_fd_sc_hs__tap_1 PHY_89 (  );
sky130_fd_sc_hs__tap_1 PHY_90 (  );
sky130_fd_sc_hs__tap_1 PHY_91 (  );
sky130_fd_sc_hs__tap_1 PHY_92 (  );
sky130_fd_sc_hs__tap_1 PHY_93 (  );
sky130_fd_sc_hs__tap_1 PHY_94 (  );
sky130_fd_sc_hs__tap_1 PHY_95 (  );
sky130_fd_sc_hs__tap_1 PHY_96 (  );
sky130_fd_sc_hs__tap_1 PHY_97 (  );
sky130_fd_sc_hs__tap_1 PHY_98 (  );
sky130_fd_sc_hs__tap_1 PHY_99 (  );
sky130_fd_sc_hs__tap_1 PHY_100 (  );
sky130_fd_sc_hs__tap_1 PHY_101 (  );
sky130_fd_sc_hs__tap_1 PHY_102 (  );
sky130_fd_sc_hs__tap_1 PHY_103 (  );
sky130_fd_sc_hs__tap_1 PHY_104 (  );
sky130_fd_sc_hs__tap_1 PHY_105 (  );
sky130_fd_sc_hs__tap_1 PHY_106 (  );
sky130_fd_sc_hs__tap_1 PHY_107 (  );
sky130_fd_sc_hs__tap_1 PHY_108 (  );
sky130_fd_sc_hs__tap_1 PHY_109 (  );
sky130_fd_sc_hs__tap_1 PHY_110 (  );
sky130_fd_sc_hs__tap_1 PHY_111 (  );
sky130_fd_sc_hs__tap_1 PHY_112 (  );
sky130_fd_sc_hs__tap_1 PHY_113 (  );
sky130_fd_sc_hs__tap_1 PHY_114 (  );
sky130_fd_sc_hs__tap_1 PHY_115 (  );
sky130_fd_sc_hs__tap_1 PHY_116 (  );
sky130_fd_sc_hs__tap_1 PHY_117 (  );
sky130_fd_sc_hs__tap_1 PHY_118 (  );
sky130_fd_sc_hs__tap_1 PHY_119 (  );
sky130_fd_sc_hs__tap_1 PHY_120 (  );
sky130_fd_sc_hs__tap_1 PHY_121 (  );
sky130_fd_sc_hs__tap_1 PHY_122 (  );
sky130_fd_sc_hs__tap_1 PHY_123 (  );
sky130_fd_sc_hs__tap_1 PHY_124 (  );
sky130_fd_sc_hs__tap_1 PHY_125 (  );
sky130_fd_sc_hs__tap_1 PHY_126 (  );
sky130_fd_sc_hs__tap_1 PHY_127 (  );
sky130_fd_sc_hs__tap_1 PHY_128 (  );
sky130_fd_sc_hs__tap_1 PHY_129 (  );
sky130_fd_sc_hs__tap_1 PHY_130 (  );
sky130_fd_sc_hs__tap_1 PHY_131 (  );
sky130_fd_sc_hs__tap_1 PHY_132 (  );
sky130_fd_sc_hs__tap_1 PHY_133 (  );
sky130_fd_sc_hs__tap_1 PHY_134 (  );
sky130_fd_sc_hs__tap_1 PHY_135 (  );
sky130_fd_sc_hs__tap_1 PHY_136 (  );
sky130_fd_sc_hs__tap_1 PHY_137 (  );
sky130_fd_sc_hs__tap_1 PHY_138 (  );
sky130_fd_sc_hs__tap_1 PHY_139 (  );
sky130_fd_sc_hs__tap_1 PHY_140 (  );
sky130_fd_sc_hs__tap_1 PHY_141 (  );
sky130_fd_sc_hs__tap_1 PHY_142 (  );
sky130_fd_sc_hs__tap_1 PHY_143 (  );
sky130_fd_sc_hs__tap_1 PHY_144 (  );
sky130_fd_sc_hs__tap_1 PHY_145 (  );
sky130_fd_sc_hs__tap_1 PHY_146 (  );
sky130_fd_sc_hs__tap_1 PHY_147 (  );
sky130_fd_sc_hs__tap_1 PHY_148 (  );
sky130_fd_sc_hs__tap_1 PHY_149 (  );
sky130_fd_sc_hs__tap_1 PHY_150 (  );
sky130_fd_sc_hs__tap_1 PHY_151 (  );
sky130_fd_sc_hs__tap_1 PHY_152 (  );
sky130_fd_sc_hs__tap_1 PHY_153 (  );
sky130_fd_sc_hs__tap_1 PHY_154 (  );
sky130_fd_sc_hs__tap_1 PHY_155 (  );
sky130_fd_sc_hs__tap_1 PHY_156 (  );
sky130_fd_sc_hs__tap_1 PHY_157 (  );
sky130_fd_sc_hs__tap_1 PHY_158 (  );
sky130_fd_sc_hs__tap_1 PHY_159 (  );
sky130_fd_sc_hs__tap_1 PHY_160 (  );
sky130_fd_sc_hs__tap_1 PHY_161 (  );
sky130_fd_sc_hs__tap_1 PHY_162 (  );
sky130_fd_sc_hs__tap_1 PHY_163 (  );
sky130_fd_sc_hs__tap_1 PHY_164 (  );
sky130_fd_sc_hs__tap_1 PHY_165 (  );
sky130_fd_sc_hs__tap_1 PHY_166 (  );
sky130_fd_sc_hs__tap_1 PHY_167 (  );
sky130_fd_sc_hs__tap_1 PHY_168 (  );
sky130_fd_sc_hs__tap_1 PHY_169 (  );
sky130_fd_sc_hs__tap_1 PHY_170 (  );
sky130_fd_sc_hs__tap_1 PHY_171 (  );
sky130_fd_sc_hs__tap_1 PHY_172 (  );
sky130_fd_sc_hs__tap_1 PHY_173 (  );
sky130_fd_sc_hs__tap_1 PHY_174 (  );
sky130_fd_sc_hs__tap_1 PHY_175 (  );
sky130_fd_sc_hs__tap_1 PHY_176 (  );
sky130_fd_sc_hs__tap_1 PHY_177 (  );
sky130_fd_sc_hs__tap_1 PHY_178 (  );
sky130_fd_sc_hs__tap_1 PHY_179 (  );
sky130_fd_sc_hs__tap_1 PHY_180 (  );
sky130_fd_sc_hs__tap_1 PHY_181 (  );
sky130_fd_sc_hs__tap_1 PHY_182 (  );
sky130_fd_sc_hs__tap_1 PHY_183 (  );
sky130_fd_sc_hs__tap_1 PHY_184 (  );
sky130_fd_sc_hs__tap_1 PHY_185 (  );
sky130_fd_sc_hs__tap_1 PHY_186 (  );
sky130_fd_sc_hs__tap_1 PHY_187 (  );
sky130_fd_sc_hs__tap_1 PHY_188 (  );
sky130_fd_sc_hs__tap_1 PHY_189 (  );
sky130_fd_sc_hs__tap_1 PHY_190 (  );
sky130_fd_sc_hs__tap_1 PHY_191 (  );
sky130_fd_sc_hs__tap_1 PHY_192 (  );
sky130_fd_sc_hs__tap_1 PHY_193 (  );
sky130_fd_sc_hs__tap_1 PHY_194 (  );
sky130_fd_sc_hs__tap_1 PHY_195 (  );
sky130_fd_sc_hs__tap_1 PHY_196 (  );
sky130_fd_sc_hs__tap_1 PHY_197 (  );
sky130_fd_sc_hs__tap_1 PHY_198 (  );
sky130_fd_sc_hs__tap_1 PHY_199 (  );
sky130_fd_sc_hs__tap_1 PHY_200 (  );
sky130_fd_sc_hs__tap_1 PHY_201 (  );
sky130_fd_sc_hs__tap_1 PHY_202 (  );
sky130_fd_sc_hs__tap_1 PHY_203 (  );
sky130_fd_sc_hs__tap_1 PHY_204 (  );
sky130_fd_sc_hs__tap_1 PHY_205 (  );
sky130_fd_sc_hs__tap_1 PHY_206 (  );
sky130_fd_sc_hs__tap_1 PHY_207 (  );
sky130_fd_sc_hs__tap_1 PHY_208 (  );
sky130_fd_sc_hs__tap_1 PHY_209 (  );
sky130_fd_sc_hs__tap_1 PHY_210 (  );
sky130_fd_sc_hs__tap_1 PHY_211 (  );
sky130_fd_sc_hs__tap_1 PHY_212 (  );
sky130_fd_sc_hs__tap_1 PHY_213 (  );
sky130_fd_sc_hs__tap_1 PHY_214 (  );
sky130_fd_sc_hs__tap_1 PHY_215 (  );
sky130_fd_sc_hs__tap_1 PHY_216 (  );
sky130_fd_sc_hs__tap_1 PHY_217 (  );
sky130_fd_sc_hs__tap_1 PHY_218 (  );
sky130_fd_sc_hs__tap_1 PHY_219 (  );
sky130_fd_sc_hs__tap_1 PHY_220 (  );
sky130_fd_sc_hs__tap_1 PHY_221 (  );
sky130_fd_sc_hs__tap_1 PHY_222 (  );
sky130_fd_sc_hs__tap_1 PHY_223 (  );
sky130_fd_sc_hs__tap_1 PHY_224 (  );
sky130_fd_sc_hs__tap_1 PHY_225 (  );
sky130_fd_sc_hs__tap_1 PHY_226 (  );
sky130_fd_sc_hs__tap_1 PHY_227 (  );
sky130_fd_sc_hs__tap_1 PHY_228 (  );
sky130_fd_sc_hs__tap_1 PHY_229 (  );
sky130_fd_sc_hs__tap_1 PHY_230 (  );
sky130_fd_sc_hs__tap_1 PHY_231 (  );
sky130_fd_sc_hs__tap_1 PHY_232 (  );
sky130_fd_sc_hs__tap_1 PHY_233 (  );
sky130_fd_sc_hs__tap_1 PHY_234 (  );
sky130_fd_sc_hs__tap_1 PHY_235 (  );
sky130_fd_sc_hs__tap_1 PHY_236 (  );
sky130_fd_sc_hs__tap_1 PHY_237 (  );
sky130_fd_sc_hs__tap_1 PHY_238 (  );
sky130_fd_sc_hs__tap_1 PHY_239 (  );
sky130_fd_sc_hs__tap_1 PHY_240 (  );
sky130_fd_sc_hs__tap_1 PHY_241 (  );
sky130_fd_sc_hs__tap_1 PHY_242 (  );
sky130_fd_sc_hs__tap_1 PHY_243 (  );
sky130_fd_sc_hs__tap_1 PHY_244 (  );
sky130_fd_sc_hs__tap_1 PHY_245 (  );
sky130_fd_sc_hs__tap_1 PHY_246 (  );
sky130_fd_sc_hs__tap_1 PHY_247 (  );
sky130_fd_sc_hs__tap_1 PHY_248 (  );
sky130_fd_sc_hs__tap_1 PHY_249 (  );
sky130_fd_sc_hs__tap_1 PHY_250 (  );
sky130_fd_sc_hs__tap_1 PHY_251 (  );
sky130_fd_sc_hs__tap_1 PHY_252 (  );
sky130_fd_sc_hs__tap_1 PHY_253 (  );
sky130_fd_sc_hs__tap_1 PHY_254 (  );
sky130_fd_sc_hs__tap_1 PHY_255 (  );
sky130_fd_sc_hs__tap_1 PHY_256 (  );
sky130_fd_sc_hs__tap_1 PHY_257 (  );
sky130_fd_sc_hs__tap_1 PHY_258 (  );
sky130_fd_sc_hs__tap_1 PHY_259 (  );
sky130_fd_sc_hs__tap_1 PHY_260 (  );
sky130_fd_sc_hs__tap_1 PHY_261 (  );
sky130_fd_sc_hs__tap_1 PHY_262 (  );
sky130_fd_sc_hs__tap_1 PHY_263 (  );
sky130_fd_sc_hs__tap_1 PHY_264 (  );
sky130_fd_sc_hs__tap_1 PHY_265 (  );
sky130_fd_sc_hs__tap_1 PHY_266 (  );
sky130_fd_sc_hs__tap_1 PHY_267 (  );
sky130_fd_sc_hs__tap_1 PHY_268 (  );
sky130_fd_sc_hs__tap_1 PHY_269 (  );
sky130_fd_sc_hs__tap_1 PHY_270 (  );
sky130_fd_sc_hs__tap_1 PHY_271 (  );
sky130_fd_sc_hs__tap_1 PHY_272 (  );
sky130_fd_sc_hs__tap_1 PHY_273 (  );
sky130_fd_sc_hs__tap_1 PHY_274 (  );
sky130_fd_sc_hs__tap_1 PHY_275 (  );
sky130_fd_sc_hs__tap_1 PHY_276 (  );
sky130_fd_sc_hs__tap_1 PHY_277 (  );
sky130_fd_sc_hs__tap_1 PHY_278 (  );
sky130_fd_sc_hs__tap_1 PHY_279 (  );
sky130_fd_sc_hs__tap_1 PHY_280 (  );
sky130_fd_sc_hs__tap_1 PHY_281 (  );
sky130_fd_sc_hs__tap_1 PHY_282 (  );
sky130_fd_sc_hs__tap_1 PHY_283 (  );
sky130_fd_sc_hs__tap_1 PHY_284 (  );
sky130_fd_sc_hs__tap_1 PHY_285 (  );
sky130_fd_sc_hs__tap_1 PHY_286 (  );
sky130_fd_sc_hs__tap_1 PHY_287 (  );
sky130_fd_sc_hs__tap_1 PHY_288 (  );
sky130_fd_sc_hs__tap_1 PHY_289 (  );
sky130_fd_sc_hs__tap_1 PHY_290 (  );
sky130_fd_sc_hs__tap_1 PHY_291 (  );
sky130_fd_sc_hs__tap_1 PHY_292 (  );
sky130_fd_sc_hs__tap_1 PHY_293 (  );
sky130_fd_sc_hs__tap_1 PHY_294 (  );
sky130_fd_sc_hs__tap_1 PHY_295 (  );
sky130_fd_sc_hs__tap_1 PHY_296 (  );
sky130_fd_sc_hs__tap_1 PHY_297 (  );
sky130_fd_sc_hs__tap_1 PHY_298 (  );
sky130_fd_sc_hs__tap_1 PHY_299 (  );
sky130_fd_sc_hs__tap_1 PHY_300 (  );
sky130_fd_sc_hs__tap_1 PHY_301 (  );
sky130_fd_sc_hs__tap_1 PHY_302 (  );
sky130_fd_sc_hs__tap_1 PHY_303 (  );
sky130_fd_sc_hs__tap_1 PHY_304 (  );
sky130_fd_sc_hs__tap_1 PHY_305 (  );
sky130_fd_sc_hs__tap_1 PHY_306 (  );
sky130_fd_sc_hs__tap_1 PHY_307 (  );
sky130_fd_sc_hs__tap_1 PHY_308 (  );
sky130_fd_sc_hs__tap_1 PHY_309 (  );
sky130_fd_sc_hs__tap_1 PHY_310 (  );
sky130_fd_sc_hs__tap_1 PHY_311 (  );
sky130_fd_sc_hs__tap_1 PHY_312 (  );
sky130_fd_sc_hs__tap_1 PHY_313 (  );
sky130_fd_sc_hs__tap_1 PHY_314 (  );
sky130_fd_sc_hs__tap_1 PHY_315 (  );
sky130_fd_sc_hs__tap_1 PHY_316 (  );
sky130_fd_sc_hs__tap_1 PHY_317 (  );
sky130_fd_sc_hs__tap_1 PHY_318 (  );
sky130_fd_sc_hs__tap_1 PHY_319 (  );
sky130_fd_sc_hs__tap_1 PHY_320 (  );
sky130_fd_sc_hs__tap_1 PHY_321 (  );
sky130_fd_sc_hs__tap_1 PHY_322 (  );
sky130_fd_sc_hs__tap_1 PHY_323 (  );
sky130_fd_sc_hs__tap_1 PHY_324 (  );
sky130_fd_sc_hs__tap_1 PHY_325 (  );
sky130_fd_sc_hs__tap_1 PHY_326 (  );
sky130_fd_sc_hs__tap_1 PHY_327 (  );
sky130_fd_sc_hs__tap_1 PHY_328 (  );
sky130_fd_sc_hs__tap_1 PHY_329 (  );
sky130_fd_sc_hs__tap_1 PHY_330 (  );
sky130_fd_sc_hs__tap_1 PHY_331 (  );
sky130_fd_sc_hs__tap_1 PHY_332 (  );
sky130_fd_sc_hs__tap_1 PHY_333 (  );
sky130_fd_sc_hs__tap_1 PHY_334 (  );
sky130_fd_sc_hs__tap_1 PHY_335 (  );
sky130_fd_sc_hs__tap_1 PHY_336 (  );
sky130_fd_sc_hs__tap_1 PHY_337 (  );
sky130_fd_sc_hs__tap_1 PHY_338 (  );
sky130_fd_sc_hs__tap_1 PHY_339 (  );
sky130_fd_sc_hs__tap_1 PHY_340 (  );
sky130_fd_sc_hs__tap_1 PHY_341 (  );
sky130_fd_sc_hs__tap_1 PHY_342 (  );
sky130_fd_sc_hs__tap_1 PHY_343 (  );
sky130_fd_sc_hs__tap_1 PHY_344 (  );
sky130_fd_sc_hs__tap_1 PHY_345 (  );
sky130_fd_sc_hs__tap_1 PHY_346 (  );
sky130_fd_sc_hs__tap_1 PHY_347 (  );
sky130_fd_sc_hs__tap_1 PHY_348 (  );
sky130_fd_sc_hs__tap_1 PHY_349 (  );
sky130_fd_sc_hs__tap_1 PHY_350 (  );
sky130_fd_sc_hs__tap_1 PHY_351 (  );
sky130_fd_sc_hs__tap_1 PHY_352 (  );
sky130_fd_sc_hs__tap_1 PHY_353 (  );
sky130_fd_sc_hs__tap_1 PHY_354 (  );
sky130_fd_sc_hs__tap_1 PHY_355 (  );
sky130_fd_sc_hs__tap_1 PHY_356 (  );
sky130_fd_sc_hs__tap_1 PHY_357 (  );
sky130_fd_sc_hs__tap_1 PHY_358 (  );
sky130_fd_sc_hs__tap_1 PHY_359 (  );
sky130_fd_sc_hs__tap_1 PHY_360 (  );
sky130_fd_sc_hs__tap_1 PHY_361 (  );
sky130_fd_sc_hs__tap_1 PHY_362 (  );
sky130_fd_sc_hs__tap_1 PHY_363 (  );
sky130_fd_sc_hs__tap_1 PHY_364 (  );
sky130_fd_sc_hs__tap_1 PHY_365 (  );
sky130_fd_sc_hs__tap_1 PHY_366 (  );
sky130_fd_sc_hs__tap_1 PHY_367 (  );
sky130_fd_sc_hs__tap_1 PHY_368 (  );
sky130_fd_sc_hs__tap_1 PHY_369 (  );
sky130_fd_sc_hs__tap_1 PHY_370 (  );
sky130_fd_sc_hs__tap_1 PHY_371 (  );
sky130_fd_sc_hs__tap_1 PHY_372 (  );
sky130_fd_sc_hs__tap_1 PHY_373 (  );
sky130_fd_sc_hs__tap_1 PHY_374 (  );
sky130_fd_sc_hs__tap_1 PHY_375 (  );
sky130_fd_sc_hs__tap_1 PHY_376 (  );
sky130_fd_sc_hs__tap_1 PHY_377 (  );
sky130_fd_sc_hs__tap_1 PHY_378 (  );
sky130_fd_sc_hs__tap_1 PHY_379 (  );
sky130_fd_sc_hs__tap_1 PHY_380 (  );
sky130_fd_sc_hs__tap_1 PHY_381 (  );
sky130_fd_sc_hs__tap_1 PHY_382 (  );
sky130_fd_sc_hs__tap_1 PHY_383 (  );
sky130_fd_sc_hs__tap_1 PHY_384 (  );
sky130_fd_sc_hs__tap_1 PHY_385 (  );
sky130_fd_sc_hs__tap_1 PHY_386 (  );
sky130_fd_sc_hs__tap_1 PHY_387 (  );
sky130_fd_sc_hs__tap_1 PHY_388 (  );
sky130_fd_sc_hs__tap_1 PHY_389 (  );
sky130_fd_sc_hs__tap_1 PHY_390 (  );
sky130_fd_sc_hs__tap_1 PHY_391 (  );
sky130_fd_sc_hs__tap_1 PHY_392 (  );
sky130_fd_sc_hs__tap_1 PHY_393 (  );
sky130_fd_sc_hs__tap_1 PHY_394 (  );
sky130_fd_sc_hs__tap_1 PHY_395 (  );
sky130_fd_sc_hs__tap_1 PHY_396 (  );
sky130_fd_sc_hs__tap_1 PHY_397 (  );
sky130_fd_sc_hs__tap_1 PHY_398 (  );
sky130_fd_sc_hs__tap_1 PHY_399 (  );
sky130_fd_sc_hs__tap_1 PHY_400 (  );
sky130_fd_sc_hs__tap_1 PHY_401 (  );
sky130_fd_sc_hs__tap_1 PHY_402 (  );
sky130_fd_sc_hs__tap_1 PHY_403 (  );
sky130_fd_sc_hs__tap_1 PHY_404 (  );
sky130_fd_sc_hs__tap_1 PHY_405 (  );
sky130_fd_sc_hs__tap_1 PHY_406 (  );
sky130_fd_sc_hs__tap_1 PHY_407 (  );
sky130_fd_sc_hs__tap_1 PHY_408 (  );
sky130_fd_sc_hs__tap_1 PHY_409 (  );
sky130_fd_sc_hs__tap_1 PHY_410 (  );
sky130_fd_sc_hs__tap_1 PHY_411 (  );
sky130_fd_sc_hs__tap_1 PHY_412 (  );
sky130_fd_sc_hs__tap_1 PHY_413 (  );
sky130_fd_sc_hs__tap_1 PHY_414 (  );
sky130_fd_sc_hs__tap_1 PHY_415 (  );
sky130_fd_sc_hs__tap_1 PHY_416 (  );
sky130_fd_sc_hs__tap_1 PHY_417 (  );
sky130_fd_sc_hs__tap_1 PHY_418 (  );
sky130_fd_sc_hs__tap_1 PHY_419 (  );
sky130_fd_sc_hs__tap_1 PHY_420 (  );
sky130_fd_sc_hs__tap_1 PHY_421 (  );
sky130_fd_sc_hs__tap_1 PHY_422 (  );
sky130_fd_sc_hs__tap_1 PHY_423 (  );
sky130_fd_sc_hs__tap_1 PHY_424 (  );
sky130_fd_sc_hs__tap_1 PHY_425 (  );
sky130_fd_sc_hs__tap_1 PHY_426 (  );
sky130_fd_sc_hs__tap_1 PHY_427 (  );
sky130_fd_sc_hs__tap_1 PHY_428 (  );
sky130_fd_sc_hs__tap_1 PHY_429 (  );
sky130_fd_sc_hs__tap_1 PHY_430 (  );
sky130_fd_sc_hs__tap_1 PHY_431 (  );
sky130_fd_sc_hs__tap_1 PHY_432 (  );
sky130_fd_sc_hs__tap_1 PHY_433 (  );
sky130_fd_sc_hs__tap_1 PHY_434 (  );
sky130_fd_sc_hs__tap_1 PHY_435 (  );
sky130_fd_sc_hs__tap_1 PHY_436 (  );
sky130_fd_sc_hs__tap_1 PHY_437 (  );
sky130_fd_sc_hs__tap_1 PHY_438 (  );
sky130_fd_sc_hs__tap_1 PHY_439 (  );
sky130_fd_sc_hs__tap_1 PHY_440 (  );
sky130_fd_sc_hs__tap_1 PHY_441 (  );
sky130_fd_sc_hs__tap_1 PHY_442 (  );
sky130_fd_sc_hs__tap_1 PHY_443 (  );
sky130_fd_sc_hs__tap_1 PHY_444 (  );
sky130_fd_sc_hs__tap_1 PHY_445 (  );
sky130_fd_sc_hs__tap_1 PHY_446 (  );
sky130_fd_sc_hs__tap_1 PHY_447 (  );
sky130_fd_sc_hs__tap_1 PHY_448 (  );
sky130_fd_sc_hs__tap_1 PHY_449 (  );
sky130_fd_sc_hs__tap_1 PHY_450 (  );
sky130_fd_sc_hs__tap_1 PHY_451 (  );
sky130_fd_sc_hs__tap_1 PHY_452 (  );
sky130_fd_sc_hs__tap_1 PHY_453 (  );
sky130_fd_sc_hs__tap_1 PHY_454 (  );
sky130_fd_sc_hs__tap_1 PHY_455 (  );
sky130_fd_sc_hs__tap_1 PHY_456 (  );
sky130_fd_sc_hs__tap_1 PHY_457 (  );
sky130_fd_sc_hs__tap_1 PHY_458 (  );
sky130_fd_sc_hs__tap_1 PHY_459 (  );
sky130_fd_sc_hs__tap_1 PHY_460 (  );
sky130_fd_sc_hs__tap_1 PHY_461 (  );
sky130_fd_sc_hs__tap_1 PHY_462 (  );
sky130_fd_sc_hs__tap_1 PHY_463 (  );
sky130_fd_sc_hs__tap_1 PHY_464 (  );
sky130_fd_sc_hs__tap_1 PHY_465 (  );
sky130_fd_sc_hs__tap_1 PHY_466 (  );
sky130_fd_sc_hs__tap_1 PHY_467 (  );
sky130_fd_sc_hs__tap_1 PHY_468 (  );
sky130_fd_sc_hs__tap_1 PHY_469 (  );
sky130_fd_sc_hs__tap_1 PHY_470 (  );
sky130_fd_sc_hs__tap_1 PHY_471 (  );
sky130_fd_sc_hs__tap_1 PHY_472 (  );
sky130_fd_sc_hs__tap_1 PHY_473 (  );
sky130_fd_sc_hs__tap_1 PHY_474 (  );
sky130_fd_sc_hs__tap_1 PHY_475 (  );
sky130_fd_sc_hs__tap_1 PHY_476 (  );
sky130_fd_sc_hs__tap_1 PHY_477 (  );
sky130_fd_sc_hs__tap_1 PHY_478 (  );
sky130_fd_sc_hs__tap_1 PHY_479 (  );
sky130_fd_sc_hs__tap_1 PHY_480 (  );
sky130_fd_sc_hs__tap_1 PHY_481 (  );
sky130_fd_sc_hs__tap_1 PHY_482 (  );
sky130_fd_sc_hs__tap_1 PHY_483 (  );
sky130_fd_sc_hs__tap_1 PHY_484 (  );
sky130_fd_sc_hs__tap_1 PHY_485 (  );
sky130_fd_sc_hs__tap_1 PHY_486 (  );
sky130_fd_sc_hs__tap_1 PHY_487 (  );
sky130_fd_sc_hs__tap_1 PHY_488 (  );
sky130_fd_sc_hs__tap_1 PHY_489 (  );
sky130_fd_sc_hs__tap_1 PHY_490 (  );
sky130_fd_sc_hs__tap_1 PHY_491 (  );
sky130_fd_sc_hs__tap_1 PHY_492 (  );
sky130_fd_sc_hs__tap_1 PHY_493 (  );
sky130_fd_sc_hs__tap_1 PHY_494 (  );
sky130_fd_sc_hs__tap_1 PHY_495 (  );
sky130_fd_sc_hs__tap_1 PHY_496 (  );
sky130_fd_sc_hs__tap_1 PHY_497 (  );
sky130_fd_sc_hs__tap_1 PHY_498 (  );
sky130_fd_sc_hs__tap_1 PHY_499 (  );
sky130_fd_sc_hs__tap_1 PHY_500 (  );
sky130_fd_sc_hs__tap_1 PHY_501 (  );
sky130_fd_sc_hs__tap_1 PHY_502 (  );
sky130_fd_sc_hs__tap_1 PHY_503 (  );
sky130_fd_sc_hs__tap_1 PHY_504 (  );
sky130_fd_sc_hs__tap_1 PHY_505 (  );
sky130_fd_sc_hs__tap_1 PHY_506 (  );
sky130_fd_sc_hs__tap_1 PHY_507 (  );
sky130_fd_sc_hs__tap_1 PHY_508 (  );
sky130_fd_sc_hs__tap_1 PHY_509 (  );
sky130_fd_sc_hs__tap_1 PHY_510 (  );
sky130_fd_sc_hs__tap_1 PHY_511 (  );
sky130_fd_sc_hs__tap_1 PHY_512 (  );
sky130_fd_sc_hs__tap_1 PHY_513 (  );
sky130_fd_sc_hs__tap_1 PHY_514 (  );
sky130_fd_sc_hs__tap_1 PHY_515 (  );
sky130_fd_sc_hs__tap_1 PHY_516 (  );
sky130_fd_sc_hs__tap_1 PHY_517 (  );
sky130_fd_sc_hs__tap_1 PHY_518 (  );
sky130_fd_sc_hs__tap_1 PHY_519 (  );
sky130_fd_sc_hs__tap_1 PHY_520 (  );
sky130_fd_sc_hs__tap_1 PHY_521 (  );
sky130_fd_sc_hs__tap_1 PHY_522 (  );
sky130_fd_sc_hs__tap_1 PHY_523 (  );
sky130_fd_sc_hs__tap_1 PHY_524 (  );
sky130_fd_sc_hs__tap_1 PHY_525 (  );
sky130_fd_sc_hs__tap_1 PHY_526 (  );
sky130_fd_sc_hs__tap_1 PHY_527 (  );
sky130_fd_sc_hs__tap_1 PHY_528 (  );
sky130_fd_sc_hs__tap_1 PHY_529 (  );
sky130_fd_sc_hs__tap_1 PHY_530 (  );
sky130_fd_sc_hs__tap_1 PHY_531 (  );
sky130_fd_sc_hs__tap_1 PHY_532 (  );
sky130_fd_sc_hs__tap_1 PHY_533 (  );
sky130_fd_sc_hs__tap_1 PHY_534 (  );
sky130_fd_sc_hs__tap_1 PHY_535 (  );
sky130_fd_sc_hs__tap_1 PHY_536 (  );
sky130_fd_sc_hs__tap_1 PHY_537 (  );
sky130_fd_sc_hs__tap_1 PHY_538 (  );
sky130_fd_sc_hs__tap_1 PHY_539 (  );
sky130_fd_sc_hs__tap_1 PHY_540 (  );
sky130_fd_sc_hs__tap_1 PHY_541 (  );
sky130_fd_sc_hs__tap_1 PHY_542 (  );
sky130_fd_sc_hs__tap_1 PHY_543 (  );
sky130_fd_sc_hs__tap_1 PHY_544 (  );
sky130_fd_sc_hs__tap_1 PHY_545 (  );
sky130_fd_sc_hs__tap_1 PHY_546 (  );
sky130_fd_sc_hs__tap_1 PHY_547 (  );
sky130_fd_sc_hs__tap_1 PHY_548 (  );
sky130_fd_sc_hs__tap_1 PHY_549 (  );
sky130_fd_sc_hs__tap_1 PHY_550 (  );
sky130_fd_sc_hs__tap_1 PHY_551 (  );
sky130_fd_sc_hs__tap_1 PHY_552 (  );
sky130_fd_sc_hs__tap_1 PHY_553 (  );
sky130_fd_sc_hs__tap_1 PHY_554 (  );
sky130_fd_sc_hs__tap_1 PHY_555 (  );
sky130_fd_sc_hs__tap_1 PHY_556 (  );
sky130_fd_sc_hs__tap_1 PHY_557 (  );
sky130_fd_sc_hs__tap_1 PHY_558 (  );
sky130_fd_sc_hs__tap_1 PHY_559 (  );
sky130_fd_sc_hs__tap_1 PHY_560 (  );
sky130_fd_sc_hs__tap_1 PHY_561 (  );
sky130_fd_sc_hs__tap_1 PHY_562 (  );
sky130_fd_sc_hs__tap_1 PHY_563 (  );
sky130_fd_sc_hs__tap_1 PHY_564 (  );
sky130_fd_sc_hs__tap_1 PHY_565 (  );
sky130_fd_sc_hs__tap_1 PHY_566 (  );
sky130_fd_sc_hs__tap_1 PHY_567 (  );
sky130_fd_sc_hs__tap_1 PHY_568 (  );
sky130_fd_sc_hs__tap_1 PHY_569 (  );
sky130_fd_sc_hs__tap_1 PHY_570 (  );
sky130_fd_sc_hs__tap_1 PHY_571 (  );
sky130_fd_sc_hs__tap_1 PHY_572 (  );
sky130_fd_sc_hs__tap_1 PHY_573 (  );
sky130_fd_sc_hs__tap_1 PHY_574 (  );
sky130_fd_sc_hs__tap_1 PHY_575 (  );
sky130_fd_sc_hs__tap_1 PHY_576 (  );
sky130_fd_sc_hs__tap_1 PHY_577 (  );
sky130_fd_sc_hs__tap_1 PHY_578 (  );
sky130_fd_sc_hs__tap_1 PHY_579 (  );
sky130_fd_sc_hs__tap_1 PHY_580 (  );
sky130_fd_sc_hs__tap_1 PHY_581 (  );
sky130_fd_sc_hs__tap_1 PHY_582 (  );
sky130_fd_sc_hs__tap_1 PHY_583 (  );
sky130_fd_sc_hs__tap_1 PHY_584 (  );
sky130_fd_sc_hs__tap_1 PHY_585 (  );
sky130_fd_sc_hs__tap_1 PHY_586 (  );
sky130_fd_sc_hs__tap_1 PHY_587 (  );
sky130_fd_sc_hs__tap_1 PHY_588 (  );
sky130_fd_sc_hs__tap_1 PHY_589 (  );
sky130_fd_sc_hs__tap_1 PHY_590 (  );
sky130_fd_sc_hs__tap_1 PHY_591 (  );
sky130_fd_sc_hs__tap_1 PHY_592 (  );
sky130_fd_sc_hs__tap_1 PHY_593 (  );
sky130_fd_sc_hs__tap_1 PHY_594 (  );
sky130_fd_sc_hs__tap_1 PHY_595 (  );
sky130_fd_sc_hs__tap_1 PHY_596 (  );
sky130_fd_sc_hs__tap_1 PHY_597 (  );
sky130_fd_sc_hs__tap_1 PHY_598 (  );
sky130_fd_sc_hs__tap_1 PHY_599 (  );
sky130_fd_sc_hs__tap_1 PHY_600 (  );
sky130_fd_sc_hs__tap_1 PHY_601 (  );
sky130_fd_sc_hs__tap_1 PHY_602 (  );
sky130_fd_sc_hs__tap_1 PHY_603 (  );
sky130_fd_sc_hs__tap_1 PHY_604 (  );
sky130_fd_sc_hs__tap_1 PHY_605 (  );
sky130_fd_sc_hs__tap_1 PHY_606 (  );
sky130_fd_sc_hs__tap_1 PHY_607 (  );
sky130_fd_sc_hs__tap_1 PHY_608 (  );
sky130_fd_sc_hs__tap_1 PHY_609 (  );
sky130_fd_sc_hs__tap_1 PHY_610 (  );
sky130_fd_sc_hs__tap_1 PHY_611 (  );
sky130_fd_sc_hs__tap_1 PHY_612 (  );
sky130_fd_sc_hs__tap_1 PHY_613 (  );
sky130_fd_sc_hs__tap_1 PHY_614 (  );
sky130_fd_sc_hs__tap_1 PHY_615 (  );
sky130_fd_sc_hs__tap_1 PHY_616 (  );
sky130_fd_sc_hs__tap_1 PHY_617 (  );
sky130_fd_sc_hs__tap_1 PHY_618 (  );
sky130_fd_sc_hs__tap_1 PHY_619 (  );
sky130_fd_sc_hs__tap_1 PHY_620 (  );
sky130_fd_sc_hs__tap_1 PHY_621 (  );
sky130_fd_sc_hs__tap_1 PHY_622 (  );
sky130_fd_sc_hs__tap_1 PHY_623 (  );
sky130_fd_sc_hs__tap_1 PHY_624 (  );
sky130_fd_sc_hs__tap_1 PHY_625 (  );
sky130_fd_sc_hs__tap_1 PHY_626 (  );
sky130_fd_sc_hs__tap_1 PHY_627 (  );
sky130_fd_sc_hs__tap_1 PHY_628 (  );
sky130_fd_sc_hs__tap_1 PHY_629 (  );
sky130_fd_sc_hs__tap_1 PHY_630 (  );
sky130_fd_sc_hs__tap_1 PHY_631 (  );
sky130_fd_sc_hs__tap_1 PHY_632 (  );
sky130_fd_sc_hs__tap_1 PHY_633 (  );
sky130_fd_sc_hs__tap_1 PHY_634 (  );
sky130_fd_sc_hs__tap_1 PHY_635 (  );
sky130_fd_sc_hs__tap_1 PHY_636 (  );
sky130_fd_sc_hs__tap_1 PHY_637 (  );
sky130_fd_sc_hs__tap_1 PHY_638 (  );
sky130_fd_sc_hs__tap_1 PHY_639 (  );
sky130_fd_sc_hs__tap_1 PHY_640 (  );
sky130_fd_sc_hs__tap_1 PHY_641 (  );
sky130_fd_sc_hs__tap_1 PHY_642 (  );
sky130_fd_sc_hs__tap_1 PHY_643 (  );
sky130_fd_sc_hs__tap_1 PHY_644 (  );
sky130_fd_sc_hs__tap_1 PHY_645 (  );
sky130_fd_sc_hs__tap_1 PHY_646 (  );
sky130_fd_sc_hs__tap_1 PHY_647 (  );
sky130_fd_sc_hs__tap_1 PHY_648 (  );
sky130_fd_sc_hs__tap_1 PHY_649 (  );
sky130_fd_sc_hs__tap_1 PHY_650 (  );
sky130_fd_sc_hs__tap_1 PHY_651 (  );
sky130_fd_sc_hs__tap_1 PHY_652 (  );
sky130_fd_sc_hs__tap_1 PHY_653 (  );
sky130_fd_sc_hs__tap_1 PHY_654 (  );
sky130_fd_sc_hs__tap_1 PHY_655 (  );
sky130_fd_sc_hs__tap_1 PHY_656 (  );
sky130_fd_sc_hs__tap_1 PHY_657 (  );
sky130_fd_sc_hs__tap_1 PHY_658 (  );
sky130_fd_sc_hs__tap_1 PHY_659 (  );
sky130_fd_sc_hs__tap_1 PHY_660 (  );
sky130_fd_sc_hs__tap_1 PHY_661 (  );
sky130_fd_sc_hs__tap_1 PHY_662 (  );
sky130_fd_sc_hs__tap_1 PHY_663 (  );
sky130_fd_sc_hs__tap_1 PHY_664 (  );
sky130_fd_sc_hs__tap_1 PHY_665 (  );
sky130_fd_sc_hs__tap_1 PHY_666 (  );
sky130_fd_sc_hs__tap_1 PHY_667 (  );
sky130_fd_sc_hs__tap_1 PHY_668 (  );
sky130_fd_sc_hs__tap_1 PHY_669 (  );
sky130_fd_sc_hs__tap_1 PHY_670 (  );
sky130_fd_sc_hs__tap_1 PHY_671 (  );
sky130_fd_sc_hs__tap_1 PHY_672 (  );
sky130_fd_sc_hs__tap_1 PHY_673 (  );
sky130_fd_sc_hs__tap_1 PHY_674 (  );
sky130_fd_sc_hs__tap_1 PHY_675 (  );
sky130_fd_sc_hs__tap_1 PHY_676 (  );
sky130_fd_sc_hs__tap_1 PHY_677 (  );
sky130_fd_sc_hs__tap_1 PHY_678 (  );
sky130_fd_sc_hs__tap_1 PHY_679 (  );
sky130_fd_sc_hs__tap_1 PHY_680 (  );
sky130_fd_sc_hs__tap_1 PHY_681 (  );
sky130_fd_sc_hs__tap_1 PHY_682 (  );
sky130_fd_sc_hs__tap_1 PHY_683 (  );
sky130_fd_sc_hs__tap_1 PHY_684 (  );
sky130_fd_sc_hs__tap_1 PHY_685 (  );
sky130_fd_sc_hs__tap_1 PHY_686 (  );
sky130_fd_sc_hs__tap_1 PHY_687 (  );
sky130_fd_sc_hs__tap_1 PHY_688 (  );
sky130_fd_sc_hs__tap_1 PHY_689 (  );
sky130_fd_sc_hs__tap_1 PHY_690 (  );
sky130_fd_sc_hs__tap_1 PHY_691 (  );
sky130_fd_sc_hs__tap_1 PHY_692 (  );
sky130_fd_sc_hs__tap_1 PHY_693 (  );
sky130_fd_sc_hs__tap_1 PHY_694 (  );
sky130_fd_sc_hs__tap_1 PHY_695 (  );
sky130_fd_sc_hs__tap_1 PHY_696 (  );
sky130_fd_sc_hs__tap_1 PHY_697 (  );
sky130_fd_sc_hs__tap_1 PHY_698 (  );
sky130_fd_sc_hs__tap_1 PHY_699 (  );
sky130_fd_sc_hs__tap_1 PHY_700 (  );
sky130_fd_sc_hs__tap_1 PHY_701 (  );
sky130_fd_sc_hs__tap_1 PHY_702 (  );
sky130_fd_sc_hs__tap_1 PHY_703 (  );
sky130_fd_sc_hs__tap_1 PHY_704 (  );
sky130_fd_sc_hs__tap_1 PHY_705 (  );
sky130_fd_sc_hs__tap_1 PHY_706 (  );
sky130_fd_sc_hs__tap_1 PHY_707 (  );
sky130_fd_sc_hs__tap_1 PHY_708 (  );
sky130_fd_sc_hs__tap_1 PHY_709 (  );
sky130_fd_sc_hs__tap_1 PHY_710 (  );
sky130_fd_sc_hs__tap_1 PHY_711 (  );
sky130_fd_sc_hs__tap_1 PHY_712 (  );
sky130_fd_sc_hs__tap_1 PHY_713 (  );
sky130_fd_sc_hs__tap_1 PHY_714 (  );
sky130_fd_sc_hs__tap_1 PHY_715 (  );
sky130_fd_sc_hs__tap_1 PHY_716 (  );
sky130_fd_sc_hs__tap_1 PHY_717 (  );
sky130_fd_sc_hs__tap_1 PHY_718 (  );
sky130_fd_sc_hs__tap_1 PHY_719 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_0 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_1 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_2 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_3 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_4 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_5 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_6 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_7 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_8 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_9 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_10 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_11 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_12 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_13 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_14 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_15 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_16 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_17 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_18 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_19 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_20 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_21 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_22 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_23 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_24 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_25 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_26 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_27 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_28 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_29 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_30 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_31 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_32 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_33 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_34 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_35 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_36 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_37 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_38 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_39 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_40 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_41 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_42 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_43 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_44 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_45 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_46 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_47 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_48 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_49 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_50 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_51 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_52 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_53 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_54 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_55 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_56 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_57 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_58 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_59 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_60 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_61 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_62 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_63 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_64 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_65 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_66 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_67 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_68 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_69 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_70 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_71 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_72 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_73 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_74 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_75 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_76 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_77 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_78 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_79 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_80 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_81 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_82 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_83 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_84 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_85 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_86 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_87 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_88 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_89 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_90 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_91 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_92 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_93 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_94 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_95 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_96 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_97 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_98 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_99 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_100 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_101 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_102 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_103 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_104 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_105 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_106 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_107 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_108 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_109 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_110 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_111 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_112 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_113 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_114 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_115 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_116 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_117 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_118 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_119 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_120 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_121 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_122 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_123 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_124 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_125 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_126 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_127 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_128 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_129 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_130 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_131 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_132 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_133 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_134 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_135 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_136 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_137 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_138 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_139 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_140 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_141 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_142 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_143 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_144 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_145 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_146 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_147 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_148 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_149 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_150 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_151 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_152 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_153 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_154 (  );
sky130_fd_sc_hs__fill_1 ENDCAP_155 (  );
sky130_fd_sc_hs__buf_1 clk_86_buf ( .A(clk_61 ), .X(clk_86 ) );
sky130_fd_sc_hs__buf_1 clk_85_buf ( .A(clk_60 ), .X(clk_85 ) );
sky130_fd_sc_hs__buf_1 clk_84_buf ( .A(clk_59 ), .X(clk_84 ) );
sky130_fd_sc_hs__buf_1 clk_83_buf ( .A(clk_59 ), .X(clk_83 ) );
sky130_fd_sc_hs__buf_1 clk_82_buf ( .A(clk_56 ), .X(clk_82 ) );
sky130_fd_sc_hs__buf_1 clk_81_buf ( .A(clk_55 ), .X(clk_81 ) );
sky130_fd_sc_hs__buf_1 clk_80_buf ( .A(clk_55 ), .X(clk_80 ) );
sky130_fd_sc_hs__buf_1 clk_79_buf ( .A(clk_54 ), .X(clk_79 ) );
sky130_fd_sc_hs__buf_1 clk_78_buf ( .A(clk_54 ), .X(clk_78 ) );
sky130_fd_sc_hs__buf_1 clk_77_buf ( .A(clk_53 ), .X(clk_77 ) );
sky130_fd_sc_hs__buf_1 clk_76_buf ( .A(clk_52 ), .X(clk_76 ) );
sky130_fd_sc_hs__buf_1 clk_75_buf ( .A(clk_51 ), .X(clk_75 ) );
sky130_fd_sc_hs__buf_1 clk_74_buf ( .A(clk_51 ), .X(clk_74 ) );
sky130_fd_sc_hs__buf_1 clk_73_buf ( .A(clk_50 ), .X(clk_73 ) );
sky130_fd_sc_hs__buf_1 clk_72_buf ( .A(clk_50 ), .X(clk_72 ) );
sky130_fd_sc_hs__buf_1 clk_71_buf ( .A(clk_49 ), .X(clk_71 ) );
sky130_fd_sc_hs__buf_1 clk_70_buf ( .A(clk_49 ), .X(clk_70 ) );
sky130_fd_sc_hs__buf_1 clk_69_buf ( .A(clk_48 ), .X(clk_69 ) );
sky130_fd_sc_hs__buf_1 clk_68_buf ( .A(clk_48 ), .X(clk_68 ) );
sky130_fd_sc_hs__buf_1 clk_67_buf ( .A(clk_47 ), .X(clk_67 ) );
sky130_fd_sc_hs__buf_1 clk_66_buf ( .A(clk_47 ), .X(clk_66 ) );
sky130_fd_sc_hs__buf_1 clk_65_buf ( .A(clk_46 ), .X(clk_65 ) );
sky130_fd_sc_hs__buf_1 clk_64_buf ( .A(clk_46 ), .X(clk_64 ) );
sky130_fd_sc_hs__buf_1 clk_63_buf ( .A(clk_45 ), .X(clk_63 ) );
sky130_fd_sc_hs__buf_1 clk_62_buf ( .A(clk_44 ), .X(clk_62 ) );
sky130_fd_sc_hs__buf_1 clk_61_buf ( .A(clk_43 ), .X(clk_61 ) );
sky130_fd_sc_hs__buf_1 clk_60_buf ( .A(clk_43 ), .X(clk_60 ) );
sky130_fd_sc_hs__buf_1 clk_59_buf ( .A(clk_42 ), .X(clk_59 ) );
sky130_fd_sc_hs__buf_1 clk_58_buf ( .A(clk_41 ), .X(clk_58 ) );
sky130_fd_sc_hs__buf_1 clk_57_buf ( .A(clk_40 ), .X(clk_57 ) );
sky130_fd_sc_hs__buf_1 clk_56_buf ( .A(clk_39 ), .X(clk_56 ) );
sky130_fd_sc_hs__buf_1 clk_55_buf ( .A(clk_38 ), .X(clk_55 ) );
sky130_fd_sc_hs__buf_1 clk_54_buf ( .A(clk_37 ), .X(clk_54 ) );
sky130_fd_sc_hs__buf_1 clk_53_buf ( .A(clk_36 ), .X(clk_53 ) );
sky130_fd_sc_hs__buf_1 clk_52_buf ( .A(clk_36 ), .X(clk_52 ) );
sky130_fd_sc_hs__buf_1 clk_51_buf ( .A(clk_35 ), .X(clk_51 ) );
sky130_fd_sc_hs__buf_1 clk_50_buf ( .A(clk_35 ), .X(clk_50 ) );
sky130_fd_sc_hs__buf_1 clk_49_buf ( .A(clk_34 ), .X(clk_49 ) );
sky130_fd_sc_hs__buf_1 clk_48_buf ( .A(clk_34 ), .X(clk_48 ) );
sky130_fd_sc_hs__buf_1 clk_47_buf ( .A(clk_33 ), .X(clk_47 ) );
sky130_fd_sc_hs__buf_1 clk_46_buf ( .A(clk_33 ), .X(clk_46 ) );
sky130_fd_sc_hs__buf_1 clk_45_buf ( .A(clk_32 ), .X(clk_45 ) );
sky130_fd_sc_hs__buf_1 clk_44_buf ( .A(clk_32 ), .X(clk_44 ) );
sky130_fd_sc_hs__buf_1 clk_43_buf ( .A(clk_31 ), .X(clk_43 ) );
sky130_fd_sc_hs__buf_1 clk_42_buf ( .A(clk_30 ), .X(clk_42 ) );
sky130_fd_sc_hs__buf_1 clk_41_buf ( .A(clk_29 ), .X(clk_41 ) );
sky130_fd_sc_hs__buf_1 clk_40_buf ( .A(clk_29 ), .X(clk_40 ) );
sky130_fd_sc_hs__buf_1 clk_39_buf ( .A(clk_28 ), .X(clk_39 ) );
sky130_fd_sc_hs__buf_1 clk_38_buf ( .A(clk_27 ), .X(clk_38 ) );
sky130_fd_sc_hs__buf_1 clk_37_buf ( .A(clk_27 ), .X(clk_37 ) );
sky130_fd_sc_hs__buf_1 clk_36_buf ( .A(clk_26 ), .X(clk_36 ) );
sky130_fd_sc_hs__buf_1 clk_35_buf ( .A(clk_25 ), .X(clk_35 ) );
sky130_fd_sc_hs__buf_1 clk_34_buf ( .A(clk_24 ), .X(clk_34 ) );
sky130_fd_sc_hs__buf_1 clk_33_buf ( .A(clk_23 ), .X(clk_33 ) );
sky130_fd_sc_hs__buf_1 clk_32_buf ( .A(clk_22 ), .X(clk_32 ) );
sky130_fd_sc_hs__buf_1 clk_31_buf ( .A(clk_21 ), .X(clk_31 ) );
sky130_fd_sc_hs__buf_1 clk_30_buf ( .A(clk_20 ), .X(clk_30 ) );
sky130_fd_sc_hs__buf_1 clk_29_buf ( .A(clk_19 ), .X(clk_29 ) );
sky130_fd_sc_hs__buf_1 clk_28_buf ( .A(clk_18 ), .X(clk_28 ) );
sky130_fd_sc_hs__buf_1 clk_27_buf ( .A(clk_17 ), .X(clk_27 ) );
sky130_fd_sc_hs__buf_1 clk_26_buf ( .A(clk_17 ), .X(clk_26 ) );
sky130_fd_sc_hs__buf_1 clk_25_buf ( .A(clk_16 ), .X(clk_25 ) );
sky130_fd_sc_hs__buf_1 clk_24_buf ( .A(clk_16 ), .X(clk_24 ) );
sky130_fd_sc_hs__buf_1 clk_23_buf ( .A(clk_15 ), .X(clk_23 ) );
sky130_fd_sc_hs__buf_1 clk_22_buf ( .A(clk_15 ), .X(clk_22 ) );
sky130_fd_sc_hs__buf_1 clk_21_buf ( .A(clk_14 ), .X(clk_21 ) );
sky130_fd_sc_hs__buf_1 clk_20_buf ( .A(clk_14 ), .X(clk_20 ) );
sky130_fd_sc_hs__buf_1 clk_19_buf ( .A(clk_13 ), .X(clk_19 ) );
sky130_fd_sc_hs__buf_1 clk_18_buf ( .A(clk_13 ), .X(clk_18 ) );
sky130_fd_sc_hs__buf_1 clk_17_buf ( .A(clk_12 ), .X(clk_17 ) );
sky130_fd_sc_hs__buf_1 clk_16_buf ( .A(clk_11 ), .X(clk_16 ) );
sky130_fd_sc_hs__buf_1 clk_15_buf ( .A(clk_10 ), .X(clk_15 ) );
sky130_fd_sc_hs__buf_1 clk_14_buf ( .A(clk_9 ), .X(clk_14 ) );
sky130_fd_sc_hs__buf_1 clk_13_buf ( .A(clk_8 ), .X(clk_13 ) );
sky130_fd_sc_hs__buf_1 clk_12_buf ( .A(clk_7 ), .X(clk_12 ) );
sky130_fd_sc_hs__buf_1 clk_11_buf ( .A(clk_6 ), .X(clk_11 ) );
sky130_fd_sc_hs__buf_1 clk_10_buf ( .A(clk_6 ), .X(clk_10 ) );
sky130_fd_sc_hs__buf_1 clk_9_buf ( .A(clk_5 ), .X(clk_9 ) );
sky130_fd_sc_hs__buf_1 clk_8_buf ( .A(clk_5 ), .X(clk_8 ) );
sky130_fd_sc_hs__buf_1 clk_7_buf ( .A(clk_4 ), .X(clk_7 ) );
sky130_fd_sc_hs__buf_1 clk_6_buf ( .A(clk_3 ), .X(clk_6 ) );
sky130_fd_sc_hs__buf_1 clk_5_buf ( .A(clk_2 ), .X(clk_5 ) );
sky130_fd_sc_hs__buf_1 clk_4_buf ( .A(clk_2 ), .X(clk_4 ) );
sky130_fd_sc_hs__buf_1 clk_3_buf ( .A(clk_1 ), .X(clk_3 ) );
sky130_fd_sc_hs__buf_1 clk_2_buf ( .A(clk_0 ), .X(clk_2 ) );
sky130_fd_sc_hs__buf_1 clk_1_buf ( .A(clk_0 ), .X(clk_1 ) );
sky130_fd_sc_hs__buf_1 clk_0_buf ( .A(clk ), .X(clk_0 ) );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_0 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_8 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_9 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_10 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_11 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_12 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_13 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_14 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_15 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_16 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_17 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_18 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_19 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_20 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_21 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_22 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_23 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_24 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_25 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_26 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_27 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_28 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_29 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_30 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_31 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_32 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_33 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_34 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_35 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_36 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_37 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_38 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_39 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_40 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_41 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_42 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_43 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_44 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_45 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_46 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_47 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_48 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_49 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_50 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_51 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_52 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_53 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_54 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_55 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_56 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_57 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_58 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_59 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_60 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_61 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_62 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_63 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_64 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_65 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_66 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_67 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_68 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_69 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_70 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_71 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_72 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_73 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_74 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_75 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_76 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_77 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_78 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_79 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_80 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_81 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_82 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_83 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_84 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_85 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_86 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_87 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_88 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_89 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_90 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_91 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_92 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_93 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_94 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_95 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_96 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_97 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_98 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_99 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_100 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_101 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_102 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_103 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_104 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_105 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_106 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_107 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_108 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_109 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_110 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_111 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_112 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_113 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_114 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_115 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_116 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_117 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_118 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_119 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_120 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_121 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_122 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_123 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_124 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_125 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_126 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_127 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_128 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_129 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_130 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_131 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_132 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_133 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_134 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_135 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_136 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_137 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_138 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_139 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_140 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_141 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_142 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_143 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_144 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_145 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_146 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_147 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_148 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_149 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_150 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_151 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_152 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_153 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_154 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_155 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_156 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_157 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_158 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_159 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_160 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_161 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_162 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_163 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_164 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_165 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_166 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_167 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_168 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_169 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_170 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_171 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_172 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_173 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_174 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_175 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_176 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_177 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_178 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_179 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_180 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_181 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_182 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_183 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_184 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_185 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_186 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_187 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_188 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_189 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_190 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_191 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_192 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_193 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_194 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_195 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_196 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_197 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_198 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_199 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_200 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_201 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_202 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_203 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_204 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_205 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_206 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_207 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_208 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_209 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_210 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_211 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_212 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_213 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_214 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_215 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_216 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_217 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_218 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_219 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_220 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_221 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_222 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_223 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_224 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_225 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_226 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_227 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_228 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_229 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_230 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_231 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_232 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_233 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_234 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_235 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_236 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_237 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_238 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_239 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_240 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_241 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_242 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_243 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_244 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_245 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_246 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_247 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_248 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_249 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_250 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_251 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_252 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_253 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_254 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_255 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_256 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_257 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_258 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_259 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_260 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_261 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_262 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_263 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_264 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_265 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_266 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_267 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_268 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_269 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_270 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_271 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_272 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_273 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_274 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_275 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_276 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_277 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_278 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_279 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_280 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_281 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_282 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_283 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_284 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_285 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_286 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_287 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_288 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_289 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_290 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_291 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_292 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_293 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_294 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_295 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_296 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_297 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_298 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_299 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_300 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_301 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_302 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_303 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_304 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_305 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_306 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_307 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_308 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_309 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_310 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_311 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_312 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_313 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_314 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_315 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_316 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_317 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_318 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_319 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_320 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_321 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_322 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_323 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_324 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_325 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_326 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_327 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_328 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_329 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_330 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_331 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_332 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_333 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_334 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_335 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_336 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_337 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_338 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_339 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_340 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_341 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_342 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_343 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_344 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_345 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_346 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_347 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_348 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_349 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_350 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_351 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_352 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_353 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_354 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_355 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_356 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_357 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_358 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_359 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_360 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_361 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_362 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_363 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_364 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_365 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_366 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_367 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_368 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_369 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_370 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_371 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_372 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_373 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_374 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_375 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_376 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_377 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_378 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_379 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_380 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_381 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_382 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_383 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_384 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_385 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_386 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_387 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_388 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_389 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_390 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_391 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_392 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_393 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_394 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_395 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_396 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_397 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_398 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_399 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_400 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_401 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_402 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_403 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_404 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_405 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_406 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_407 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_408 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_409 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_410 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_411 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_412 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_413 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_414 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_415 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_416 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_417 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_418 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_419 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_420 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_421 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_422 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_423 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_424 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_425 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_426 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_427 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_428 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_429 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_430 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_431 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_432 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_433 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_434 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_435 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_436 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_437 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_438 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_439 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_440 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_441 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_442 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_443 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_444 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_445 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_446 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_447 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_448 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_449 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_450 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_451 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_452 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_453 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_454 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_455 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_456 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_457 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_458 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_459 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_460 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_461 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_462 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_463 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_464 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_465 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_466 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_467 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_468 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_469 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_470 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_471 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_472 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_473 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_474 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_475 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_476 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_477 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_478 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_479 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_480 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_481 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_482 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_483 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_484 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_485 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_486 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_487 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_488 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_489 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_490 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_491 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_492 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_493 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_494 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_495 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_496 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_497 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_498 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_499 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_500 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_501 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_502 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_503 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_504 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_505 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_506 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_507 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_508 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_509 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_510 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_511 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_512 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_513 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_514 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_515 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_516 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_517 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_518 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_519 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_520 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_521 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_522 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_523 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_524 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_525 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_526 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_527 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_528 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_529 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_530 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_531 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_532 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_533 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_534 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_535 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_536 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_537 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_538 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_539 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_540 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_541 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_542 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_543 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_544 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_545 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_546 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_547 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_548 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_549 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_550 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_551 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_552 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_553 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_554 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_555 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_556 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_557 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_558 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_559 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_560 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_561 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_562 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_563 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_564 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_565 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_566 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_567 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_568 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_569 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_570 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_571 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_572 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_573 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_574 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_575 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_576 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_577 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_578 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_579 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_580 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_581 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_582 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_583 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_584 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_585 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_586 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_587 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_588 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_589 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_590 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_591 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_592 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_593 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_594 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_595 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_596 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_597 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_598 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_599 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_600 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_601 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_602 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_603 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_604 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_605 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_606 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_607 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_608 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_609 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_610 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_611 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_612 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_613 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_614 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_615 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_616 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_617 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_618 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_619 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_620 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_621 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_622 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_623 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_624 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_625 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_626 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_627 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_628 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_629 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_630 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_631 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_632 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_633 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_634 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_635 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_636 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_637 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_638 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_639 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_640 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_641 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_642 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_643 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_644 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_645 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_646 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_647 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_648 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_649 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_650 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_651 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_652 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_653 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_654 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_655 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_656 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_657 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_658 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_659 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_660 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_661 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_662 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_663 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_664 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_665 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_666 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_667 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_668 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_669 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_670 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_671 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_672 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_673 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_674 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_675 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_676 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_677 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_678 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_679 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_680 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_681 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_682 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_683 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_684 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_685 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_686 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_687 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_688 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_689 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_690 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_691 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_692 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_693 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_694 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_695 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_696 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_697 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_698 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_699 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_700 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_701 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_702 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_703 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_704 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_705 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_706 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_707 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_708 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_709 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_710 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_711 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_712 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_713 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_714 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_715 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_716 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_717 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_718 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_719 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_720 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_721 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_722 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_723 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_724 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_725 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_726 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_727 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_728 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_729 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_730 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_731 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_732 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_733 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_734 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_735 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_736 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_737 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_738 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_739 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_740 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_741 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_742 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_743 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_744 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_745 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_746 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_747 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_748 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_749 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_750 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_751 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_752 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_753 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_754 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_755 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_756 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_757 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_758 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_759 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_760 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_761 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_762 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_763 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_764 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_765 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_766 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_767 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_768 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_769 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_770 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_771 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_772 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_773 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_774 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_775 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_776 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_777 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_778 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_779 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_780 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_781 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_782 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_783 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_784 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_785 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_786 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_787 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_788 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_789 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_790 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_791 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_792 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_793 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_794 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_795 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_796 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_797 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_798 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_799 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_800 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_801 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_802 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_803 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_804 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_805 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_806 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_807 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_808 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_809 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_810 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_811 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_812 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_813 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_814 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_815 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_816 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_817 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_818 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_819 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_820 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_821 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_822 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_823 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_824 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_825 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_826 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_827 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_828 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_829 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_830 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_831 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_832 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_833 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_834 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_835 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_836 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_837 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_838 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_839 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_840 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_841 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_842 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_843 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_844 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_845 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_846 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_847 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_848 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_849 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_850 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_851 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_852 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_853 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_854 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_855 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_856 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_857 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_858 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_859 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_860 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_861 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_862 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_863 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_864 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_865 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_866 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_867 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_868 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_869 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_870 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_871 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_872 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_873 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_874 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_875 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_876 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_877 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_878 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_879 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_880 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_881 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_882 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_883 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_884 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_885 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_886 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_887 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_888 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_889 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_890 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_891 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_892 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_893 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_894 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_895 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_896 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_897 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_898 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_899 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_900 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_901 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_902 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_903 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_904 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_905 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_906 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_907 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_908 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_909 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_910 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_911 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_912 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_913 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_914 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_915 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_916 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_917 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_918 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_919 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_920 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_921 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_922 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_923 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_924 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_925 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_926 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_927 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_928 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_929 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_930 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_931 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_932 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_933 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_934 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_935 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_936 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_937 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_938 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_939 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_940 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_941 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_942 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_943 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_944 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_945 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_946 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_947 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_948 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_949 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_950 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_951 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_952 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_953 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_954 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_955 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_956 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_957 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_958 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_959 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_960 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_961 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_962 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_963 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_964 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_965 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_966 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_967 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_968 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_969 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_970 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_971 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_972 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_973 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_974 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_975 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_976 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_977 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_978 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_979 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_980 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_981 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_982 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_983 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_984 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_985 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_986 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_987 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_988 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_989 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_990 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_991 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_992 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_993 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_994 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_995 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_996 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_997 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_998 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_999 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1000 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1001 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1002 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1003 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1004 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1005 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1006 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1007 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1008 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1009 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1010 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1011 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1012 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1013 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1014 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1015 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1016 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1017 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1018 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1019 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1020 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1021 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1022 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1023 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1024 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1025 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1026 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1027 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1028 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1029 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1030 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1031 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1032 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1033 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1034 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1035 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1036 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1037 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1038 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1039 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1040 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1041 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1042 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1043 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1044 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1045 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1046 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1047 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1048 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1049 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1050 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1051 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1052 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1053 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1054 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1055 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1056 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1057 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1058 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1059 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1060 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1061 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1062 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1063 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1064 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1065 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1066 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1067 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1068 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1069 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1070 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1071 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1072 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1073 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1074 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1075 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1076 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1077 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1078 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1079 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1080 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1081 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1082 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1083 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1084 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1085 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1086 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1087 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1088 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1089 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1090 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1091 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1092 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1093 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1094 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1095 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1096 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1097 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1098 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1099 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1100 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1101 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1102 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1103 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1104 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1105 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1106 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1107 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1108 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1109 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1110 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1111 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1112 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1113 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1114 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1115 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1116 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1117 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1118 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1119 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1120 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1121 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1122 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1123 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1124 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1125 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1126 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1127 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1128 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1129 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1130 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1131 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1132 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1133 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1134 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1135 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1136 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1137 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1138 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1139 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1140 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1141 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1142 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1143 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1144 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1145 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1146 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1147 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1148 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1149 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1150 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1151 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1152 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1153 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1154 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1155 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1156 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1157 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1158 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1159 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1160 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1161 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1162 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1163 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1164 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1165 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1166 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1167 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1168 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1169 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1170 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1171 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1172 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1173 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1174 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1175 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1176 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1177 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1178 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1179 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1180 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1181 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1182 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1183 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1184 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1185 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1186 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1187 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1188 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1189 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1190 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1191 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1192 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1193 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1194 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1195 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1196 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1197 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1198 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1199 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1200 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1201 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1202 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1203 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1204 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1205 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1206 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1207 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1208 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1209 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1210 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1211 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1212 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1213 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1214 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1215 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1216 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1217 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1218 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1219 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1220 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1221 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1222 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1223 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1224 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1225 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1226 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1227 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1228 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1229 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1230 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1231 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1232 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1233 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1234 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1235 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1236 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1237 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1238 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1239 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1240 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1241 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1242 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1243 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1244 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1245 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1246 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1247 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1248 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1249 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1250 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1251 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1252 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1253 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1254 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1255 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1256 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1257 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1258 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1259 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1260 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1261 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1262 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1263 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1264 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1265 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1266 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1267 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1268 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1269 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1270 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1271 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1272 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1273 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1274 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1275 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1276 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1277 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1278 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1279 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1280 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1281 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1282 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1283 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1284 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1285 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1286 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1287 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1288 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1289 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1290 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1291 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1292 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1293 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1294 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1295 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1296 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1297 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1298 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1299 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1300 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1301 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1302 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1303 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1304 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1305 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1306 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1307 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1308 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1309 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1310 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1311 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1312 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1313 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1314 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1315 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1316 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1317 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1318 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1319 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1320 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1321 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1322 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1323 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1324 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1325 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1326 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1327 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1328 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1329 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1330 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1331 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1332 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1333 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1334 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1335 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1336 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1337 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1338 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1339 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1340 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1341 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1342 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1343 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1344 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1345 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1346 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1347 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1348 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1349 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1350 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1351 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1352 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1353 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1354 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1355 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1356 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1357 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1358 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1359 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1360 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1361 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1362 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1363 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1364 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1365 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1366 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1367 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1368 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1369 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1370 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1371 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1372 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1373 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1374 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1375 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1376 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1377 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1378 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1379 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1380 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1381 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1382 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1383 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1384 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1385 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1386 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1387 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1388 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1389 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1390 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1391 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1392 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1393 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1394 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1395 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1396 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1397 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1398 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1399 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1400 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1401 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1402 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1403 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1404 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1405 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1406 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1407 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1408 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1409 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1410 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1411 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1412 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1413 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1414 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1415 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1416 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1417 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1418 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1419 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1420 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1421 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1422 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1423 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1424 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1425 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1426 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1427 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1428 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1429 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1430 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1431 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1432 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1433 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1434 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1435 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1436 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1437 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1438 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1439 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1440 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1441 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1442 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1443 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1444 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1445 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1446 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1447 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1448 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1449 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1450 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1451 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1452 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1453 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1454 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1455 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1456 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1457 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1458 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1459 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1460 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1461 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1462 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1463 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1464 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1465 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1466 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1467 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1468 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1469 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1470 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1471 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1472 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1473 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1474 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1475 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1476 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1477 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1478 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1479 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1480 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1481 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1482 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1483 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1484 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1485 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1486 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1487 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1488 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1489 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1490 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1491 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1492 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1493 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1494 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1495 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1496 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1497 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1498 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1499 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1500 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1501 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1502 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1503 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1504 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1505 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1506 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1507 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1508 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1509 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1510 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1511 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1512 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1513 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1514 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1515 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1516 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1517 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1518 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1519 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1520 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1521 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1522 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1523 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1524 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1525 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1526 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1527 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1528 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1529 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1530 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1531 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1532 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1533 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1534 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1535 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1536 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1537 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1538 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1539 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1540 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1541 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1542 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1543 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1544 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1545 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1546 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1547 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1548 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1549 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1550 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1551 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1552 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1553 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1554 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1555 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1556 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1557 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1558 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1559 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1560 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1561 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1562 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1563 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1564 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1565 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1566 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1567 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1568 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1569 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1570 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1571 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1572 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1573 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1574 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1575 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1576 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1577 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1578 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1579 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1580 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1581 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1582 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1583 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1584 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1585 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1586 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1587 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1588 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1589 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1590 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1591 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1592 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1593 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1594 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1595 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1596 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1597 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1598 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1599 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1600 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1601 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1602 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1603 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1604 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1605 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1606 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1607 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1608 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1609 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1610 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1611 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1612 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1613 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1614 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1615 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1616 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1617 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1618 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1619 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1620 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1621 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1622 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1623 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1624 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1625 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1626 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1627 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1628 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1629 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1630 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1631 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1632 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1633 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1634 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1635 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1636 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1637 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1638 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1639 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1640 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1641 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1642 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1643 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1644 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1645 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1646 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1647 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1648 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1649 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1650 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1651 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1652 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1653 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1654 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1655 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1656 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1657 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1658 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1659 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1660 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1661 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1662 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1663 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1664 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1665 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1666 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1667 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1668 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1669 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1670 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1671 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1672 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1673 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1674 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1675 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1676 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1677 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1678 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1679 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1680 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1681 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1682 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1683 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1684 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1685 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1686 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1687 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1688 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1689 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1690 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1691 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1692 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1693 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1694 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1695 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1696 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1697 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1698 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1699 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1700 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1701 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1702 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1703 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1704 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1705 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1706 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1707 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1708 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1709 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1710 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1711 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1712 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1713 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1714 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1715 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1716 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1717 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1718 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1719 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1720 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1721 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1722 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1723 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1724 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1725 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1726 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1727 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1728 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1729 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1730 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1731 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1732 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1733 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1734 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1735 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1736 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1737 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1738 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1739 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1740 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1741 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1742 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1743 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1744 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1745 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1746 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1747 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1748 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1749 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1750 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1751 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1752 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1753 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1754 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1755 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1756 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1757 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1758 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1759 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1760 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1761 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1762 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1763 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1764 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1765 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1766 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1767 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1768 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1769 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1770 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1771 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1772 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1773 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1774 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1775 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1776 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1777 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1778 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1779 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1780 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1781 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1782 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1783 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1784 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1785 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1786 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1787 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1788 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1789 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1790 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1791 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1792 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1793 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1794 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1795 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1796 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1797 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1798 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1799 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1800 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1801 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1802 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1803 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1804 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1805 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1806 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1807 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1808 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1809 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1810 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1811 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1812 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1813 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1814 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1815 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1816 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1817 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1818 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1819 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1820 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1821 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1822 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1823 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1824 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1825 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1826 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1827 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1828 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1829 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1830 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1831 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1832 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1833 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1834 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1835 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1836 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1837 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1838 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1839 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1840 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1841 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1842 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1843 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1844 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1845 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1846 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1847 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1848 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1849 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1850 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1851 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1852 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1853 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1854 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1855 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1856 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1857 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1858 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1859 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1860 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1861 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1862 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1863 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1864 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1865 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1866 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1867 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1868 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1869 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1870 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1871 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1872 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1873 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1874 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1875 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1876 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1877 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1878 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1879 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1880 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1881 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1882 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1883 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1884 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1885 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1886 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1887 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1888 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1889 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1890 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1891 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1892 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1893 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1894 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1895 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1896 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1897 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1898 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1899 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1900 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1901 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1902 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1903 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1904 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1905 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1906 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1907 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1908 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1909 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1910 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1911 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1912 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1913 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1914 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1915 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1916 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1917 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1918 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1919 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1920 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1921 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1922 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1923 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1924 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1925 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1926 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1927 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1928 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1929 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1930 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1931 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1932 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1933 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1934 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1935 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1936 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1937 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1938 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1939 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1940 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1941 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1942 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1943 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1944 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1945 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1946 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1947 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1948 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1949 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1950 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1951 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1952 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1953 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1954 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1955 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1956 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1957 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1958 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1959 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1960 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1961 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1962 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1963 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1964 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1965 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1966 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1967 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1968 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1969 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1970 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1971 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1972 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1973 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1974 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1975 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1976 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1977 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1978 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1979 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1980 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1981 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1982 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1983 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1984 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1985 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1986 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1987 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1988 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1989 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1990 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1991 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1992 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1993 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1994 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1995 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_1996 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_1997 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_1998 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_1999 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2000 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2001 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2002 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2003 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2004 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2005 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2006 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2007 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2008 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2009 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2010 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2011 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2012 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2013 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2014 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2015 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2016 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2017 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2018 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2019 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2020 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2021 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2022 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2023 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2024 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2025 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2026 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2027 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2028 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2029 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2030 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2031 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2032 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2033 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2034 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2035 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2036 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2037 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2038 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2039 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2040 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2041 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2042 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2043 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2044 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2045 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2046 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2047 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2048 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2049 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2050 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2051 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2052 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2053 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2054 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2055 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2056 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2057 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2058 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2059 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2060 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2061 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2062 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2063 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2064 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2065 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2066 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2067 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2068 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2069 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2070 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2071 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2072 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2073 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2074 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2075 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2076 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2077 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2078 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2079 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2080 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2081 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2082 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2083 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2084 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2085 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2086 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2087 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2088 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2089 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2090 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2091 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2092 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2093 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2094 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2095 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2096 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2097 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2098 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2099 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2100 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2101 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2102 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2103 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2104 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2105 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2106 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2107 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2108 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2109 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2110 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2111 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2112 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2113 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2114 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2115 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2116 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2117 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2118 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2119 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2120 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2121 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2122 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2123 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2124 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2125 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2126 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2127 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2128 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2129 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2130 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2131 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2132 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2133 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2134 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2135 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2136 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2137 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2138 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2139 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2140 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2141 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2142 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2143 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2144 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2145 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2146 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2147 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2148 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2149 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2150 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2151 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2152 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2153 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2154 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2155 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2156 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2157 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2158 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2159 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2160 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2161 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2162 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2163 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2164 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2165 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2166 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2167 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2168 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2169 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2170 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2171 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2172 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2173 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2174 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2175 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2176 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2177 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2178 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2179 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2180 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2181 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2182 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2183 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2184 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2185 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2186 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2187 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2188 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2189 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2190 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2191 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2192 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2193 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2194 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2195 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2196 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2197 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2198 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2199 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2200 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2201 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2202 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2203 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2204 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2205 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2206 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2207 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2208 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2209 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2210 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2211 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2212 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2213 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2214 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2215 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2216 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2217 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2218 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2219 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2220 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2221 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2222 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2223 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2224 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2225 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2226 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2227 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2228 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2229 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2230 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2231 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2232 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2233 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2234 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2235 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2236 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2237 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2238 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2239 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2240 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2241 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2242 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2243 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2244 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2245 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2246 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2247 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2248 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2249 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2250 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2251 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2252 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2253 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2254 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2255 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2256 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2257 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2258 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2259 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2260 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2261 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2262 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2263 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2264 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2265 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2266 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2267 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2268 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2269 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2270 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2271 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2272 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2273 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2274 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2275 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2276 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2277 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2278 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2279 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2280 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2281 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2282 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2283 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2284 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2285 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2286 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2287 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2288 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2289 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2290 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2291 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2292 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2293 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2294 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2295 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2296 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2297 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2298 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2299 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2300 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2301 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2302 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2303 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2304 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2305 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2306 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2307 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2308 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2309 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2310 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2311 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2312 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2313 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2314 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2315 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2316 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2317 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2318 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2319 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2320 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2321 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2322 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2323 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2324 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2325 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2326 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2327 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2328 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2329 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2330 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2331 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2332 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2333 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2334 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2335 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2336 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2337 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2338 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2339 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2340 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2341 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2342 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2343 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2344 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2345 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2346 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2347 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2348 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2349 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2350 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2351 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2352 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2353 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2354 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2355 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2356 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2357 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2358 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2359 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2360 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2361 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2362 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2363 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2364 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2365 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2366 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2367 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2368 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2369 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2370 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2371 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2372 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2373 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2374 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2375 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2376 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2377 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2378 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2379 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2380 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2381 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2382 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2383 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2384 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2385 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2386 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2387 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2388 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2389 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2390 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2391 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2392 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2393 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2394 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2395 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2396 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2397 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2398 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2399 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2400 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2401 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2402 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2403 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2404 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2405 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2406 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2407 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2408 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2409 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2410 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2411 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2412 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2413 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2414 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2415 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2416 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2417 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2418 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2419 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2420 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2421 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2422 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2423 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2424 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2425 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2426 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2427 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2428 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2429 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2430 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2431 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2432 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2433 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2434 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2435 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2436 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2437 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2438 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2439 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2440 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2441 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2442 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2443 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2444 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2445 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2446 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2447 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2448 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2449 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2450 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2451 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2452 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2453 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2454 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2455 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2456 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2457 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2458 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2459 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2460 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2461 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2462 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2463 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2464 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2465 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2466 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2467 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2468 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2469 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2470 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2471 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2472 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2473 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2474 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2475 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2476 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2477 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2478 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2479 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2480 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2481 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2482 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2483 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2484 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2485 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2486 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2487 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2488 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2489 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2490 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2491 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2492 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2493 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2494 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2495 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2496 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2497 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2498 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2499 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2500 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2501 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2502 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2503 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2504 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2505 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2506 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2507 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2508 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2509 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2510 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2511 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2512 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2513 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2514 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2515 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2516 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2517 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2518 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2519 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2520 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2521 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2522 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2523 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2524 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2525 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2526 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2527 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2528 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2529 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2530 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2531 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2532 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2533 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2534 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2535 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2536 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2537 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2538 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2539 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2540 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2541 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2542 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2543 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2544 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2545 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2546 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2547 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2548 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2549 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2550 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2551 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2552 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2553 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2554 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2555 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2556 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2557 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2558 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2559 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2560 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2561 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2562 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2563 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2564 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2565 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2566 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2567 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2568 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2569 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2570 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2571 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2572 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2573 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2574 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2575 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2576 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2577 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2578 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2579 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2580 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2581 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2582 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2583 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2584 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2585 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2586 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2587 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2588 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2589 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2590 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2591 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2592 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2593 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2594 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2595 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2596 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2597 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2598 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2599 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2600 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2601 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2602 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2603 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2604 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2605 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2606 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2607 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2608 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2609 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2610 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2611 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2612 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2613 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2614 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2615 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2616 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2617 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2618 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2619 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2620 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2621 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2622 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2623 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2624 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2625 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2626 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2627 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2628 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2629 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2630 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2631 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2632 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2633 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2634 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2635 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2636 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2637 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2638 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2639 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2640 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2641 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2642 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2643 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2644 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2645 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2646 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2647 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2648 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2649 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2650 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2651 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2652 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2653 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2654 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2655 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2656 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2657 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2658 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2659 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2660 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2661 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2662 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2663 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2664 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2665 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2666 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2667 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2668 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2669 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2670 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2671 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2672 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2673 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2674 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2675 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2676 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2677 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2678 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2679 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2680 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2681 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2682 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2683 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2684 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2685 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2686 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2687 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2688 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2689 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2690 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2691 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2692 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2693 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2694 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2695 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2696 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2697 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2698 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2699 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2700 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2701 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2702 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2703 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2704 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2705 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2706 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2707 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2708 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2709 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2710 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2711 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2712 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2713 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2714 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2715 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2716 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2717 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2718 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2719 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2720 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2721 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2722 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2723 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2724 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2725 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2726 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2727 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2728 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2729 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2730 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2731 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2732 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2733 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2734 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2735 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2736 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2737 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2738 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2739 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2740 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2741 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2742 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2743 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2744 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2745 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2746 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2747 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2748 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2749 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2750 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2751 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2752 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2753 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2754 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2755 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2756 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2757 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2758 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2759 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2760 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2761 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2762 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2763 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2764 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2765 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2766 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2767 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2768 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2769 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2770 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2771 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2772 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2773 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2774 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2775 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2776 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2777 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2778 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2779 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2780 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2781 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2782 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2783 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2784 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2785 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2786 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2787 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2788 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2789 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2790 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2791 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2792 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2793 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2794 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2795 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2796 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2797 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2798 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2799 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2800 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2801 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2802 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2803 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2804 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2805 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2806 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2807 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2808 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2809 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2810 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2811 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2812 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2813 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2814 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2815 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2816 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2817 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2818 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2819 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2820 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2821 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2822 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2823 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2824 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2825 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2826 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2827 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2828 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2829 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2830 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2831 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2832 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2833 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2834 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2835 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2836 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2837 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2838 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2839 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2840 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2841 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2842 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2843 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2844 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2845 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2846 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2847 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2848 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2849 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2850 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2851 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2852 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2853 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2854 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2855 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2856 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2857 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2858 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2859 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2860 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2861 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2862 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2863 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2864 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2865 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2866 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2867 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2868 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2869 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2870 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2871 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2872 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2873 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2874 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2875 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2876 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2877 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2878 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2879 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2880 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2881 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2882 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2883 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2884 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2885 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2886 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2887 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2888 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2889 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2890 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2891 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2892 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2893 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2894 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2895 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2896 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2897 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2898 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2899 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2900 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2901 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2902 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2903 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2904 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2905 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2906 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2907 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2908 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2909 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2910 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2911 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2912 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2913 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2914 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2915 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2916 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2917 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2918 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2919 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2920 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2921 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2922 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2923 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2924 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2925 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2926 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2927 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2928 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2929 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2930 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2931 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2932 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2933 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2934 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2935 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2936 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2937 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2938 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2939 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2940 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2941 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2942 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2943 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2944 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2945 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2946 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2947 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2948 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2949 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2950 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2951 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2952 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2953 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2954 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2955 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2956 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2957 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2958 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2959 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2960 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2961 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2962 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2963 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2964 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2965 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2966 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2967 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2968 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2969 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2970 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2971 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2972 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2973 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2974 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2975 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2976 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2977 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2978 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2979 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2980 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2981 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2982 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2983 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2984 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2985 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2986 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2987 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2988 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2989 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2990 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2991 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2992 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2993 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2994 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2995 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_2996 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_2997 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_2998 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_2999 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3000 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3001 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3002 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3003 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3004 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3005 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3006 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3007 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3008 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3009 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3010 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3011 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3012 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3013 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3014 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3015 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3016 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3017 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3018 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3019 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3020 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3021 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3022 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3023 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3024 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3025 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3026 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3027 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3028 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3029 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3030 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3031 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3032 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3033 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3034 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3035 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3036 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3037 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3038 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3039 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3040 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3041 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3042 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3043 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3044 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3045 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3046 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3047 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3048 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3049 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3050 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3051 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3052 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3053 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3054 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3055 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3056 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3057 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3058 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3059 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3060 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3061 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3062 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3063 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3064 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3065 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3066 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3067 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3068 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3069 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3070 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3071 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3072 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3073 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3074 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3075 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3076 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3077 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3078 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3079 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3080 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3081 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3082 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3083 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3084 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3085 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3086 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3087 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3088 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3089 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3090 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3091 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3092 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3093 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3094 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3095 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3096 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3097 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3098 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3099 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3100 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3101 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3102 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3103 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3104 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3105 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3106 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3107 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3108 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3109 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3110 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3111 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3112 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3113 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3114 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3115 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3116 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3117 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3118 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3119 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3120 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3121 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3122 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3123 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3124 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3125 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3126 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3127 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3128 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3129 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3130 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3131 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3132 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3133 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3134 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3135 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3136 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3137 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3138 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3139 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3140 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3141 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3142 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3143 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3144 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3145 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3146 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3147 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3148 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3149 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3150 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3151 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3152 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3153 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3154 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3155 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3156 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3157 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3158 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3159 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3160 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3161 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3162 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3163 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3164 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3165 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3166 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3167 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3168 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3169 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3170 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3171 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3172 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3173 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3174 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3175 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3176 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3177 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3178 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3179 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3180 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3181 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3182 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3183 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3184 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3185 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3186 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3187 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3188 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3189 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3190 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3191 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3192 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3193 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3194 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3195 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3196 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3197 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3198 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3199 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3200 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3201 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3202 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3203 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3204 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3205 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3206 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3207 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3208 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3209 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3210 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3211 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3212 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3213 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3214 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3215 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3216 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3217 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3218 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3219 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3220 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3221 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3222 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3223 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3224 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3225 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3226 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3227 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3228 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3229 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3230 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3231 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3232 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3233 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3234 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3235 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3236 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3237 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3238 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3239 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3240 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3241 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3242 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3243 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3244 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3245 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3246 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3247 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3248 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3249 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3250 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3251 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3252 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3253 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3254 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3255 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3256 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3257 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3258 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3259 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3260 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3261 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3262 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3263 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3264 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3265 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3266 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3267 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3268 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3269 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3270 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3271 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3272 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3273 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3274 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3275 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3276 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3277 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3278 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3279 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3280 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3281 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3282 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3283 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3284 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3285 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3286 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3287 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3288 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3289 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3290 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3291 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3292 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3293 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3294 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3295 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3296 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3297 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3298 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3299 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3300 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3301 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3302 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3303 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3304 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3305 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3306 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3307 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3308 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3309 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3310 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3311 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3312 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3313 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3314 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3315 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3316 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3317 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3318 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3319 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3320 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3321 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3322 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3323 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3324 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3325 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3326 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3327 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3328 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3329 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3330 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3331 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3332 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3333 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3334 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3335 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3336 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3337 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3338 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3339 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3340 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3341 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3342 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3343 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3344 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3345 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3346 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3347 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3348 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3349 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3350 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3351 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3352 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3353 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3354 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3355 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3356 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3357 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3358 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3359 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3360 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3361 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3362 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3363 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3364 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3365 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3366 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3367 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3368 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3369 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3370 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3371 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3372 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3373 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3374 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3375 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3376 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3377 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3378 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3379 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3380 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3381 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3382 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3383 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3384 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3385 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3386 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3387 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3388 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3389 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3390 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3391 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3392 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3393 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3394 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3395 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3396 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3397 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3398 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3399 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3400 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3401 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3402 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3403 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3404 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3405 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3406 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3407 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3408 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3409 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3410 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3411 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3412 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3413 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3414 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3415 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3416 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3417 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3418 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3419 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3420 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3421 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3422 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3423 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3424 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3425 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3426 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3427 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3428 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3429 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3430 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3431 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3432 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3433 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3434 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3435 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3436 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3437 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3438 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3439 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3440 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3441 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3442 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3443 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3444 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3445 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3446 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3447 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3448 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3449 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3450 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3451 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3452 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3453 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3454 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3455 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3456 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3457 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3458 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3459 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3460 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3461 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3462 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3463 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3464 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3465 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3466 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3467 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3468 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3469 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3470 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3471 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3472 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3473 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3474 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3475 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3476 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3477 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3478 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3479 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3480 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3481 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3482 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3483 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3484 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3485 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3486 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3487 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3488 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3489 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3490 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3491 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3492 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3493 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3494 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3495 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3496 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3497 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3498 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3499 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3500 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3501 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3502 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3503 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3504 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3505 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3506 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3507 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3508 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3509 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3510 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3511 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3512 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3513 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3514 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3515 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3516 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3517 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3518 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3519 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3520 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3521 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3522 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3523 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3524 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3525 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3526 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3527 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3528 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3529 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3530 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3531 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3532 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3533 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3534 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3535 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3536 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3537 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3538 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3539 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3540 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3541 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3542 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3543 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3544 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3545 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3546 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3547 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3548 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3549 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3550 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3551 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3552 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3553 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3554 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3555 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3556 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3557 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3558 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3559 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3560 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3561 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3562 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3563 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3564 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3565 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3566 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3567 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3568 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3569 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3570 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3571 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3572 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3573 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3574 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3575 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3576 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3577 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3578 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3579 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3580 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3581 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3582 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3583 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3584 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3585 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3586 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3587 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3588 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3589 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3590 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3591 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3592 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3593 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3594 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3595 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3596 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3597 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3598 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3599 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3600 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3601 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3602 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3603 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3604 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3605 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3606 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3607 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3608 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3609 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3610 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3611 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3612 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3613 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3614 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3615 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3616 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3617 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3618 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3619 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3620 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3621 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3622 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3623 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3624 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3625 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3626 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3627 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3628 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3629 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3630 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3631 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3632 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3633 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3634 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3635 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3636 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3637 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3638 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3639 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3640 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3641 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3642 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3643 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3644 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3645 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3646 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3647 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3648 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3649 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3650 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3651 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3652 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3653 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3654 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3655 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3656 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3657 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3658 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3659 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3660 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3661 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3662 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3663 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3664 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3665 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3666 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3667 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3668 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3669 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3670 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3671 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3672 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3673 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3674 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3675 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3676 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3677 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3678 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3679 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3680 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3681 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3682 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3683 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3684 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3685 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3686 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3687 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3688 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3689 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3690 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3691 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3692 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3693 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3694 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3695 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3696 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3697 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3698 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3699 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3700 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3701 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3702 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3703 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3704 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3705 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3706 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3707 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3708 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3709 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3710 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3711 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3712 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3713 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3714 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3715 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3716 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3717 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3718 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3719 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3720 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3721 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3722 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3723 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3724 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3725 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3726 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3727 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3728 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3729 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3730 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3731 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3732 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3733 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3734 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3735 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3736 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3737 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3738 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3739 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3740 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3741 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3742 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3743 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3744 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3745 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3746 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3747 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3748 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3749 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3750 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3751 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3752 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3753 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3754 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3755 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3756 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3757 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3758 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3759 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3760 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3761 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3762 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3763 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3764 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3765 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3766 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3767 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3768 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3769 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3770 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3771 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3772 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3773 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3774 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3775 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3776 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3777 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3778 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3779 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3780 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3781 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3782 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3783 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3784 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3785 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3786 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3787 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3788 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3789 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3790 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3791 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3792 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3793 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3794 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3795 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3796 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3797 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3798 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3799 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3800 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3801 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3802 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3803 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3804 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3805 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3806 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3807 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3808 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3809 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3810 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3811 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3812 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3813 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3814 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3815 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3816 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3817 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3818 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3819 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3820 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3821 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3822 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3823 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3824 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3825 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3826 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3827 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3828 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3829 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3830 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3831 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3832 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3833 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3834 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3835 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3836 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3837 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3838 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3839 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3840 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3841 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3842 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3843 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3844 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3845 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3846 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3847 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3848 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3849 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3850 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3851 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3852 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3853 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3854 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3855 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3856 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3857 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3858 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3859 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3860 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3861 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3862 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3863 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3864 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3865 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3866 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3867 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3868 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3869 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3870 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3871 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3872 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3873 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3874 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3875 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3876 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3877 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3878 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3879 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3880 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3881 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3882 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3883 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3884 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3885 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3886 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3887 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3888 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3889 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3890 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3891 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3892 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3893 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3894 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3895 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3896 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3897 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3898 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3899 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3900 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3901 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3902 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3903 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3904 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3905 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3906 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3907 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3908 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3909 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3910 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3911 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3912 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3913 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3914 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3915 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3916 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3917 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3918 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3919 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3920 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3921 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3922 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3923 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3924 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3925 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3926 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3927 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3928 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3929 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3930 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3931 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3932 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3933 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3934 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3935 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3936 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3937 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3938 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3939 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3940 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3941 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3942 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3943 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3944 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3945 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3946 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3947 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3948 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3949 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3950 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3951 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3952 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3953 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3954 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3955 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3956 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3957 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3958 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3959 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3960 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3961 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3962 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3963 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3964 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3965 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3966 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3967 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3968 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3969 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3970 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3971 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3972 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3973 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3974 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3975 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3976 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3977 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3978 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3979 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3980 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3981 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3982 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3983 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3984 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3985 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3986 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3987 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3988 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3989 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_3990 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3991 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_3992 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_3993 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3994 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3995 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3996 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3997 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3998 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_3999 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4000 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4001 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4002 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4003 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4004 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4005 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4006 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4007 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4008 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4009 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4010 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4011 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4012 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4013 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4014 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4015 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4016 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4017 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4018 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4019 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4020 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4021 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4022 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4023 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4024 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4025 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4026 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4027 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4028 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4029 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4030 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4031 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4032 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4033 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4034 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4035 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4036 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4037 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4038 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4039 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4040 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4041 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4042 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4043 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4044 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4045 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4046 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4047 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4048 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4049 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4050 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4051 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4052 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4053 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4054 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4055 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4056 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4057 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4058 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4059 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4060 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4061 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4062 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4063 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4064 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4065 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4066 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4067 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4068 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4069 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4070 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4071 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4072 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4073 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4074 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4075 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4076 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4077 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4078 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4079 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4080 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4081 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4082 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4083 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4084 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4085 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4086 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4087 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4088 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4089 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4090 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4091 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4092 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4093 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4094 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4095 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4096 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4097 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4098 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4099 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4100 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4101 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4102 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4103 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4104 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4105 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4106 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4107 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4108 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4109 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4110 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4111 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4112 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4113 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4114 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4115 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4116 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4117 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4118 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4119 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4120 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4121 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4122 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4123 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4124 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4125 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4126 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4127 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4128 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4129 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4130 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4131 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4132 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4133 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4134 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4135 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4136 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4137 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4138 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4139 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4140 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4141 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4142 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4143 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4144 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4145 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4146 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4147 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4148 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4149 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4150 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4151 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4152 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4153 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4154 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4155 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4156 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4157 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4158 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4159 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4160 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4161 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4162 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4163 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4164 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4165 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4166 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4167 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4168 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4169 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4170 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4171 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4172 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4173 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4174 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4175 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4176 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4177 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4178 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4179 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4180 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4181 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4182 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4183 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4184 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4185 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4186 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4187 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4188 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4189 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4190 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4191 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4192 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4193 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4194 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4195 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4196 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4197 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4198 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4199 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4200 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4201 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4202 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4203 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4204 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4205 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4206 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4207 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4208 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4209 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4210 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4211 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4212 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4213 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4214 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4215 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4216 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4217 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4218 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4219 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4220 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4221 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4222 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4223 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4224 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4225 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4226 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4227 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4228 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4229 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4230 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4231 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4232 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4233 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4234 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4235 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4236 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4237 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4238 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4239 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4240 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4241 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4242 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4243 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4244 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4245 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4246 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4247 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4248 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4249 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4250 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4251 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4252 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4253 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4254 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4255 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4256 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4257 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4258 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4259 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4260 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4261 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4262 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4263 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4264 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4265 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4266 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4267 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4268 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4269 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4270 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4271 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4272 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4273 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4274 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4275 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4276 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4277 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4278 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4279 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4280 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4281 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4282 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4283 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4284 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4285 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4286 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4287 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4288 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4289 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4290 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4291 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4292 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4293 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4294 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4295 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4296 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4297 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4298 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4299 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4300 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4301 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4302 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4303 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4304 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4305 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4306 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4307 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4308 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4309 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4310 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4311 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4312 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4313 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4314 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4315 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4316 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4317 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4318 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4319 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4320 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4321 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4322 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4323 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4324 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4325 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4326 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4327 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4328 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4329 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4330 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4331 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4332 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4333 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4334 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4335 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4336 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4337 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4338 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4339 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4340 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4341 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4342 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4343 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4344 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4345 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4346 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4347 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4348 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4349 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4350 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4351 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4352 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4353 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4354 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4355 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4356 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4357 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4358 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4359 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4360 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4361 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4362 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4363 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4364 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4365 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4366 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4367 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4368 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4369 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4370 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4371 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4372 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4373 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4374 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4375 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4376 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4377 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4378 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4379 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4380 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4381 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4382 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4383 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4384 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4385 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4386 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4387 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4388 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4389 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4390 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4391 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4392 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4393 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4394 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4395 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4396 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4397 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4398 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4399 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4400 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4401 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4402 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4403 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4404 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4405 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4406 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4407 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4408 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4409 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4410 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4411 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4412 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4413 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4414 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4415 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4416 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4417 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4418 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4419 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4420 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4421 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4422 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4423 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4424 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4425 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4426 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4427 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4428 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4429 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4430 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4431 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4432 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4433 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4434 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4435 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4436 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4437 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4438 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4439 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4440 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4441 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4442 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4443 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4444 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4445 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4446 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4447 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4448 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4449 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4450 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4451 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4452 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4453 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4454 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4455 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4456 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4457 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4458 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4459 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4460 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4461 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4462 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4463 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4464 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4465 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4466 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4467 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4468 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4469 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4470 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4471 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4472 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4473 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4474 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4475 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4476 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4477 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4478 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4479 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4480 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4481 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4482 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4483 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4484 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4485 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4486 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4487 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4488 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4489 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4490 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4491 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4492 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4493 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4494 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4495 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4496 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4497 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4498 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4499 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4500 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4501 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4502 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4503 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4504 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4505 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4506 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4507 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4508 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4509 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4510 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4511 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4512 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4513 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4514 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4515 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4516 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4517 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4518 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4519 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4520 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4521 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4522 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4523 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4524 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4525 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4526 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4527 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4528 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4529 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4530 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4531 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4532 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4533 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4534 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4535 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4536 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4537 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4538 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4539 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4540 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4541 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4542 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4543 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4544 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4545 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4546 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4547 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4548 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4549 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4550 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4551 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4552 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4553 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4554 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4555 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4556 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4557 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4558 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4559 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4560 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4561 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4562 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4563 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4564 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4565 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4566 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4567 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4568 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4569 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4570 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4571 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4572 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4573 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4574 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4575 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4576 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4577 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4578 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4579 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4580 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4581 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4582 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4583 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4584 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4585 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4586 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4587 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4588 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4589 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4590 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4591 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4592 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4593 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4594 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4595 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4596 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4597 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4598 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4599 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4600 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4601 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4602 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4603 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4604 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4605 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4606 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4607 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4608 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4609 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4610 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4611 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4612 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4613 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4614 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4615 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4616 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4617 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4618 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4619 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4620 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4621 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4622 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4623 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4624 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4625 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4626 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4627 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4628 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4629 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4630 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4631 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4632 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4633 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4634 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4635 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4636 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4637 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4638 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4639 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4640 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4641 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4642 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4643 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4644 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4645 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4646 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4647 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4648 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4649 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4650 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4651 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4652 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4653 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4654 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4655 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4656 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4657 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4658 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4659 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4660 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4661 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4662 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4663 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4664 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4665 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4666 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4667 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4668 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4669 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4670 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4671 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4672 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4673 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4674 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4675 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4676 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4677 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4678 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4679 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4680 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4681 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4682 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4683 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4684 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4685 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4686 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4687 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4688 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4689 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4690 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4691 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4692 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4693 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4694 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4695 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4696 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4697 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4698 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4699 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4700 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4701 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4702 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4703 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4704 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4705 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4706 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4707 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4708 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4709 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4710 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4711 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4712 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4713 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4714 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4715 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4716 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4717 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4718 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4719 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4720 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4721 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4722 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4723 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4724 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4725 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4726 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4727 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4728 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4729 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4730 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4731 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4732 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4733 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4734 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4735 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4736 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4737 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4738 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4739 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4740 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4741 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4742 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4743 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4744 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4745 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4746 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4747 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4748 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4749 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4750 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4751 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4752 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4753 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4754 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4755 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4756 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4757 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4758 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4759 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4760 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4761 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4762 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4763 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4764 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4765 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4766 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4767 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4768 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4769 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4770 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4771 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4772 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4773 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4774 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4775 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4776 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4777 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4778 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4779 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4780 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4781 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4782 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4783 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4784 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4785 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4786 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4787 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4788 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4789 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4790 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4791 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4792 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4793 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4794 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4795 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4796 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4797 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4798 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4799 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4800 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4801 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4802 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4803 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4804 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4805 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4806 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4807 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4808 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4809 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4810 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4811 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4812 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4813 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4814 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4815 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4816 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4817 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4818 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4819 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4820 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4821 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4822 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4823 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4824 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4825 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4826 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4827 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4828 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4829 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4830 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4831 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4832 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4833 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4834 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4835 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4836 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4837 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4838 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4839 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4840 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4841 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4842 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4843 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4844 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4845 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4846 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4847 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4848 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4849 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4850 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4851 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4852 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4853 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4854 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4855 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4856 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4857 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4858 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4859 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4860 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4861 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4862 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4863 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4864 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4865 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4866 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4867 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4868 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4869 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4870 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4871 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4872 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4873 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4874 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4875 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4876 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4877 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4878 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4879 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4880 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4881 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4882 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4883 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4884 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4885 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4886 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4887 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4888 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4889 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4890 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4891 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4892 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4893 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4894 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4895 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4896 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4897 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4898 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4899 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4900 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4901 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4902 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4903 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4904 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4905 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4906 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4907 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4908 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4909 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4910 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4911 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4912 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4913 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4914 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4915 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4916 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4917 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4918 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4919 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4920 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4921 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4922 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4923 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4924 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4925 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4926 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4927 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4928 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4929 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4930 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4931 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4932 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4933 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4934 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4935 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4936 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4937 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4938 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4939 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4940 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4941 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4942 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4943 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4944 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4945 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4946 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4947 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4948 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4949 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4950 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4951 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4952 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4953 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4954 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4955 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4956 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4957 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4958 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4959 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4960 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4961 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4962 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4963 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4964 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4965 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4966 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4967 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4968 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4969 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4970 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4971 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4972 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4973 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4974 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4975 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4976 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4977 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4978 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4979 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4980 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4981 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4982 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4983 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4984 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4985 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4986 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4987 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4988 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4989 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4990 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4991 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4992 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4993 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4994 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_4995 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4996 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_4997 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_4998 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_4999 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5000 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5001 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5002 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5003 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5004 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5005 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5006 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5007 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5008 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5009 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5010 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5011 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5012 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5013 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5014 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5015 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5016 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5017 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5018 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5019 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5020 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5021 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5022 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5023 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5024 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5025 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5026 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5027 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5028 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5029 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5030 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5031 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5032 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5033 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5034 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5035 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5036 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5037 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5038 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5039 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5040 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5041 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5042 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5043 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5044 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5045 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5046 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5047 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5048 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5049 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5050 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5051 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5052 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5053 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5054 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5055 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5056 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5057 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5058 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5059 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5060 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5061 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5062 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5063 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5064 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5065 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5066 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5067 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5068 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5069 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5070 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5071 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5072 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5073 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5074 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5075 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5076 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5077 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5078 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5079 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5080 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5081 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5082 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5083 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5084 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5085 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5086 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5087 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5088 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5089 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5090 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5091 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5092 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5093 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5094 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5095 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5096 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5097 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5098 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5099 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5100 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5101 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5102 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5103 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5104 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5105 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5106 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5107 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5108 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5109 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5110 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5111 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5112 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5113 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5114 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5115 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5116 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5117 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5118 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5119 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5120 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5121 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5122 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5123 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5124 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5125 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5126 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5127 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5128 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5129 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5130 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5131 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5132 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5133 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5134 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5135 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5136 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5137 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5138 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5139 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5140 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5141 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5142 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5143 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5144 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5145 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5146 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5147 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5148 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5149 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5150 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5151 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5152 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5153 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5154 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5155 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5156 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5157 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5158 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5159 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5160 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5161 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5162 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5163 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5164 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5165 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5166 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5167 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5168 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5169 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5170 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5171 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5172 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5173 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5174 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5175 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5176 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5177 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5178 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5179 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5180 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5181 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5182 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5183 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5184 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5185 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5186 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5187 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5188 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5189 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5190 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5191 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5192 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5193 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5194 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5195 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5196 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5197 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5198 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5199 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5200 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5201 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5202 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5203 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5204 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5205 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5206 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5207 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5208 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5209 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5210 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5211 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5212 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5213 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5214 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5215 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5216 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5217 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5218 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5219 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5220 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5221 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5222 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5223 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5224 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5225 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5226 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5227 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5228 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5229 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5230 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5231 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5232 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5233 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5234 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5235 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5236 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5237 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5238 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5239 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5240 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5241 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5242 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5243 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5244 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5245 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5246 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5247 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5248 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5249 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5250 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5251 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5252 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5253 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5254 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5255 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5256 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5257 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5258 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5259 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5260 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5261 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5262 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5263 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5264 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5265 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5266 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5267 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5268 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5269 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5270 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5271 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5272 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5273 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5274 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5275 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5276 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5277 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5278 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5279 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5280 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5281 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5282 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5283 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5284 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5285 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5286 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5287 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5288 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5289 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5290 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5291 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5292 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5293 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5294 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5295 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5296 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5297 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5298 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5299 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5300 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5301 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5302 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5303 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5304 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5305 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5306 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5307 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5308 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5309 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5310 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5311 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5312 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5313 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5314 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5315 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5316 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5317 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5318 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5319 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5320 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5321 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5322 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5323 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5324 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5325 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5326 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5327 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5328 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5329 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5330 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5331 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5332 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5333 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5334 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5335 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5336 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5337 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5338 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5339 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5340 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5341 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5342 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5343 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5344 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5345 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5346 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5347 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5348 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5349 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5350 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5351 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5352 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5353 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5354 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5355 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5356 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5357 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5358 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5359 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5360 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5361 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5362 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5363 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5364 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5365 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5366 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5367 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5368 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5369 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5370 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5371 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5372 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5373 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5374 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5375 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5376 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5377 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5378 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5379 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5380 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5381 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5382 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5383 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5384 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5385 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5386 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5387 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5388 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5389 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5390 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5391 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5392 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5393 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5394 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5395 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5396 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5397 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5398 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5399 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5400 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5401 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5402 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5403 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5404 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5405 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5406 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5407 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5408 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5409 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5410 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5411 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5412 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5413 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5414 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5415 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5416 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5417 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5418 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5419 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5420 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5421 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5422 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5423 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5424 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5425 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5426 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5427 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5428 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5429 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5430 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5431 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5432 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5433 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5434 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5435 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5436 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5437 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5438 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5439 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5440 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5441 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5442 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5443 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5444 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5445 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5446 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5447 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5448 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5449 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5450 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5451 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5452 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5453 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5454 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5455 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5456 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5457 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5458 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5459 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5460 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5461 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5462 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5463 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5464 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5465 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5466 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5467 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5468 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5469 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5470 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5471 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5472 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5473 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5474 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5475 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5476 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5477 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5478 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5479 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5480 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5481 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5482 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5483 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5484 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5485 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5486 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5487 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5488 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5489 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5490 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5491 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5492 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5493 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5494 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5495 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5496 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5497 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5498 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5499 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5500 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5501 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5502 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5503 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5504 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5505 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5506 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5507 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5508 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5509 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5510 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5511 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5512 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5513 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5514 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5515 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5516 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5517 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5518 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5519 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5520 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5521 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5522 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5523 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5524 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5525 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5526 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5527 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5528 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5529 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5530 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5531 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5532 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5533 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5534 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5535 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5536 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5537 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5538 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5539 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5540 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5541 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5542 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5543 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5544 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5545 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5546 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5547 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5548 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5549 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5550 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5551 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5552 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5553 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5554 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5555 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5556 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5557 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5558 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5559 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5560 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5561 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5562 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5563 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5564 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5565 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5566 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5567 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5568 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5569 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5570 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5571 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5572 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5573 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5574 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5575 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5576 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5577 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5578 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5579 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5580 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5581 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5582 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5583 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5584 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5585 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5586 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5587 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5588 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5589 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5590 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5591 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5592 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5593 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5594 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5595 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5596 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5597 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5598 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5599 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5600 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5601 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5602 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5603 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5604 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5605 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5606 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5607 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5608 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5609 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5610 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5611 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5612 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5613 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5614 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5615 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5616 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5617 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5618 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5619 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5620 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5621 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5622 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5623 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5624 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5625 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5626 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5627 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5628 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5629 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5630 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5631 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5632 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5633 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5634 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5635 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5636 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5637 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5638 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5639 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5640 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5641 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5642 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5643 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5644 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5645 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5646 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5647 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5648 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5649 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5650 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5651 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5652 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5653 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5654 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5655 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5656 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5657 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5658 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5659 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5660 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5661 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5662 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5663 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5664 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5665 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5666 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5667 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5668 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5669 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5670 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5671 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5672 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5673 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5674 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5675 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5676 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5677 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5678 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5679 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5680 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5681 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5682 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5683 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5684 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5685 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5686 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5687 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5688 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5689 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5690 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5691 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5692 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5693 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5694 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5695 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5696 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5697 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5698 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5699 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5700 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5701 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5702 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5703 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5704 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5705 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5706 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5707 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5708 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5709 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5710 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5711 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5712 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5713 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5714 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5715 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5716 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5717 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5718 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5719 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5720 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5721 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5722 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5723 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5724 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5725 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5726 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5727 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5728 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5729 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5730 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5731 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5732 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5733 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5734 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5735 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5736 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5737 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5738 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5739 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5740 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5741 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5742 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5743 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5744 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5745 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5746 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5747 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5748 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5749 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5750 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5751 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5752 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5753 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5754 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5755 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5756 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5757 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5758 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5759 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5760 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5761 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5762 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5763 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5764 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5765 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5766 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5767 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5768 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5769 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5770 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5771 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5772 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5773 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5774 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5775 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5776 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5777 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5778 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5779 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5780 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5781 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5782 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5783 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5784 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5785 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5786 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5787 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5788 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5789 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5790 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5791 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5792 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5793 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5794 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5795 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5796 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5797 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5798 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5799 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5800 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5801 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5802 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5803 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5804 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5805 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5806 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5807 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5808 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5809 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5810 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5811 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5812 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5813 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5814 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5815 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5816 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5817 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5818 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5819 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5820 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5821 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5822 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5823 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5824 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5825 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5826 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5827 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5828 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5829 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5830 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5831 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5832 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5833 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5834 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5835 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5836 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5837 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5838 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5839 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5840 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5841 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5842 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5843 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5844 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5845 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5846 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5847 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5848 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5849 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5850 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5851 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5852 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5853 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5854 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5855 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5856 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5857 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5858 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5859 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5860 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5861 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5862 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5863 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5864 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5865 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5866 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5867 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5868 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5869 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5870 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5871 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5872 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5873 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5874 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5875 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5876 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5877 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5878 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5879 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5880 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5881 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5882 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5883 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5884 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5885 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5886 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5887 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5888 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5889 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5890 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5891 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5892 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5893 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5894 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5895 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5896 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5897 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5898 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5899 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5900 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5901 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5902 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5903 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5904 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5905 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5906 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5907 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5908 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5909 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5910 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5911 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5912 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5913 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5914 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5915 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5916 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5917 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5918 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5919 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5920 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5921 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5922 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5923 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5924 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5925 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5926 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5927 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5928 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5929 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5930 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5931 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5932 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5933 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5934 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5935 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5936 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5937 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5938 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5939 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5940 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5941 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5942 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5943 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5944 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5945 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5946 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5947 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5948 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5949 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5950 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5951 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5952 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5953 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5954 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5955 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5956 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5957 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5958 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5959 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5960 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5961 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5962 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5963 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5964 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5965 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5966 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5967 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5968 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5969 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5970 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5971 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5972 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5973 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5974 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5975 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5976 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5977 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5978 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5979 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5980 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5981 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5982 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5983 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5984 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5985 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5986 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_5987 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5988 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5989 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5990 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_5991 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5992 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5993 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5994 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5995 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5996 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5997 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_5998 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_5999 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6000 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6001 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6002 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6003 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6004 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6005 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6006 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6007 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6008 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6009 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6010 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6011 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6012 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6013 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6014 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6015 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6016 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6017 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6018 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6019 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6020 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6021 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6022 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6023 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6024 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6025 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6026 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6027 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6028 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6029 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6030 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6031 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6032 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6033 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6034 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6035 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6036 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6037 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6038 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6039 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6040 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6041 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6042 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6043 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6044 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6045 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6046 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6047 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6048 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6049 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6050 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6051 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6052 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6053 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6054 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6055 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6056 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6057 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6058 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6059 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6060 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6061 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6062 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6063 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6064 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6065 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6066 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6067 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6068 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6069 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6070 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6071 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6072 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6073 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6074 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6075 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6076 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6077 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6078 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6079 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6080 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6081 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6082 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6083 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6084 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6085 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6086 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6087 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6088 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6089 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6090 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6091 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6092 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6093 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6094 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6095 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6096 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6097 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6098 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6099 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6100 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6101 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6102 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6103 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6104 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6105 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6106 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6107 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6108 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6109 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6110 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6111 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6112 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6113 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6114 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6115 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6116 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6117 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6118 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6119 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6120 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6121 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6122 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6123 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6124 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6125 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6126 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6127 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6128 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6129 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6130 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6131 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6132 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6133 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6134 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6135 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6136 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6137 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6138 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6139 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6140 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6141 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6142 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6143 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6144 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6145 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6146 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6147 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6148 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6149 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6150 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6151 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6152 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6153 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6154 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6155 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6156 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6157 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6158 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6159 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6160 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6161 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6162 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6163 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6164 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6165 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6166 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6167 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6168 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6169 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6170 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6171 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6172 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6173 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6174 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6175 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6176 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6177 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6178 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6179 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6180 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6181 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6182 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6183 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6184 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6185 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6186 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6187 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6188 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6189 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6190 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6191 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6192 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6193 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6194 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6195 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6196 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6197 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6198 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6199 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6200 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6201 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6202 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6203 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6204 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6205 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6206 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6207 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6208 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6209 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6210 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6211 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6212 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6213 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6214 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6215 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6216 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6217 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6218 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6219 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6220 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6221 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6222 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6223 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6224 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6225 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6226 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6227 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6228 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6229 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6230 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6231 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6232 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6233 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6234 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6235 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6236 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6237 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6238 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6239 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6240 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6241 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6242 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6243 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6244 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6245 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6246 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6247 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6248 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6249 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6250 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6251 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6252 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6253 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6254 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6255 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6256 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6257 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6258 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6259 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6260 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6261 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6262 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6263 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6264 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6265 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6266 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6267 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6268 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6269 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6270 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6271 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6272 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6273 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6274 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6275 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6276 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6277 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6278 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6279 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6280 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6281 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6282 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6283 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6284 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6285 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6286 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6287 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6288 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6289 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6290 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6291 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6292 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6293 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6294 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6295 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6296 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6297 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6298 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6299 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6300 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6301 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6302 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6303 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6304 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6305 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6306 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6307 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6308 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6309 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6310 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6311 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6312 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6313 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6314 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6315 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6316 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6317 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6318 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6319 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6320 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6321 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6322 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6323 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6324 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6325 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6326 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6327 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6328 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6329 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6330 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6331 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6332 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6333 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6334 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6335 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6336 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6337 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6338 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6339 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6340 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6341 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6342 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6343 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6344 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6345 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6346 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6347 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6348 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6349 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6350 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6351 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6352 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6353 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6354 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6355 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6356 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6357 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6358 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6359 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6360 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6361 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6362 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6363 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6364 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6365 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6366 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6367 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6368 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6369 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6370 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6371 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6372 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6373 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6374 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6375 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6376 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6377 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6378 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6379 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6380 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6381 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6382 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6383 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6384 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6385 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6386 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6387 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6388 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6389 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6390 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6391 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6392 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6393 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6394 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6395 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6396 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6397 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6398 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6399 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6400 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6401 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6402 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6403 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6404 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6405 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6406 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6407 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6408 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6409 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6410 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6411 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6412 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6413 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6414 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6415 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6416 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6417 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6418 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6419 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6420 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6421 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6422 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6423 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6424 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6425 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6426 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6427 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6428 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6429 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6430 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6431 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6432 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6433 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6434 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6435 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6436 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6437 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6438 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6439 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6440 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6441 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6442 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6443 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6444 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6445 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6446 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6447 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6448 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6449 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6450 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6451 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6452 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6453 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6454 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6455 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6456 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6457 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6458 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6459 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6460 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6461 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6462 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6463 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6464 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6465 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6466 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6467 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6468 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6469 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6470 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6471 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6472 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6473 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6474 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6475 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6476 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6477 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6478 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6479 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6480 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6481 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6482 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6483 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6484 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6485 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6486 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6487 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6488 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6489 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6490 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6491 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6492 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6493 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6494 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6495 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6496 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6497 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6498 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6499 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6500 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6501 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6502 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6503 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6504 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6505 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6506 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6507 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6508 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6509 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6510 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6511 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6512 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6513 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6514 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6515 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6516 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6517 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6518 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6519 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6520 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6521 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6522 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6523 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6524 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6525 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6526 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6527 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6528 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6529 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6530 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6531 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6532 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6533 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6534 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6535 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6536 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6537 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6538 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6539 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6540 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6541 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6542 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6543 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6544 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6545 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6546 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6547 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6548 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6549 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6550 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6551 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6552 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6553 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6554 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6555 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6556 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6557 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6558 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6559 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6560 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6561 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6562 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6563 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6564 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6565 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6566 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6567 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6568 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6569 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6570 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6571 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6572 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6573 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6574 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6575 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6576 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6577 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6578 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6579 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6580 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6581 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6582 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6583 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6584 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6585 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6586 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6587 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6588 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6589 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6590 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6591 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6592 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6593 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6594 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6595 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6596 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6597 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6598 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6599 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6600 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6601 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6602 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6603 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6604 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6605 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6606 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6607 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6608 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6609 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6610 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6611 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6612 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6613 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6614 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6615 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6616 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6617 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6618 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6619 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6620 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6621 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6622 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6623 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6624 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6625 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6626 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6627 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6628 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6629 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6630 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6631 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6632 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6633 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6634 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6635 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6636 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6637 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6638 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6639 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6640 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6641 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6642 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6643 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6644 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6645 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6646 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6647 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6648 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6649 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6650 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6651 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6652 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6653 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6654 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6655 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6656 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6657 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6658 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6659 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6660 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6661 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6662 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6663 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6664 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6665 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6666 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6667 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6668 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6669 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6670 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6671 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6672 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6673 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6674 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6675 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6676 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6677 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6678 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6679 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6680 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6681 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6682 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6683 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6684 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6685 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6686 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6687 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6688 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6689 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6690 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6691 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6692 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6693 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6694 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6695 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6696 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6697 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6698 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6699 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6700 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6701 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6702 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6703 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6704 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6705 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6706 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6707 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6708 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6709 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6710 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6711 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6712 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6713 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6714 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6715 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6716 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6717 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6718 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6719 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6720 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6721 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6722 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6723 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6724 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6725 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6726 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6727 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6728 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6729 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6730 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6731 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6732 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6733 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6734 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6735 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6736 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6737 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6738 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6739 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6740 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6741 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6742 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6743 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6744 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6745 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6746 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6747 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6748 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6749 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6750 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6751 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6752 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6753 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6754 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6755 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6756 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6757 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6758 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6759 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6760 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6761 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6762 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6763 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6764 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6765 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6766 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6767 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6768 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6769 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6770 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6771 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6772 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6773 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6774 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6775 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6776 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6777 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6778 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6779 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6780 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6781 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6782 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6783 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6784 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6785 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6786 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6787 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6788 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6789 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6790 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6791 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6792 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6793 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6794 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6795 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6796 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6797 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6798 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6799 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6800 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6801 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6802 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6803 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6804 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6805 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6806 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6807 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6808 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6809 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6810 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6811 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6812 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6813 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6814 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6815 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6816 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6817 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6818 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6819 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6820 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6821 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6822 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6823 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6824 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6825 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6826 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6827 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6828 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6829 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6830 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6831 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6832 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6833 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6834 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6835 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6836 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6837 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6838 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6839 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6840 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6841 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6842 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6843 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6844 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6845 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6846 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6847 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6848 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6849 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6850 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6851 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6852 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6853 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6854 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6855 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6856 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6857 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6858 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6859 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6860 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6861 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6862 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6863 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6864 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6865 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6866 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6867 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6868 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6869 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6870 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6871 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6872 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6873 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6874 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6875 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6876 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6877 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6878 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6879 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6880 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6881 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6882 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6883 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6884 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6885 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6886 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6887 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6888 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6889 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6890 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6891 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6892 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6893 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6894 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6895 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6896 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6897 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6898 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6899 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6900 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6901 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6902 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6903 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6904 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6905 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6906 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6907 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6908 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6909 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6910 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6911 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6912 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6913 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6914 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6915 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6916 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6917 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6918 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6919 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6920 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6921 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6922 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6923 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6924 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6925 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6926 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6927 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6928 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6929 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6930 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6931 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6932 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6933 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6934 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6935 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6936 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6937 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6938 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6939 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6940 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6941 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6942 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6943 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6944 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6945 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6946 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6947 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6948 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6949 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6950 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6951 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6952 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6953 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6954 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6955 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6956 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6957 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6958 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6959 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6960 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6961 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6962 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6963 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6964 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6965 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6966 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6967 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6968 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6969 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6970 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6971 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6972 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6973 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6974 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6975 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6976 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6977 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6978 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6979 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6980 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_6981 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_6982 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6983 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6984 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6985 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6986 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6987 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6988 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6989 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6990 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6991 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6992 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6993 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6994 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6995 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6996 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6997 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_6998 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_6999 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7000 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7001 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7002 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7003 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7004 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7005 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7006 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7007 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7008 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7009 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7010 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7011 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7012 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7013 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7014 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7015 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_7016 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_7017 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_7018 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7019 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7020 (  );
sky130_fd_sc_hs__fill_1 sky130_fd_sc_hs__fill_1_7021 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_7022 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7023 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7024 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7025 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7026 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7027 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7028 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7029 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7030 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7031 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7032 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7033 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7034 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7035 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7036 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7037 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7038 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7039 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7040 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7041 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7042 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7043 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7044 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7045 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7046 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7047 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7048 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7049 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7050 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7051 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7052 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7053 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7054 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7055 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7056 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7057 (  );
sky130_fd_sc_hs__fill_4 sky130_fd_sc_hs__fill_4_7058 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7059 (  );
sky130_fd_sc_hs__fill_8 sky130_fd_sc_hs__fill_8_7060 (  );
sky130_fd_sc_hs__fill_2 sky130_fd_sc_hs__fill_2_7061 (  );

endmodule
