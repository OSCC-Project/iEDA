//Generate the verilog at 2023-03-24T11:22:18
module gcd (
clk,
req_msg[0],
req_msg[1],
req_msg[2],
req_msg[3],
req_msg[4],
req_msg[5],
req_msg[6],
req_msg[7],
req_msg[8],
req_msg[9],
req_msg[10],
req_msg[11],
req_msg[12],
req_msg[13],
req_msg[14],
req_msg[15],
req_msg[16],
req_msg[17],
req_msg[18],
req_msg[19],
req_msg[20],
req_msg[21],
req_msg[22],
req_msg[23],
req_msg[24],
req_msg[25],
req_msg[26],
req_msg[27],
req_msg[28],
req_msg[29],
req_msg[30],
req_msg[31],
req_rdy,
req_val,
reset,
resp_msg[0],
resp_msg[1],
resp_msg[2],
resp_msg[3],
resp_msg[4],
resp_msg[5],
resp_msg[6],
resp_msg[7],
resp_msg[8],
resp_msg[9],
resp_msg[10],
resp_msg[11],
resp_msg[12],
resp_msg[13],
resp_msg[14],
resp_msg[15],
resp_rdy,
resp_val
);

input clk ;
input req_msg[0] ;
input req_msg[1] ;
input req_msg[2] ;
input req_msg[3] ;
input req_msg[4] ;
input req_msg[5] ;
input req_msg[6] ;
input req_msg[7] ;
input req_msg[8] ;
input req_msg[9] ;
input req_msg[10] ;
input req_msg[11] ;
input req_msg[12] ;
input req_msg[13] ;
input req_msg[14] ;
input req_msg[15] ;
input req_msg[16] ;
input req_msg[17] ;
input req_msg[18] ;
input req_msg[19] ;
input req_msg[20] ;
input req_msg[21] ;
input req_msg[22] ;
input req_msg[23] ;
input req_msg[24] ;
input req_msg[25] ;
input req_msg[26] ;
input req_msg[27] ;
input req_msg[28] ;
input req_msg[29] ;
input req_msg[30] ;
input req_msg[31] ;
output req_rdy ;
input req_val ;
input reset ;
output resp_msg[0] ;
output resp_msg[1] ;
output resp_msg[2] ;
output resp_msg[3] ;
output resp_msg[4] ;
output resp_msg[5] ;
output resp_msg[6] ;
output resp_msg[7] ;
output resp_msg[8] ;
output resp_msg[9] ;
output resp_msg[10] ;
output resp_msg[11] ;
output resp_msg[12] ;
output resp_msg[13] ;
output resp_msg[14] ;
output resp_msg[15] ;
input resp_rdy ;
output resp_val ;

wire \ctrl$a_mux_sel[0] ;
wire \ctrl$a_mux_sel[1] ;
wire ctrl$a_reg_en ;
wire ctrl$b_mux_sel ;
wire ctrl$b_reg_en ;
wire ctrl$is_a_lt_b ;
wire ctrl$is_b_zero ;
wire \ctrl/_00_ ;
wire \ctrl/_01_ ;
wire \ctrl/_02_ ;
wire \ctrl/_03_ ;
wire \ctrl/_04_ ;
wire \ctrl/_05_ ;
wire \ctrl/_06_ ;
wire \ctrl/_07_ ;
wire \ctrl/_08_ ;
wire \ctrl/_09_ ;
wire \ctrl/_10_ ;
wire \ctrl/_11_ ;
wire \ctrl/_12_ ;
wire \ctrl/_13_ ;
wire \ctrl/_14_ ;
wire \ctrl/_15_ ;
wire \ctrl/_16_ ;
wire \ctrl/curr_state__0[0] ;
wire \ctrl/curr_state__0[1] ;
wire \ctrl/next_state__0[0] ;
wire \ctrl/next_state__0[1] ;
wire \ctrl/state/_00_ ;
wire \ctrl/state/_01_ ;
wire \ctrl/state/_02_ ;
wire \ctrl/state/_03_ ;
wire \ctrl/state/_04_ ;
wire \ctrl/state/_05_ ;
wire \ctrl/state/_06_ ;
wire \dpath/a_lt_b$in0[0] ;
wire \dpath/a_lt_b$in0[10] ;
wire \dpath/a_lt_b$in0[11] ;
wire \dpath/a_lt_b$in0[12] ;
wire \dpath/a_lt_b$in0[13] ;
wire \dpath/a_lt_b$in0[14] ;
wire \dpath/a_lt_b$in0[15] ;
wire \dpath/a_lt_b$in0[1] ;
wire \dpath/a_lt_b$in0[2] ;
wire \dpath/a_lt_b$in0[3] ;
wire \dpath/a_lt_b$in0[4] ;
wire \dpath/a_lt_b$in0[5] ;
wire \dpath/a_lt_b$in0[6] ;
wire \dpath/a_lt_b$in0[7] ;
wire \dpath/a_lt_b$in0[8] ;
wire \dpath/a_lt_b$in0[9] ;
wire \dpath/a_lt_b$in1[0] ;
wire \dpath/a_lt_b$in1[10] ;
wire \dpath/a_lt_b$in1[11] ;
wire \dpath/a_lt_b$in1[12] ;
wire \dpath/a_lt_b$in1[13] ;
wire \dpath/a_lt_b$in1[14] ;
wire \dpath/a_lt_b$in1[15] ;
wire \dpath/a_lt_b$in1[1] ;
wire \dpath/a_lt_b$in1[2] ;
wire \dpath/a_lt_b$in1[3] ;
wire \dpath/a_lt_b$in1[4] ;
wire \dpath/a_lt_b$in1[5] ;
wire \dpath/a_lt_b$in1[6] ;
wire \dpath/a_lt_b$in1[7] ;
wire \dpath/a_lt_b$in1[8] ;
wire \dpath/a_lt_b$in1[9] ;
wire \dpath/a_mux$out[0] ;
wire \dpath/a_mux$out[10] ;
wire \dpath/a_mux$out[11] ;
wire \dpath/a_mux$out[12] ;
wire \dpath/a_mux$out[13] ;
wire \dpath/a_mux$out[14] ;
wire \dpath/a_mux$out[15] ;
wire \dpath/a_mux$out[1] ;
wire \dpath/a_mux$out[2] ;
wire \dpath/a_mux$out[3] ;
wire \dpath/a_mux$out[4] ;
wire \dpath/a_mux$out[5] ;
wire \dpath/a_mux$out[6] ;
wire \dpath/a_mux$out[7] ;
wire \dpath/a_mux$out[8] ;
wire \dpath/a_mux$out[9] ;
wire \dpath/b_mux$out[0] ;
wire \dpath/b_mux$out[10] ;
wire \dpath/b_mux$out[11] ;
wire \dpath/b_mux$out[12] ;
wire \dpath/b_mux$out[13] ;
wire \dpath/b_mux$out[14] ;
wire \dpath/b_mux$out[15] ;
wire \dpath/b_mux$out[1] ;
wire \dpath/b_mux$out[2] ;
wire \dpath/b_mux$out[3] ;
wire \dpath/b_mux$out[4] ;
wire \dpath/b_mux$out[5] ;
wire \dpath/b_mux$out[6] ;
wire \dpath/b_mux$out[7] ;
wire \dpath/b_mux$out[8] ;
wire \dpath/b_mux$out[9] ;
wire \dpath/a_lt_b/_000_ ;
wire \dpath/a_lt_b/_001_ ;
wire \dpath/a_lt_b/_002_ ;
wire \dpath/a_lt_b/_003_ ;
wire \dpath/a_lt_b/_004_ ;
wire \dpath/a_lt_b/_005_ ;
wire \dpath/a_lt_b/_006_ ;
wire \dpath/a_lt_b/_007_ ;
wire \dpath/a_lt_b/_008_ ;
wire \dpath/a_lt_b/_009_ ;
wire \dpath/a_lt_b/_010_ ;
wire \dpath/a_lt_b/_011_ ;
wire \dpath/a_lt_b/_012_ ;
wire \dpath/a_lt_b/_013_ ;
wire \dpath/a_lt_b/_014_ ;
wire \dpath/a_lt_b/_015_ ;
wire \dpath/a_lt_b/_016_ ;
wire \dpath/a_lt_b/_017_ ;
wire \dpath/a_lt_b/_018_ ;
wire \dpath/a_lt_b/_019_ ;
wire \dpath/a_lt_b/_020_ ;
wire \dpath/a_lt_b/_021_ ;
wire \dpath/a_lt_b/_022_ ;
wire \dpath/a_lt_b/_023_ ;
wire \dpath/a_lt_b/_024_ ;
wire \dpath/a_lt_b/_025_ ;
wire \dpath/a_lt_b/_026_ ;
wire \dpath/a_lt_b/_027_ ;
wire \dpath/a_lt_b/_028_ ;
wire \dpath/a_lt_b/_029_ ;
wire \dpath/a_lt_b/_030_ ;
wire \dpath/a_lt_b/_031_ ;
wire \dpath/a_lt_b/_032_ ;
wire \dpath/a_lt_b/_033_ ;
wire \dpath/a_lt_b/_034_ ;
wire \dpath/a_lt_b/_035_ ;
wire \dpath/a_lt_b/_036_ ;
wire \dpath/a_lt_b/_037_ ;
wire \dpath/a_lt_b/_038_ ;
wire \dpath/a_lt_b/_039_ ;
wire \dpath/a_lt_b/_040_ ;
wire \dpath/a_lt_b/_041_ ;
wire \dpath/a_lt_b/_042_ ;
wire \dpath/a_lt_b/_043_ ;
wire \dpath/a_lt_b/_044_ ;
wire \dpath/a_lt_b/_045_ ;
wire \dpath/a_lt_b/_046_ ;
wire \dpath/a_lt_b/_047_ ;
wire \dpath/a_lt_b/_048_ ;
wire \dpath/a_lt_b/_049_ ;
wire \dpath/a_lt_b/_050_ ;
wire \dpath/a_lt_b/_051_ ;
wire \dpath/a_lt_b/_052_ ;
wire \dpath/a_lt_b/_053_ ;
wire \dpath/a_lt_b/_054_ ;
wire \dpath/a_lt_b/_055_ ;
wire \dpath/a_lt_b/_056_ ;
wire \dpath/a_lt_b/_057_ ;
wire \dpath/a_lt_b/_058_ ;
wire \dpath/a_lt_b/_059_ ;
wire \dpath/a_lt_b/_060_ ;
wire \dpath/a_lt_b/_061_ ;
wire \dpath/a_lt_b/_062_ ;
wire \dpath/a_lt_b/_063_ ;
wire \dpath/a_lt_b/_064_ ;
wire \dpath/a_lt_b/_065_ ;
wire \dpath/a_lt_b/_066_ ;
wire \dpath/a_lt_b/_067_ ;
wire \dpath/a_lt_b/_068_ ;
wire \dpath/a_lt_b/_069_ ;
wire \dpath/a_lt_b/_070_ ;
wire \dpath/a_lt_b/_071_ ;
wire \dpath/a_lt_b/_072_ ;
wire \dpath/a_lt_b/_073_ ;
wire \dpath/a_lt_b/_074_ ;
wire \dpath/a_lt_b/_075_ ;
wire \dpath/a_lt_b/_076_ ;
wire \dpath/a_lt_b/_077_ ;
wire \dpath/a_lt_b/_078_ ;
wire \dpath/a_lt_b/_079_ ;
wire \dpath/a_lt_b/_080_ ;
wire \dpath/a_lt_b/_081_ ;
wire \dpath/a_lt_b/_082_ ;
wire \dpath/a_lt_b/_083_ ;
wire \dpath/a_lt_b/_084_ ;
wire \dpath/a_lt_b/_085_ ;
wire \dpath/a_lt_b/_086_ ;
wire \dpath/a_lt_b/_087_ ;
wire \dpath/a_lt_b/_088_ ;
wire \dpath/a_lt_b/_089_ ;
wire \dpath/a_mux/_000_ ;
wire \dpath/a_mux/_001_ ;
wire \dpath/a_mux/_002_ ;
wire \dpath/a_mux/_003_ ;
wire \dpath/a_mux/_004_ ;
wire \dpath/a_mux/_005_ ;
wire \dpath/a_mux/_006_ ;
wire \dpath/a_mux/_007_ ;
wire \dpath/a_mux/_008_ ;
wire \dpath/a_mux/_009_ ;
wire \dpath/a_mux/_010_ ;
wire \dpath/a_mux/_011_ ;
wire \dpath/a_mux/_012_ ;
wire \dpath/a_mux/_013_ ;
wire \dpath/a_mux/_014_ ;
wire \dpath/a_mux/_015_ ;
wire \dpath/a_mux/_016_ ;
wire \dpath/a_mux/_017_ ;
wire \dpath/a_mux/_018_ ;
wire \dpath/a_mux/_019_ ;
wire \dpath/a_mux/_020_ ;
wire \dpath/a_mux/_021_ ;
wire \dpath/a_mux/_022_ ;
wire \dpath/a_mux/_023_ ;
wire \dpath/a_mux/_024_ ;
wire \dpath/a_mux/_025_ ;
wire \dpath/a_mux/_026_ ;
wire \dpath/a_mux/_027_ ;
wire \dpath/a_mux/_028_ ;
wire \dpath/a_mux/_029_ ;
wire \dpath/a_mux/_030_ ;
wire \dpath/a_mux/_031_ ;
wire \dpath/a_mux/_032_ ;
wire \dpath/a_mux/_033_ ;
wire \dpath/a_mux/_034_ ;
wire \dpath/a_mux/_035_ ;
wire \dpath/a_mux/_036_ ;
wire \dpath/a_mux/_037_ ;
wire \dpath/a_mux/_038_ ;
wire \dpath/a_mux/_039_ ;
wire \dpath/a_mux/_040_ ;
wire \dpath/a_mux/_041_ ;
wire \dpath/a_mux/_042_ ;
wire \dpath/a_mux/_043_ ;
wire \dpath/a_mux/_044_ ;
wire \dpath/a_mux/_045_ ;
wire \dpath/a_mux/_046_ ;
wire \dpath/a_mux/_047_ ;
wire \dpath/a_mux/_048_ ;
wire \dpath/a_mux/_049_ ;
wire \dpath/a_mux/_050_ ;
wire \dpath/a_mux/_051_ ;
wire \dpath/a_mux/_052_ ;
wire \dpath/a_mux/_053_ ;
wire \dpath/a_mux/_054_ ;
wire \dpath/a_mux/_055_ ;
wire \dpath/a_mux/_056_ ;
wire \dpath/a_mux/_057_ ;
wire \dpath/a_mux/_058_ ;
wire \dpath/a_mux/_059_ ;
wire \dpath/a_mux/_060_ ;
wire \dpath/a_mux/_061_ ;
wire \dpath/a_mux/_062_ ;
wire \dpath/a_mux/_063_ ;
wire \dpath/a_mux/_064_ ;
wire \dpath/a_mux/_065_ ;
wire \dpath/a_mux/_066_ ;
wire \dpath/a_mux/_067_ ;
wire \dpath/a_mux/_068_ ;
wire \dpath/a_mux/_069_ ;
wire \dpath/a_mux/_070_ ;
wire \dpath/a_mux/_071_ ;
wire \dpath/a_mux/_072_ ;
wire \dpath/a_mux/_073_ ;
wire \dpath/a_mux/_074_ ;
wire \dpath/a_mux/_075_ ;
wire \dpath/a_mux/_076_ ;
wire \dpath/a_mux/_077_ ;
wire \dpath/a_mux/_078_ ;
wire \dpath/a_mux/_079_ ;
wire \dpath/a_mux/_080_ ;
wire \dpath/a_mux/_081_ ;
wire \dpath/a_mux/_082_ ;
wire \dpath/a_mux/_083_ ;
wire \dpath/a_mux/_084_ ;
wire \dpath/a_mux/_085_ ;
wire \dpath/a_mux/_086_ ;
wire \dpath/a_mux/_087_ ;
wire \dpath/a_mux/_088_ ;
wire \dpath/a_mux/_089_ ;
wire \dpath/a_mux/_090_ ;
wire \dpath/a_mux/_091_ ;
wire \dpath/a_mux/_092_ ;
wire \dpath/a_mux/_093_ ;
wire \dpath/a_mux/_094_ ;
wire \dpath/a_mux/_095_ ;
wire \dpath/a_mux/_096_ ;
wire \dpath/a_mux/_097_ ;
wire \dpath/a_mux/_098_ ;
wire \dpath/a_mux/_099_ ;
wire \dpath/a_mux/_100_ ;
wire \dpath/a_mux/_101_ ;
wire \dpath/a_mux/_102_ ;
wire \dpath/a_mux/_103_ ;
wire \dpath/a_reg/_000_ ;
wire \dpath/a_reg/_001_ ;
wire \dpath/a_reg/_002_ ;
wire \dpath/a_reg/_003_ ;
wire \dpath/a_reg/_004_ ;
wire \dpath/a_reg/_005_ ;
wire \dpath/a_reg/_006_ ;
wire \dpath/a_reg/_007_ ;
wire \dpath/a_reg/_008_ ;
wire \dpath/a_reg/_009_ ;
wire \dpath/a_reg/_010_ ;
wire \dpath/a_reg/_011_ ;
wire \dpath/a_reg/_012_ ;
wire \dpath/a_reg/_013_ ;
wire \dpath/a_reg/_014_ ;
wire \dpath/a_reg/_015_ ;
wire \dpath/a_reg/_016_ ;
wire \dpath/a_reg/_017_ ;
wire \dpath/a_reg/_018_ ;
wire \dpath/a_reg/_019_ ;
wire \dpath/a_reg/_020_ ;
wire \dpath/a_reg/_021_ ;
wire \dpath/a_reg/_022_ ;
wire \dpath/a_reg/_023_ ;
wire \dpath/a_reg/_024_ ;
wire \dpath/a_reg/_025_ ;
wire \dpath/a_reg/_026_ ;
wire \dpath/a_reg/_027_ ;
wire \dpath/a_reg/_028_ ;
wire \dpath/a_reg/_029_ ;
wire \dpath/a_reg/_030_ ;
wire \dpath/a_reg/_031_ ;
wire \dpath/a_reg/_032_ ;
wire \dpath/a_reg/_033_ ;
wire \dpath/a_reg/_034_ ;
wire \dpath/a_reg/_035_ ;
wire \dpath/a_reg/_036_ ;
wire \dpath/a_reg/_037_ ;
wire \dpath/a_reg/_038_ ;
wire \dpath/a_reg/_039_ ;
wire \dpath/a_reg/_040_ ;
wire \dpath/a_reg/_041_ ;
wire \dpath/a_reg/_042_ ;
wire \dpath/a_reg/_043_ ;
wire \dpath/a_reg/_044_ ;
wire \dpath/a_reg/_045_ ;
wire \dpath/a_reg/_046_ ;
wire \dpath/a_reg/_047_ ;
wire \dpath/a_reg/_048_ ;
wire \dpath/a_reg/_049_ ;
wire \dpath/a_reg/_050_ ;
wire \dpath/a_reg/_051_ ;
wire \dpath/a_reg/_052_ ;
wire \dpath/a_reg/_053_ ;
wire \dpath/a_reg/_054_ ;
wire \dpath/a_reg/_055_ ;
wire \dpath/a_reg/_056_ ;
wire \dpath/a_reg/_057_ ;
wire \dpath/a_reg/_058_ ;
wire \dpath/a_reg/_059_ ;
wire \dpath/a_reg/_060_ ;
wire \dpath/a_reg/_061_ ;
wire \dpath/a_reg/_062_ ;
wire \dpath/a_reg/_063_ ;
wire \dpath/a_reg/_064_ ;
wire \dpath/a_reg/_065_ ;
wire \dpath/b_mux/_000_ ;
wire \dpath/b_mux/_001_ ;
wire \dpath/b_mux/_002_ ;
wire \dpath/b_mux/_003_ ;
wire \dpath/b_mux/_004_ ;
wire \dpath/b_mux/_005_ ;
wire \dpath/b_mux/_006_ ;
wire \dpath/b_mux/_007_ ;
wire \dpath/b_mux/_008_ ;
wire \dpath/b_mux/_009_ ;
wire \dpath/b_mux/_010_ ;
wire \dpath/b_mux/_011_ ;
wire \dpath/b_mux/_012_ ;
wire \dpath/b_mux/_013_ ;
wire \dpath/b_mux/_014_ ;
wire \dpath/b_mux/_015_ ;
wire \dpath/b_mux/_016_ ;
wire \dpath/b_mux/_017_ ;
wire \dpath/b_mux/_018_ ;
wire \dpath/b_mux/_019_ ;
wire \dpath/b_mux/_020_ ;
wire \dpath/b_mux/_021_ ;
wire \dpath/b_mux/_022_ ;
wire \dpath/b_mux/_023_ ;
wire \dpath/b_mux/_024_ ;
wire \dpath/b_mux/_025_ ;
wire \dpath/b_mux/_026_ ;
wire \dpath/b_mux/_027_ ;
wire \dpath/b_mux/_028_ ;
wire \dpath/b_mux/_029_ ;
wire \dpath/b_mux/_030_ ;
wire \dpath/b_mux/_031_ ;
wire \dpath/b_mux/_032_ ;
wire \dpath/b_mux/_033_ ;
wire \dpath/b_mux/_034_ ;
wire \dpath/b_mux/_035_ ;
wire \dpath/b_mux/_036_ ;
wire \dpath/b_mux/_037_ ;
wire \dpath/b_mux/_038_ ;
wire \dpath/b_mux/_039_ ;
wire \dpath/b_mux/_040_ ;
wire \dpath/b_mux/_041_ ;
wire \dpath/b_mux/_042_ ;
wire \dpath/b_mux/_043_ ;
wire \dpath/b_mux/_044_ ;
wire \dpath/b_mux/_045_ ;
wire \dpath/b_mux/_046_ ;
wire \dpath/b_mux/_047_ ;
wire \dpath/b_mux/_048_ ;
wire \dpath/b_mux/_049_ ;
wire \dpath/b_reg/_000_ ;
wire \dpath/b_reg/_001_ ;
wire \dpath/b_reg/_002_ ;
wire \dpath/b_reg/_003_ ;
wire \dpath/b_reg/_004_ ;
wire \dpath/b_reg/_005_ ;
wire \dpath/b_reg/_006_ ;
wire \dpath/b_reg/_007_ ;
wire \dpath/b_reg/_008_ ;
wire \dpath/b_reg/_009_ ;
wire \dpath/b_reg/_010_ ;
wire \dpath/b_reg/_011_ ;
wire \dpath/b_reg/_012_ ;
wire \dpath/b_reg/_013_ ;
wire \dpath/b_reg/_014_ ;
wire \dpath/b_reg/_015_ ;
wire \dpath/b_reg/_016_ ;
wire \dpath/b_reg/_017_ ;
wire \dpath/b_reg/_018_ ;
wire \dpath/b_reg/_019_ ;
wire \dpath/b_reg/_020_ ;
wire \dpath/b_reg/_021_ ;
wire \dpath/b_reg/_022_ ;
wire \dpath/b_reg/_023_ ;
wire \dpath/b_reg/_024_ ;
wire \dpath/b_reg/_025_ ;
wire \dpath/b_reg/_026_ ;
wire \dpath/b_reg/_027_ ;
wire \dpath/b_reg/_028_ ;
wire \dpath/b_reg/_029_ ;
wire \dpath/b_reg/_030_ ;
wire \dpath/b_reg/_031_ ;
wire \dpath/b_reg/_032_ ;
wire \dpath/b_reg/_033_ ;
wire \dpath/b_reg/_034_ ;
wire \dpath/b_reg/_035_ ;
wire \dpath/b_reg/_036_ ;
wire \dpath/b_reg/_037_ ;
wire \dpath/b_reg/_038_ ;
wire \dpath/b_reg/_039_ ;
wire \dpath/b_reg/_040_ ;
wire \dpath/b_reg/_041_ ;
wire \dpath/b_reg/_042_ ;
wire \dpath/b_reg/_043_ ;
wire \dpath/b_reg/_044_ ;
wire \dpath/b_reg/_045_ ;
wire \dpath/b_reg/_046_ ;
wire \dpath/b_reg/_047_ ;
wire \dpath/b_reg/_048_ ;
wire \dpath/b_reg/_049_ ;
wire \dpath/b_reg/_050_ ;
wire \dpath/b_reg/_051_ ;
wire \dpath/b_reg/_052_ ;
wire \dpath/b_reg/_053_ ;
wire \dpath/b_reg/_054_ ;
wire \dpath/b_reg/_055_ ;
wire \dpath/b_reg/_056_ ;
wire \dpath/b_reg/_057_ ;
wire \dpath/b_reg/_058_ ;
wire \dpath/b_reg/_059_ ;
wire \dpath/b_reg/_060_ ;
wire \dpath/b_reg/_061_ ;
wire \dpath/b_reg/_062_ ;
wire \dpath/b_reg/_063_ ;
wire \dpath/b_reg/_064_ ;
wire \dpath/b_reg/_065_ ;
wire \dpath/b_zero/_00_ ;
wire \dpath/b_zero/_01_ ;
wire \dpath/b_zero/_02_ ;
wire \dpath/b_zero/_03_ ;
wire \dpath/b_zero/_04_ ;
wire \dpath/b_zero/_05_ ;
wire \dpath/b_zero/_06_ ;
wire \dpath/b_zero/_07_ ;
wire \dpath/b_zero/_08_ ;
wire \dpath/b_zero/_09_ ;
wire \dpath/b_zero/_10_ ;
wire \dpath/b_zero/_11_ ;
wire \dpath/b_zero/_12_ ;
wire \dpath/b_zero/_13_ ;
wire \dpath/b_zero/_14_ ;
wire \dpath/b_zero/_15_ ;
wire \dpath/b_zero/_16_ ;
wire \dpath/b_zero/_17_ ;
wire \dpath/b_zero/_18_ ;
wire \dpath/b_zero/_19_ ;
wire \dpath/b_zero/_20_ ;
wire \dpath/b_zero/_21_ ;
wire \dpath/b_zero/_22_ ;
wire \dpath/b_zero/_23_ ;
wire \dpath/b_zero/_24_ ;
wire \dpath/sub/_000_ ;
wire \dpath/sub/_001_ ;
wire \dpath/sub/_002_ ;
wire \dpath/sub/_003_ ;
wire \dpath/sub/_004_ ;
wire \dpath/sub/_005_ ;
wire \dpath/sub/_006_ ;
wire \dpath/sub/_007_ ;
wire \dpath/sub/_008_ ;
wire \dpath/sub/_009_ ;
wire \dpath/sub/_010_ ;
wire \dpath/sub/_011_ ;
wire \dpath/sub/_012_ ;
wire \dpath/sub/_013_ ;
wire \dpath/sub/_014_ ;
wire \dpath/sub/_015_ ;
wire \dpath/sub/_016_ ;
wire \dpath/sub/_017_ ;
wire \dpath/sub/_018_ ;
wire \dpath/sub/_019_ ;
wire \dpath/sub/_020_ ;
wire \dpath/sub/_021_ ;
wire \dpath/sub/_022_ ;
wire \dpath/sub/_023_ ;
wire \dpath/sub/_024_ ;
wire \dpath/sub/_025_ ;
wire \dpath/sub/_026_ ;
wire \dpath/sub/_027_ ;
wire \dpath/sub/_028_ ;
wire \dpath/sub/_029_ ;
wire \dpath/sub/_030_ ;
wire \dpath/sub/_031_ ;
wire \dpath/sub/_032_ ;
wire \dpath/sub/_033_ ;
wire \dpath/sub/_034_ ;
wire \dpath/sub/_035_ ;
wire \dpath/sub/_036_ ;
wire \dpath/sub/_037_ ;
wire \dpath/sub/_038_ ;
wire \dpath/sub/_039_ ;
wire \dpath/sub/_040_ ;
wire \dpath/sub/_041_ ;
wire \dpath/sub/_042_ ;
wire \dpath/sub/_043_ ;
wire \dpath/sub/_044_ ;
wire \dpath/sub/_045_ ;
wire \dpath/sub/_046_ ;
wire \dpath/sub/_047_ ;
wire \dpath/sub/_048_ ;
wire \dpath/sub/_049_ ;
wire \dpath/sub/_050_ ;
wire \dpath/sub/_051_ ;
wire \dpath/sub/_052_ ;
wire \dpath/sub/_053_ ;
wire \dpath/sub/_054_ ;
wire \dpath/sub/_055_ ;
wire \dpath/sub/_056_ ;
wire \dpath/sub/_057_ ;
wire \dpath/sub/_058_ ;
wire \dpath/sub/_059_ ;
wire \dpath/sub/_060_ ;
wire \dpath/sub/_061_ ;
wire \dpath/sub/_062_ ;
wire \dpath/sub/_063_ ;
wire \dpath/sub/_064_ ;
wire \dpath/sub/_065_ ;
wire \dpath/sub/_066_ ;
wire \dpath/sub/_067_ ;
wire \dpath/sub/_068_ ;
wire \dpath/sub/_069_ ;
wire \dpath/sub/_070_ ;
wire \dpath/sub/_071_ ;
wire \dpath/sub/_072_ ;
wire \dpath/sub/_073_ ;
wire \dpath/sub/_074_ ;
wire \dpath/sub/_075_ ;
wire \dpath/sub/_076_ ;
wire \dpath/sub/_077_ ;
wire \dpath/sub/_078_ ;
wire \dpath/sub/_079_ ;
wire \dpath/sub/_080_ ;
wire \dpath/sub/_081_ ;
wire \dpath/sub/_082_ ;
wire \dpath/sub/_083_ ;
wire \dpath/sub/_084_ ;
wire \dpath/sub/_085_ ;
wire \dpath/sub/_086_ ;
wire \dpath/sub/_087_ ;
wire \dpath/sub/_088_ ;
wire \dpath/sub/_089_ ;
wire \dpath/sub/_090_ ;
wire \dpath/sub/_091_ ;
wire \dpath/sub/_092_ ;
wire \dpath/sub/_093_ ;
wire \dpath/sub/_094_ ;
wire \dpath/sub/_095_ ;
wire \dpath/sub/_096_ ;
wire \dpath/sub/_097_ ;
wire \dpath/sub/_098_ ;
wire \dpath/sub/_099_ ;
wire \dpath/sub/_100_ ;
wire \dpath/sub/_101_ ;
wire \dpath/sub/_102_ ;
wire \dpath/sub/_103_ ;
wire \dpath/sub/_104_ ;
wire \dpath/sub/_105_ ;
wire \dpath/sub/_106_ ;
wire \dpath/sub/_107_ ;
wire \dpath/sub/_108_ ;
wire \dpath/sub/_109_ ;
wire \dpath/sub/_110_ ;
wire \dpath/sub/_111_ ;
wire \dpath/sub/_112_ ;
wire \dpath/sub/_113_ ;
wire \dpath/sub/_114_ ;
wire \dpath/sub/_115_ ;
wire \dpath/sub/_116_ ;
wire \dpath/sub/_117_ ;
wire \dpath/sub/_118_ ;
wire \dpath/sub/_119_ ;
wire \dpath/sub/_120_ ;
wire req_rdy ;
wire resp_val ;
wire req_val ;
wire resp_rdy ;
wire reset ;
wire clk ;
wire \resp_msg[0] ;
wire \req_msg[16] ;
wire \resp_msg[1] ;
wire \req_msg[17] ;
wire \resp_msg[2] ;
wire \req_msg[18] ;
wire \resp_msg[3] ;
wire \req_msg[19] ;
wire \resp_msg[4] ;
wire \req_msg[20] ;
wire \resp_msg[5] ;
wire \req_msg[21] ;
wire \resp_msg[6] ;
wire \req_msg[22] ;
wire \resp_msg[7] ;
wire \req_msg[23] ;
wire \resp_msg[8] ;
wire \req_msg[24] ;
wire \resp_msg[9] ;
wire \req_msg[25] ;
wire \resp_msg[10] ;
wire \req_msg[26] ;
wire \resp_msg[11] ;
wire \req_msg[27] ;
wire \resp_msg[12] ;
wire \req_msg[28] ;
wire \resp_msg[13] ;
wire \req_msg[29] ;
wire \resp_msg[14] ;
wire \req_msg[30] ;
wire \resp_msg[15] ;
wire \req_msg[31] ;
wire \req_msg[0] ;
wire \req_msg[1] ;
wire \req_msg[2] ;
wire \req_msg[3] ;
wire \req_msg[4] ;
wire \req_msg[5] ;
wire \req_msg[6] ;
wire \req_msg[7] ;
wire \req_msg[8] ;
wire \req_msg[9] ;
wire \req_msg[10] ;
wire \req_msg[11] ;
wire \req_msg[12] ;
wire \req_msg[13] ;
wire \req_msg[14] ;
wire \req_msg[15] ;
wire clk_86 ;
wire clk_85 ;
wire clk_84 ;
wire clk_83 ;
wire clk_82 ;
wire clk_81 ;
wire clk_80 ;
wire clk_79 ;
wire clk_78 ;
wire clk_77 ;
wire clk_76 ;
wire clk_75 ;
wire clk_74 ;
wire clk_73 ;
wire clk_72 ;
wire clk_71 ;
wire clk_70 ;
wire clk_69 ;
wire clk_68 ;
wire clk_67 ;
wire clk_66 ;
wire clk_65 ;
wire clk_64 ;
wire clk_63 ;
wire clk_62 ;
wire clk_61 ;
wire clk_60 ;
wire clk_59 ;
wire clk_58 ;
wire clk_57 ;
wire clk_56 ;
wire clk_55 ;
wire clk_54 ;
wire clk_53 ;
wire clk_52 ;
wire clk_51 ;
wire clk_50 ;
wire clk_49 ;
wire clk_48 ;
wire clk_47 ;
wire clk_46 ;
wire clk_45 ;
wire clk_44 ;
wire clk_43 ;
wire clk_42 ;
wire clk_41 ;
wire clk_40 ;
wire clk_39 ;
wire clk_38 ;
wire clk_37 ;
wire clk_36 ;
wire clk_35 ;
wire clk_34 ;
wire clk_33 ;
wire clk_32 ;
wire clk_31 ;
wire clk_30 ;
wire clk_29 ;
wire clk_28 ;
wire clk_27 ;
wire clk_26 ;
wire clk_25 ;
wire clk_24 ;
wire clk_23 ;
wire clk_22 ;
wire clk_21 ;
wire clk_20 ;
wire clk_19 ;
wire clk_18 ;
wire clk_17 ;
wire clk_16 ;
wire clk_15 ;
wire clk_14 ;
wire clk_13 ;
wire clk_12 ;
wire clk_11 ;
wire clk_10 ;
wire clk_9 ;
wire clk_8 ;
wire clk_7 ;
wire clk_6 ;
wire clk_5 ;
wire clk_4 ;
wire clk_3 ;
wire clk_2 ;
wire clk_1 ;
wire clk_0 ;

sky130_fd_sc_hs__nor2_1 \ctrl/_17_ ( .A(\ctrl/_05_ ), .B(\ctrl/_06_ ), .Y(\ctrl/_03_ ) );
sky130_fd_sc_hs__and2b_1 \ctrl/_18_ ( .A_N(\ctrl/_05_ ), .B(\ctrl/_06_ ), .X(\ctrl/_16_ ) );
sky130_fd_sc_hs__nor3b_1 \ctrl/_19_ ( .A(\ctrl/_06_ ), .B(\ctrl/_07_ ), .C_N(\ctrl/_05_ ), .Y(\ctrl/_00_ ) );
sky130_fd_sc_hs__and3b_1 \ctrl/_20_ ( .A_N(\ctrl/_06_ ), .B(\ctrl/_05_ ), .C(\ctrl/_07_ ), .X(\ctrl/_01_ ) );
sky130_fd_sc_hs__nor3b_1 \ctrl/_21_ ( .A(\ctrl/_05_ ), .B(\ctrl/_06_ ), .C_N(\ctrl/_14_ ), .Y(\ctrl/_09_ ) );
sky130_fd_sc_hs__nor2b_4 \ctrl/_22_ ( .A(\ctrl/_07_ ), .B_N(\ctrl/_08_ ), .Y(\ctrl/_10_ ) );
sky130_fd_sc_hs__inv_1 \ctrl/_23_ ( .A(\ctrl/_06_ ), .Y(\ctrl/_02_ ) );
sky130_fd_sc_hs__nand3_2 \ctrl/_24_ ( .A(\ctrl/_10_ ), .B(\ctrl/_05_ ), .C(\ctrl/_02_ ), .Y(\ctrl/_11_ ) );
sky130_fd_sc_hs__o21a_1 \ctrl/_25_ ( .A1(\ctrl/_05_ ), .A2(\ctrl/_09_ ), .B1(\ctrl/_11_ ), .X(\ctrl/_12_ ) );
sky130_fd_sc_hs__a22oi_1 \ctrl/_26_ ( .A1(\ctrl/_15_ ), .A2(\ctrl/_16_ ), .B1(\ctrl/_11_ ), .B2(\ctrl/_02_ ), .Y(\ctrl/_13_ ) );
sky130_fd_sc_hs__o21bai_1 \ctrl/_27_ ( .A1(\ctrl/_05_ ), .A2(\ctrl/_06_ ), .B1_N(\ctrl/_01_ ), .Y(\ctrl/_04_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/_28_ ( .A(ctrl$b_mux_sel ), .X(req_rdy ) );
sky130_fd_sc_hs__buf_1 \ctrl/_29_ ( .A(\ctrl/curr_state__0[0] ), .X(\ctrl/_05_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/_30_ ( .A(\ctrl/curr_state__0[1] ), .X(\ctrl/_06_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/_31_ ( .A(\ctrl/_03_ ), .X(ctrl$b_mux_sel ) );
sky130_fd_sc_hs__buf_1 \ctrl/_32_ ( .A(\ctrl/_16_ ), .X(resp_val ) );
sky130_fd_sc_hs__buf_1 \ctrl/_33_ ( .A(ctrl$is_a_lt_b ), .X(\ctrl/_07_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/_34_ ( .A(\ctrl/_00_ ), .X(\ctrl$a_mux_sel[0] ) );
sky130_fd_sc_hs__buf_1 \ctrl/_35_ ( .A(\ctrl/_01_ ), .X(\ctrl$a_mux_sel[1] ) );
sky130_fd_sc_hs__buf_1 \ctrl/_36_ ( .A(req_val ), .X(\ctrl/_14_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/_37_ ( .A(ctrl$is_b_zero ), .X(\ctrl/_08_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/_38_ ( .A(resp_rdy ), .X(\ctrl/_15_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/_39_ ( .A(\ctrl/_12_ ), .X(\ctrl/next_state__0[0] ) );
sky130_fd_sc_hs__buf_1 \ctrl/_40_ ( .A(\ctrl/_13_ ), .X(\ctrl/next_state__0[1] ) );
sky130_fd_sc_hs__buf_1 \ctrl/_41_ ( .A(\ctrl/_04_ ), .X(ctrl$b_reg_en ) );
sky130_fd_sc_hs__buf_1 \ctrl/_42_ ( .A(\ctrl/_02_ ), .X(ctrl$a_reg_en ) );
sky130_fd_sc_hs__nor2b_2 \ctrl/state/_07_ ( .A(\ctrl/state/_06_ ), .B_N(\ctrl/state/_04_ ), .Y(\ctrl/state/_02_ ) );
sky130_fd_sc_hs__nor2b_2 \ctrl/state/_08_ ( .A(\ctrl/state/_06_ ), .B_N(\ctrl/state/_05_ ), .Y(\ctrl/state/_03_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/state/_09_ ( .A(\ctrl/next_state__0[0] ), .X(\ctrl/state/_04_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/state/_10_ ( .A(reset ), .X(\ctrl/state/_06_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/state/_11_ ( .A(\ctrl/state/_02_ ), .X(\ctrl/state/_00_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/state/_12_ ( .A(\ctrl/next_state__0[1] ), .X(\ctrl/state/_05_ ) );
sky130_fd_sc_hs__buf_1 \ctrl/state/_13_ ( .A(\ctrl/state/_03_ ), .X(\ctrl/state/_01_ ) );
sky130_fd_sc_hs__dfxtp_1 \ctrl/state/_14_ ( .D(\ctrl/state/_00_ ), .Q(\ctrl/curr_state__0[0] ), .CLK(clk_85 ) );
sky130_fd_sc_hs__dfxtp_1 \ctrl/state/_15_ ( .D(\ctrl/state/_01_ ), .Q(\ctrl/curr_state__0[1] ), .CLK(clk_85 ) );
sky130_fd_sc_hs__nor2b_2 \dpath/a_lt_b/_090_ ( .A(\dpath/a_lt_b/_025_ ), .B_N(\dpath/a_lt_b/_009_ ), .Y(\dpath/a_lt_b/_032_ ) );
sky130_fd_sc_hs__nand2b_2 \dpath/a_lt_b/_091_ ( .A_N(\dpath/a_lt_b/_009_ ), .B(\dpath/a_lt_b/_025_ ), .Y(\dpath/a_lt_b/_033_ ) );
sky130_fd_sc_hs__and3b_1 \dpath/a_lt_b/_092_ ( .A_N(\dpath/a_lt_b/_024_ ), .B(\dpath/a_lt_b/_033_ ), .C(\dpath/a_lt_b/_008_ ), .X(\dpath/a_lt_b/_034_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/a_lt_b/_093_ ( .A(\dpath/a_lt_b/_024_ ), .B(\dpath/a_lt_b/_008_ ), .Y(\dpath/a_lt_b/_035_ ) );
sky130_fd_sc_hs__and3b_1 \dpath/a_lt_b/_094_ ( .A_N(\dpath/a_lt_b/_032_ ), .B(\dpath/a_lt_b/_035_ ), .C(\dpath/a_lt_b/_033_ ), .X(\dpath/a_lt_b/_036_ ) );
sky130_fd_sc_hs__inv_8 \dpath/a_lt_b/_095_ ( .A(\dpath/a_lt_b/_023_ ), .Y(\dpath/a_lt_b/_037_ ) );
sky130_fd_sc_hs__nand2b_4 \dpath/a_lt_b/_096_ ( .A_N(\dpath/a_lt_b/_000_ ), .B(\dpath/a_lt_b/_016_ ), .Y(\dpath/a_lt_b/_038_ ) );
sky130_fd_sc_hs__maj3_1 \dpath/a_lt_b/_097_ ( .A(\dpath/a_lt_b/_037_ ), .B(\dpath/a_lt_b/_038_ ), .C(\dpath/a_lt_b/_007_ ), .X(\dpath/a_lt_b/_039_ ) );
sky130_fd_sc_hs__and2_1 \dpath/a_lt_b/_098_ ( .A(\dpath/a_lt_b/_036_ ), .B(\dpath/a_lt_b/_039_ ), .X(\dpath/a_lt_b/_040_ ) );
sky130_fd_sc_hs__inv_1 \dpath/a_lt_b/_099_ ( .A(\dpath/a_lt_b/_026_ ), .Y(\dpath/a_lt_b/_041_ ) );
sky130_fd_sc_hs__nor2b_1 \dpath/a_lt_b/_100_ ( .A(\dpath/a_lt_b/_027_ ), .B_N(\dpath/a_lt_b/_011_ ), .Y(\dpath/a_lt_b/_042_ ) );
sky130_fd_sc_hs__a21o_1 \dpath/a_lt_b/_101_ ( .A1(\dpath/a_lt_b/_010_ ), .A2(\dpath/a_lt_b/_041_ ), .B1(\dpath/a_lt_b/_042_ ), .X(\dpath/a_lt_b/_043_ ) );
sky130_fd_sc_hs__nor2b_4 \dpath/a_lt_b/_102_ ( .A(\dpath/a_lt_b/_013_ ), .B_N(\dpath/a_lt_b/_029_ ), .Y(\dpath/a_lt_b/_044_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/a_lt_b/_103_ ( .A(\dpath/a_lt_b/_028_ ), .B(\dpath/a_lt_b/_012_ ), .Y(\dpath/a_lt_b/_045_ ) );
sky130_fd_sc_hs__nand2b_1 \dpath/a_lt_b/_104_ ( .A_N(\dpath/a_lt_b/_029_ ), .B(\dpath/a_lt_b/_013_ ), .Y(\dpath/a_lt_b/_046_ ) );
sky130_fd_sc_hs__and3b_1 \dpath/a_lt_b/_105_ ( .A_N(\dpath/a_lt_b/_044_ ), .B(\dpath/a_lt_b/_045_ ), .C(\dpath/a_lt_b/_046_ ), .X(\dpath/a_lt_b/_047_ ) );
sky130_fd_sc_hs__nor2b_4 \dpath/a_lt_b/_106_ ( .A(\dpath/a_lt_b/_011_ ), .B_N(\dpath/a_lt_b/_027_ ), .Y(\dpath/a_lt_b/_048_ ) );
sky130_fd_sc_hs__o21ba_1 \dpath/a_lt_b/_107_ ( .A1(\dpath/a_lt_b/_010_ ), .A2(\dpath/a_lt_b/_041_ ), .B1_N(\dpath/a_lt_b/_048_ ), .X(\dpath/a_lt_b/_049_ ) );
sky130_fd_sc_hs__and3b_1 \dpath/a_lt_b/_108_ ( .A_N(\dpath/a_lt_b/_043_ ), .B(\dpath/a_lt_b/_047_ ), .C(\dpath/a_lt_b/_049_ ), .X(\dpath/a_lt_b/_050_ ) );
sky130_fd_sc_hs__o31ai_1 \dpath/a_lt_b/_109_ ( .A1(\dpath/a_lt_b/_032_ ), .A2(\dpath/a_lt_b/_034_ ), .A3(\dpath/a_lt_b/_040_ ), .B1(\dpath/a_lt_b/_050_ ), .Y(\dpath/a_lt_b/_051_ ) );
sky130_fd_sc_hs__nor2b_2 \dpath/a_lt_b/_110_ ( .A(\dpath/a_lt_b/_028_ ), .B_N(\dpath/a_lt_b/_012_ ), .Y(\dpath/a_lt_b/_052_ ) );
sky130_fd_sc_hs__nor2b_1 \dpath/a_lt_b/_111_ ( .A(\dpath/a_lt_b/_052_ ), .B_N(\dpath/a_lt_b/_046_ ), .Y(\dpath/a_lt_b/_053_ ) );
sky130_fd_sc_hs__or2_1 \dpath/a_lt_b/_112_ ( .A(\dpath/a_lt_b/_044_ ), .B(\dpath/a_lt_b/_053_ ), .X(\dpath/a_lt_b/_054_ ) );
sky130_fd_sc_hs__nand3b_1 \dpath/a_lt_b/_113_ ( .A_N(\dpath/a_lt_b/_048_ ), .B(\dpath/a_lt_b/_047_ ), .C(\dpath/a_lt_b/_043_ ), .Y(\dpath/a_lt_b/_055_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/a_lt_b/_114_ ( .A(\dpath/a_lt_b/_020_ ), .B_N(\dpath/a_lt_b/_004_ ), .X(\dpath/a_lt_b/_056_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/a_lt_b/_115_ ( .A(\dpath/a_lt_b/_019_ ), .B_N(\dpath/a_lt_b/_003_ ), .X(\dpath/a_lt_b/_057_ ) );
sky130_fd_sc_hs__nand2_2 \dpath/a_lt_b/_116_ ( .A(\dpath/a_lt_b/_056_ ), .B(\dpath/a_lt_b/_057_ ), .Y(\dpath/a_lt_b/_058_ ) );
sky130_fd_sc_hs__and2b_2 \dpath/a_lt_b/_117_ ( .A_N(\dpath/a_lt_b/_005_ ), .B(\dpath/a_lt_b/_021_ ), .X(\dpath/a_lt_b/_059_ ) );
sky130_fd_sc_hs__nor2b_2 \dpath/a_lt_b/_118_ ( .A(\dpath/a_lt_b/_006_ ), .B_N(\dpath/a_lt_b/_022_ ), .Y(\dpath/a_lt_b/_060_ ) );
sky130_fd_sc_hs__nand2b_2 \dpath/a_lt_b/_119_ ( .A_N(\dpath/a_lt_b/_021_ ), .B(\dpath/a_lt_b/_005_ ), .Y(\dpath/a_lt_b/_061_ ) );
sky130_fd_sc_hs__nand2b_4 \dpath/a_lt_b/_120_ ( .A_N(\dpath/a_lt_b/_022_ ), .B(\dpath/a_lt_b/_006_ ), .Y(\dpath/a_lt_b/_062_ ) );
sky130_fd_sc_hs__nand3b_1 \dpath/a_lt_b/_121_ ( .A_N(\dpath/a_lt_b/_060_ ), .B(\dpath/a_lt_b/_061_ ), .C(\dpath/a_lt_b/_062_ ), .Y(\dpath/a_lt_b/_063_ ) );
sky130_fd_sc_hs__nor2_2 \dpath/a_lt_b/_122_ ( .A(\dpath/a_lt_b/_059_ ), .B(\dpath/a_lt_b/_063_ ), .Y(\dpath/a_lt_b/_064_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/a_lt_b/_123_ ( .A(\dpath/a_lt_b/_004_ ), .B_N(\dpath/a_lt_b/_020_ ), .X(\dpath/a_lt_b/_065_ ) );
sky130_fd_sc_hs__or2b_4 \dpath/a_lt_b/_124_ ( .A(\dpath/a_lt_b/_003_ ), .B_N(\dpath/a_lt_b/_019_ ), .X(\dpath/a_lt_b/_066_ ) );
sky130_fd_sc_hs__nand3_2 \dpath/a_lt_b/_125_ ( .A(\dpath/a_lt_b/_064_ ), .B(\dpath/a_lt_b/_065_ ), .C(\dpath/a_lt_b/_066_ ), .Y(\dpath/a_lt_b/_067_ ) );
sky130_fd_sc_hs__or2_1 \dpath/a_lt_b/_126_ ( .A(\dpath/a_lt_b/_058_ ), .B(\dpath/a_lt_b/_067_ ), .X(\dpath/a_lt_b/_068_ ) );
sky130_fd_sc_hs__inv_1 \dpath/a_lt_b/_127_ ( .A(\dpath/a_lt_b/_001_ ), .Y(\dpath/a_lt_b/_069_ ) );
sky130_fd_sc_hs__nor2b_4 \dpath/a_lt_b/_128_ ( .A(\dpath/a_lt_b/_018_ ), .B_N(\dpath/a_lt_b/_002_ ), .Y(\dpath/a_lt_b/_070_ ) );
sky130_fd_sc_hs__nor2b_4 \dpath/a_lt_b/_129_ ( .A(\dpath/a_lt_b/_017_ ), .B_N(\dpath/a_lt_b/_001_ ), .Y(\dpath/a_lt_b/_071_ ) );
sky130_fd_sc_hs__nor2b_2 \dpath/a_lt_b/_130_ ( .A(\dpath/a_lt_b/_002_ ), .B_N(\dpath/a_lt_b/_018_ ), .Y(\dpath/a_lt_b/_072_ ) );
sky130_fd_sc_hs__or3_1 \dpath/a_lt_b/_131_ ( .A(\dpath/a_lt_b/_070_ ), .B(\dpath/a_lt_b/_071_ ), .C(\dpath/a_lt_b/_072_ ), .X(\dpath/a_lt_b/_073_ ) );
sky130_fd_sc_hs__a21oi_4 \dpath/a_lt_b/_132_ ( .A1(\dpath/a_lt_b/_017_ ), .A2(\dpath/a_lt_b/_069_ ), .B1(\dpath/a_lt_b/_073_ ), .Y(\dpath/a_lt_b/_074_ ) );
sky130_fd_sc_hs__and2b_2 \dpath/a_lt_b/_133_ ( .A_N(\dpath/a_lt_b/_015_ ), .B(\dpath/a_lt_b/_031_ ), .X(\dpath/a_lt_b/_075_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/a_lt_b/_134_ ( .A(\dpath/a_lt_b/_014_ ), .B(\dpath/a_lt_b/_030_ ), .Y(\dpath/a_lt_b/_076_ ) );
sky130_fd_sc_hs__or2b_2 \dpath/a_lt_b/_135_ ( .A(\dpath/a_lt_b/_031_ ), .B_N(\dpath/a_lt_b/_015_ ), .X(\dpath/a_lt_b/_077_ ) );
sky130_fd_sc_hs__and3b_1 \dpath/a_lt_b/_136_ ( .A_N(\dpath/a_lt_b/_075_ ), .B(\dpath/a_lt_b/_076_ ), .C(\dpath/a_lt_b/_077_ ), .X(\dpath/a_lt_b/_078_ ) );
sky130_fd_sc_hs__nand3b_1 \dpath/a_lt_b/_137_ ( .A_N(\dpath/a_lt_b/_068_ ), .B(\dpath/a_lt_b/_074_ ), .C(\dpath/a_lt_b/_078_ ), .Y(\dpath/a_lt_b/_079_ ) );
sky130_fd_sc_hs__a31o_1 \dpath/a_lt_b/_138_ ( .A1(\dpath/a_lt_b/_051_ ), .A2(\dpath/a_lt_b/_054_ ), .A3(\dpath/a_lt_b/_055_ ), .B1(\dpath/a_lt_b/_079_ ), .X(\dpath/a_lt_b/_080_ ) );
sky130_fd_sc_hs__nor3b_1 \dpath/a_lt_b/_139_ ( .A(\dpath/a_lt_b/_070_ ), .B(\dpath/a_lt_b/_072_ ), .C_N(\dpath/a_lt_b/_071_ ), .Y(\dpath/a_lt_b/_081_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/a_lt_b/_140_ ( .A(\dpath/a_lt_b/_030_ ), .B_N(\dpath/a_lt_b/_014_ ), .X(\dpath/a_lt_b/_082_ ) );
sky130_fd_sc_hs__a21oi_1 \dpath/a_lt_b/_141_ ( .A1(\dpath/a_lt_b/_077_ ), .A2(\dpath/a_lt_b/_082_ ), .B1(\dpath/a_lt_b/_075_ ), .Y(\dpath/a_lt_b/_083_ ) );
sky130_fd_sc_hs__and2_1 \dpath/a_lt_b/_142_ ( .A(\dpath/a_lt_b/_074_ ), .B(\dpath/a_lt_b/_083_ ), .X(\dpath/a_lt_b/_084_ ) );
sky130_fd_sc_hs__nor2_1 \dpath/a_lt_b/_143_ ( .A(\dpath/a_lt_b/_058_ ), .B(\dpath/a_lt_b/_067_ ), .Y(\dpath/a_lt_b/_085_ ) );
sky130_fd_sc_hs__o31ai_1 \dpath/a_lt_b/_144_ ( .A1(\dpath/a_lt_b/_070_ ), .A2(\dpath/a_lt_b/_081_ ), .A3(\dpath/a_lt_b/_084_ ), .B1(\dpath/a_lt_b/_085_ ), .Y(\dpath/a_lt_b/_086_ ) );
sky130_fd_sc_hs__a21o_1 \dpath/a_lt_b/_145_ ( .A1(\dpath/a_lt_b/_061_ ), .A2(\dpath/a_lt_b/_062_ ), .B1(\dpath/a_lt_b/_060_ ), .X(\dpath/a_lt_b/_087_ ) );
sky130_fd_sc_hs__nand3_1 \dpath/a_lt_b/_146_ ( .A(\dpath/a_lt_b/_064_ ), .B(\dpath/a_lt_b/_058_ ), .C(\dpath/a_lt_b/_065_ ), .Y(\dpath/a_lt_b/_088_ ) );
sky130_fd_sc_hs__and4_1 \dpath/a_lt_b/_147_ ( .A(\dpath/a_lt_b/_080_ ), .B(\dpath/a_lt_b/_086_ ), .C(\dpath/a_lt_b/_087_ ), .D(\dpath/a_lt_b/_088_ ), .X(\dpath/a_lt_b/_089_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_148_ ( .A(\dpath/a_lt_b$in0[8] ), .X(\dpath/a_lt_b/_014_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_149_ ( .A(\dpath/a_lt_b$in1[8] ), .X(\dpath/a_lt_b/_030_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_150_ ( .A(\dpath/a_lt_b$in1[7] ), .X(\dpath/a_lt_b/_029_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_151_ ( .A(\dpath/a_lt_b$in0[7] ), .X(\dpath/a_lt_b/_013_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_152_ ( .A(\dpath/a_lt_b$in1[6] ), .X(\dpath/a_lt_b/_028_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_153_ ( .A(\dpath/a_lt_b$in0[6] ), .X(\dpath/a_lt_b/_012_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_154_ ( .A(\dpath/a_lt_b$in1[5] ), .X(\dpath/a_lt_b/_027_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_155_ ( .A(\dpath/a_lt_b$in0[5] ), .X(\dpath/a_lt_b/_011_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_156_ ( .A(\dpath/a_lt_b$in0[4] ), .X(\dpath/a_lt_b/_010_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_157_ ( .A(\dpath/a_lt_b$in1[4] ), .X(\dpath/a_lt_b/_026_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_158_ ( .A(\dpath/a_lt_b$in1[3] ), .X(\dpath/a_lt_b/_025_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_159_ ( .A(\dpath/a_lt_b$in0[3] ), .X(\dpath/a_lt_b/_009_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_160_ ( .A(\dpath/a_lt_b$in1[2] ), .X(\dpath/a_lt_b/_024_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_161_ ( .A(\dpath/a_lt_b$in0[2] ), .X(\dpath/a_lt_b/_008_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_162_ ( .A(\dpath/a_lt_b$in1[1] ), .X(\dpath/a_lt_b/_023_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_163_ ( .A(\dpath/a_lt_b$in0[1] ), .X(\dpath/a_lt_b/_007_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_164_ ( .A(\dpath/a_lt_b$in1[0] ), .X(\dpath/a_lt_b/_016_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_165_ ( .A(\dpath/a_lt_b$in0[0] ), .X(\dpath/a_lt_b/_000_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_166_ ( .A(\dpath/a_lt_b/_089_ ), .X(ctrl$is_a_lt_b ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_167_ ( .A(\dpath/a_lt_b$in1[15] ), .X(\dpath/a_lt_b/_022_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_168_ ( .A(\dpath/a_lt_b$in0[15] ), .X(\dpath/a_lt_b/_006_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_169_ ( .A(\dpath/a_lt_b$in1[14] ), .X(\dpath/a_lt_b/_021_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_170_ ( .A(\dpath/a_lt_b$in0[14] ), .X(\dpath/a_lt_b/_005_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_171_ ( .A(\dpath/a_lt_b$in1[13] ), .X(\dpath/a_lt_b/_020_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_172_ ( .A(\dpath/a_lt_b$in0[13] ), .X(\dpath/a_lt_b/_004_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_173_ ( .A(\dpath/a_lt_b$in0[12] ), .X(\dpath/a_lt_b/_003_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_174_ ( .A(\dpath/a_lt_b$in1[12] ), .X(\dpath/a_lt_b/_019_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_175_ ( .A(\dpath/a_lt_b$in1[11] ), .X(\dpath/a_lt_b/_018_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_176_ ( .A(\dpath/a_lt_b$in0[11] ), .X(\dpath/a_lt_b/_002_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_177_ ( .A(\dpath/a_lt_b$in1[10] ), .X(\dpath/a_lt_b/_017_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_178_ ( .A(\dpath/a_lt_b$in0[10] ), .X(\dpath/a_lt_b/_001_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_179_ ( .A(\dpath/a_lt_b$in1[9] ), .X(\dpath/a_lt_b/_031_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_lt_b/_180_ ( .A(\dpath/a_lt_b$in0[9] ), .X(\dpath/a_lt_b/_015_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_104_ ( .A(\dpath/a_mux/_000_ ), .Y(\dpath/a_mux/_062_ ) );
sky130_fd_sc_hs__xor2_4 \dpath/a_mux/_105_ ( .A(\dpath/a_mux/_102_ ), .B(\dpath/a_mux/_103_ ), .X(\dpath/a_mux/_063_ ) );
sky130_fd_sc_hs__buf_4 \dpath/a_mux/_106_ ( .A(\dpath/a_mux/_063_ ), .X(\dpath/a_mux/_064_ ) );
sky130_fd_sc_hs__and2b_4 \dpath/a_mux/_107_ ( .A_N(\dpath/a_mux/_103_ ), .B(\dpath/a_mux/_102_ ), .X(\dpath/a_mux/_065_ ) );
sky130_fd_sc_hs__buf_16 \dpath/a_mux/_108_ ( .A(\dpath/a_mux/_065_ ), .X(\dpath/a_mux/_066_ ) );
sky130_fd_sc_hs__and2b_4 \dpath/a_mux/_109_ ( .A_N(\dpath/a_mux/_102_ ), .B(\dpath/a_mux/_103_ ), .X(\dpath/a_mux/_067_ ) );
sky130_fd_sc_hs__buf_8 \dpath/a_mux/_110_ ( .A(\dpath/a_mux/_067_ ), .X(\dpath/a_mux/_068_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_111_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_016_ ), .B1(\dpath/a_mux/_032_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_069_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_112_ ( .A1(\dpath/a_mux/_062_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_069_ ), .Y(\dpath/a_mux/_086_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_113_ ( .A(\dpath/a_mux/_007_ ), .Y(\dpath/a_mux/_070_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_114_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_023_ ), .B1(\dpath/a_mux/_039_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_071_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_115_ ( .A1(\dpath/a_mux/_070_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_071_ ), .Y(\dpath/a_mux/_093_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_116_ ( .A(\dpath/a_mux/_008_ ), .Y(\dpath/a_mux/_072_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_117_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_024_ ), .B1(\dpath/a_mux/_040_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_073_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_118_ ( .A1(\dpath/a_mux/_072_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_073_ ), .Y(\dpath/a_mux/_094_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_119_ ( .A(\dpath/a_mux/_009_ ), .Y(\dpath/a_mux/_074_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_120_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_025_ ), .B1(\dpath/a_mux/_041_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_075_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_121_ ( .A1(\dpath/a_mux/_074_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_075_ ), .Y(\dpath/a_mux/_095_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_122_ ( .A(\dpath/a_mux/_010_ ), .Y(\dpath/a_mux/_076_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_123_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_026_ ), .B1(\dpath/a_mux/_042_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_077_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_124_ ( .A1(\dpath/a_mux/_076_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_077_ ), .Y(\dpath/a_mux/_096_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_125_ ( .A(\dpath/a_mux/_011_ ), .Y(\dpath/a_mux/_078_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_126_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_027_ ), .B1(\dpath/a_mux/_043_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_079_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_127_ ( .A1(\dpath/a_mux/_078_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_079_ ), .Y(\dpath/a_mux/_097_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_128_ ( .A(\dpath/a_mux/_012_ ), .Y(\dpath/a_mux/_080_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_129_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_028_ ), .B1(\dpath/a_mux/_044_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_081_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_130_ ( .A1(\dpath/a_mux/_080_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_081_ ), .Y(\dpath/a_mux/_098_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_131_ ( .A(\dpath/a_mux/_013_ ), .Y(\dpath/a_mux/_082_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_132_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_029_ ), .B1(\dpath/a_mux/_045_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_083_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_133_ ( .A1(\dpath/a_mux/_082_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_083_ ), .Y(\dpath/a_mux/_099_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_134_ ( .A(\dpath/a_mux/_014_ ), .Y(\dpath/a_mux/_084_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_135_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_030_ ), .B1(\dpath/a_mux/_046_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_085_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_136_ ( .A1(\dpath/a_mux/_084_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_085_ ), .Y(\dpath/a_mux/_100_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_137_ ( .A(\dpath/a_mux/_015_ ), .Y(\dpath/a_mux/_048_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_138_ ( .A1(\dpath/a_mux/_066_ ), .A2(\dpath/a_mux/_031_ ), .B1(\dpath/a_mux/_047_ ), .B2(\dpath/a_mux/_068_ ), .Y(\dpath/a_mux/_049_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_139_ ( .A1(\dpath/a_mux/_048_ ), .A2(\dpath/a_mux/_064_ ), .B1(\dpath/a_mux/_049_ ), .Y(\dpath/a_mux/_101_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_140_ ( .A(\dpath/a_mux/_001_ ), .Y(\dpath/a_mux/_050_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_141_ ( .A1(\dpath/a_mux/_065_ ), .A2(\dpath/a_mux/_017_ ), .B1(\dpath/a_mux/_033_ ), .B2(\dpath/a_mux/_067_ ), .Y(\dpath/a_mux/_051_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_142_ ( .A1(\dpath/a_mux/_050_ ), .A2(\dpath/a_mux/_063_ ), .B1(\dpath/a_mux/_051_ ), .Y(\dpath/a_mux/_087_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_143_ ( .A(\dpath/a_mux/_002_ ), .Y(\dpath/a_mux/_052_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_144_ ( .A1(\dpath/a_mux/_065_ ), .A2(\dpath/a_mux/_018_ ), .B1(\dpath/a_mux/_034_ ), .B2(\dpath/a_mux/_067_ ), .Y(\dpath/a_mux/_053_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_145_ ( .A1(\dpath/a_mux/_052_ ), .A2(\dpath/a_mux/_063_ ), .B1(\dpath/a_mux/_053_ ), .Y(\dpath/a_mux/_088_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_146_ ( .A(\dpath/a_mux/_003_ ), .Y(\dpath/a_mux/_054_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_147_ ( .A1(\dpath/a_mux/_065_ ), .A2(\dpath/a_mux/_019_ ), .B1(\dpath/a_mux/_035_ ), .B2(\dpath/a_mux/_067_ ), .Y(\dpath/a_mux/_055_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_148_ ( .A1(\dpath/a_mux/_054_ ), .A2(\dpath/a_mux/_063_ ), .B1(\dpath/a_mux/_055_ ), .Y(\dpath/a_mux/_089_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_149_ ( .A(\dpath/a_mux/_004_ ), .Y(\dpath/a_mux/_056_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_150_ ( .A1(\dpath/a_mux/_065_ ), .A2(\dpath/a_mux/_020_ ), .B1(\dpath/a_mux/_036_ ), .B2(\dpath/a_mux/_067_ ), .Y(\dpath/a_mux/_057_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_151_ ( .A1(\dpath/a_mux/_056_ ), .A2(\dpath/a_mux/_063_ ), .B1(\dpath/a_mux/_057_ ), .Y(\dpath/a_mux/_090_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_152_ ( .A(\dpath/a_mux/_005_ ), .Y(\dpath/a_mux/_058_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_153_ ( .A1(\dpath/a_mux/_065_ ), .A2(\dpath/a_mux/_021_ ), .B1(\dpath/a_mux/_037_ ), .B2(\dpath/a_mux/_067_ ), .Y(\dpath/a_mux/_059_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_154_ ( .A1(\dpath/a_mux/_058_ ), .A2(\dpath/a_mux/_063_ ), .B1(\dpath/a_mux/_059_ ), .Y(\dpath/a_mux/_091_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/a_mux/_155_ ( .A(\dpath/a_mux/_006_ ), .Y(\dpath/a_mux/_060_ ) );
sky130_fd_sc_hs__a22oi_1 \dpath/a_mux/_156_ ( .A1(\dpath/a_mux/_065_ ), .A2(\dpath/a_mux/_022_ ), .B1(\dpath/a_mux/_038_ ), .B2(\dpath/a_mux/_067_ ), .Y(\dpath/a_mux/_061_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/a_mux/_157_ ( .A1(\dpath/a_mux/_060_ ), .A2(\dpath/a_mux/_063_ ), .B1(\dpath/a_mux/_061_ ), .Y(\dpath/a_mux/_092_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_158_ ( .A(\ctrl$a_mux_sel[0] ), .X(\dpath/a_mux/_102_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_159_ ( .A(\ctrl$a_mux_sel[1] ), .X(\dpath/a_mux/_103_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_160_ ( .A(\dpath/a_lt_b$in1[0] ), .X(\dpath/a_mux/_032_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_161_ ( .A(\resp_msg[0] ), .X(\dpath/a_mux/_016_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_162_ ( .A(\req_msg[16] ), .X(\dpath/a_mux/_000_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_163_ ( .A(\dpath/a_mux/_086_ ), .X(\dpath/a_mux$out[0] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_164_ ( .A(\dpath/a_lt_b$in1[1] ), .X(\dpath/a_mux/_039_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_165_ ( .A(\resp_msg[1] ), .X(\dpath/a_mux/_023_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_166_ ( .A(\req_msg[17] ), .X(\dpath/a_mux/_007_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_167_ ( .A(\dpath/a_mux/_093_ ), .X(\dpath/a_mux$out[1] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_168_ ( .A(\dpath/a_lt_b$in1[2] ), .X(\dpath/a_mux/_040_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_169_ ( .A(\resp_msg[2] ), .X(\dpath/a_mux/_024_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_170_ ( .A(\req_msg[18] ), .X(\dpath/a_mux/_008_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_171_ ( .A(\dpath/a_mux/_094_ ), .X(\dpath/a_mux$out[2] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_172_ ( .A(\dpath/a_lt_b$in1[3] ), .X(\dpath/a_mux/_041_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_173_ ( .A(\resp_msg[3] ), .X(\dpath/a_mux/_025_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_174_ ( .A(\req_msg[19] ), .X(\dpath/a_mux/_009_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_175_ ( .A(\dpath/a_mux/_095_ ), .X(\dpath/a_mux$out[3] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_176_ ( .A(\dpath/a_lt_b$in1[4] ), .X(\dpath/a_mux/_042_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_177_ ( .A(\resp_msg[4] ), .X(\dpath/a_mux/_026_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_178_ ( .A(\req_msg[20] ), .X(\dpath/a_mux/_010_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_179_ ( .A(\dpath/a_mux/_096_ ), .X(\dpath/a_mux$out[4] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_180_ ( .A(\dpath/a_lt_b$in1[5] ), .X(\dpath/a_mux/_043_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_181_ ( .A(\resp_msg[5] ), .X(\dpath/a_mux/_027_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_182_ ( .A(\req_msg[21] ), .X(\dpath/a_mux/_011_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_183_ ( .A(\dpath/a_mux/_097_ ), .X(\dpath/a_mux$out[5] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_184_ ( .A(\dpath/a_lt_b$in1[6] ), .X(\dpath/a_mux/_044_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_185_ ( .A(\resp_msg[6] ), .X(\dpath/a_mux/_028_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_186_ ( .A(\req_msg[22] ), .X(\dpath/a_mux/_012_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_187_ ( .A(\dpath/a_mux/_098_ ), .X(\dpath/a_mux$out[6] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_188_ ( .A(\dpath/a_lt_b$in1[7] ), .X(\dpath/a_mux/_045_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_189_ ( .A(\resp_msg[7] ), .X(\dpath/a_mux/_029_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_190_ ( .A(\req_msg[23] ), .X(\dpath/a_mux/_013_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_191_ ( .A(\dpath/a_mux/_099_ ), .X(\dpath/a_mux$out[7] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_192_ ( .A(\dpath/a_lt_b$in1[8] ), .X(\dpath/a_mux/_046_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_193_ ( .A(\resp_msg[8] ), .X(\dpath/a_mux/_030_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_194_ ( .A(\req_msg[24] ), .X(\dpath/a_mux/_014_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_195_ ( .A(\dpath/a_mux/_100_ ), .X(\dpath/a_mux$out[8] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_196_ ( .A(\dpath/a_lt_b$in1[9] ), .X(\dpath/a_mux/_047_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_197_ ( .A(\resp_msg[9] ), .X(\dpath/a_mux/_031_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_198_ ( .A(\req_msg[25] ), .X(\dpath/a_mux/_015_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_199_ ( .A(\dpath/a_mux/_101_ ), .X(\dpath/a_mux$out[9] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_200_ ( .A(\dpath/a_lt_b$in1[10] ), .X(\dpath/a_mux/_033_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_201_ ( .A(\resp_msg[10] ), .X(\dpath/a_mux/_017_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_202_ ( .A(\req_msg[26] ), .X(\dpath/a_mux/_001_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_203_ ( .A(\dpath/a_mux/_087_ ), .X(\dpath/a_mux$out[10] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_204_ ( .A(\dpath/a_lt_b$in1[11] ), .X(\dpath/a_mux/_034_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_205_ ( .A(\resp_msg[11] ), .X(\dpath/a_mux/_018_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_206_ ( .A(\req_msg[27] ), .X(\dpath/a_mux/_002_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_207_ ( .A(\dpath/a_mux/_088_ ), .X(\dpath/a_mux$out[11] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_208_ ( .A(\dpath/a_lt_b$in1[12] ), .X(\dpath/a_mux/_035_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_209_ ( .A(\resp_msg[12] ), .X(\dpath/a_mux/_019_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_210_ ( .A(\req_msg[28] ), .X(\dpath/a_mux/_003_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_211_ ( .A(\dpath/a_mux/_089_ ), .X(\dpath/a_mux$out[12] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_212_ ( .A(\dpath/a_lt_b$in1[13] ), .X(\dpath/a_mux/_036_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_213_ ( .A(\resp_msg[13] ), .X(\dpath/a_mux/_020_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_214_ ( .A(\req_msg[29] ), .X(\dpath/a_mux/_004_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_215_ ( .A(\dpath/a_mux/_090_ ), .X(\dpath/a_mux$out[13] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_216_ ( .A(\dpath/a_lt_b$in1[14] ), .X(\dpath/a_mux/_037_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_217_ ( .A(\resp_msg[14] ), .X(\dpath/a_mux/_021_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_218_ ( .A(\req_msg[30] ), .X(\dpath/a_mux/_005_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_219_ ( .A(\dpath/a_mux/_091_ ), .X(\dpath/a_mux$out[14] ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_220_ ( .A(\dpath/a_lt_b$in1[15] ), .X(\dpath/a_mux/_038_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_221_ ( .A(\resp_msg[15] ), .X(\dpath/a_mux/_022_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_222_ ( .A(\req_msg[31] ), .X(\dpath/a_mux/_006_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_mux/_223_ ( .A(\dpath/a_mux/_092_ ), .X(\dpath/a_mux$out[15] ) );
sky130_fd_sc_hs__buf_16 \dpath/a_reg/_066_ ( .A(\dpath/a_reg/_032_ ), .X(\dpath/a_reg/_049_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_067_ ( .A0(\dpath/a_reg/_050_ ), .A1(\dpath/a_reg/_033_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_016_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_068_ ( .A0(\dpath/a_reg/_057_ ), .A1(\dpath/a_reg/_040_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_023_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_069_ ( .A0(\dpath/a_reg/_058_ ), .A1(\dpath/a_reg/_041_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_024_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_070_ ( .A0(\dpath/a_reg/_059_ ), .A1(\dpath/a_reg/_042_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_025_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_071_ ( .A0(\dpath/a_reg/_060_ ), .A1(\dpath/a_reg/_043_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_026_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_072_ ( .A0(\dpath/a_reg/_061_ ), .A1(\dpath/a_reg/_044_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_027_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_073_ ( .A0(\dpath/a_reg/_062_ ), .A1(\dpath/a_reg/_045_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_028_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_074_ ( .A0(\dpath/a_reg/_063_ ), .A1(\dpath/a_reg/_046_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_029_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_075_ ( .A0(\dpath/a_reg/_064_ ), .A1(\dpath/a_reg/_047_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_030_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_076_ ( .A0(\dpath/a_reg/_065_ ), .A1(\dpath/a_reg/_048_ ), .S(\dpath/a_reg/_049_ ), .X(\dpath/a_reg/_031_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_077_ ( .A0(\dpath/a_reg/_051_ ), .A1(\dpath/a_reg/_034_ ), .S(\dpath/a_reg/_032_ ), .X(\dpath/a_reg/_017_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_078_ ( .A0(\dpath/a_reg/_052_ ), .A1(\dpath/a_reg/_035_ ), .S(\dpath/a_reg/_032_ ), .X(\dpath/a_reg/_018_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_079_ ( .A0(\dpath/a_reg/_053_ ), .A1(\dpath/a_reg/_036_ ), .S(\dpath/a_reg/_032_ ), .X(\dpath/a_reg/_019_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_080_ ( .A0(\dpath/a_reg/_054_ ), .A1(\dpath/a_reg/_037_ ), .S(\dpath/a_reg/_032_ ), .X(\dpath/a_reg/_020_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_081_ ( .A0(\dpath/a_reg/_055_ ), .A1(\dpath/a_reg/_038_ ), .S(\dpath/a_reg/_032_ ), .X(\dpath/a_reg/_021_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/a_reg/_082_ ( .A0(\dpath/a_reg/_056_ ), .A1(\dpath/a_reg/_039_ ), .S(\dpath/a_reg/_032_ ), .X(\dpath/a_reg/_022_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_083_ ( .A(\dpath/a_lt_b$in0[0] ), .X(\dpath/a_reg/_050_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_084_ ( .A(\dpath/a_mux$out[0] ), .X(\dpath/a_reg/_033_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_085_ ( .A(ctrl$a_reg_en ), .X(\dpath/a_reg/_032_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_086_ ( .A(\dpath/a_reg/_016_ ), .X(\dpath/a_reg/_000_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_087_ ( .A(\dpath/a_lt_b$in0[1] ), .X(\dpath/a_reg/_057_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_088_ ( .A(\dpath/a_mux$out[1] ), .X(\dpath/a_reg/_040_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_089_ ( .A(\dpath/a_reg/_023_ ), .X(\dpath/a_reg/_007_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_090_ ( .A(\dpath/a_lt_b$in0[2] ), .X(\dpath/a_reg/_058_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_091_ ( .A(\dpath/a_mux$out[2] ), .X(\dpath/a_reg/_041_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_092_ ( .A(\dpath/a_reg/_024_ ), .X(\dpath/a_reg/_008_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_093_ ( .A(\dpath/a_lt_b$in0[3] ), .X(\dpath/a_reg/_059_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_094_ ( .A(\dpath/a_mux$out[3] ), .X(\dpath/a_reg/_042_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_095_ ( .A(\dpath/a_reg/_025_ ), .X(\dpath/a_reg/_009_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_096_ ( .A(\dpath/a_lt_b$in0[4] ), .X(\dpath/a_reg/_060_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_097_ ( .A(\dpath/a_mux$out[4] ), .X(\dpath/a_reg/_043_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_098_ ( .A(\dpath/a_reg/_026_ ), .X(\dpath/a_reg/_010_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_099_ ( .A(\dpath/a_lt_b$in0[5] ), .X(\dpath/a_reg/_061_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_100_ ( .A(\dpath/a_mux$out[5] ), .X(\dpath/a_reg/_044_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_101_ ( .A(\dpath/a_reg/_027_ ), .X(\dpath/a_reg/_011_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_102_ ( .A(\dpath/a_lt_b$in0[6] ), .X(\dpath/a_reg/_062_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_103_ ( .A(\dpath/a_mux$out[6] ), .X(\dpath/a_reg/_045_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_104_ ( .A(\dpath/a_reg/_028_ ), .X(\dpath/a_reg/_012_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_105_ ( .A(\dpath/a_lt_b$in0[7] ), .X(\dpath/a_reg/_063_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_106_ ( .A(\dpath/a_mux$out[7] ), .X(\dpath/a_reg/_046_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_107_ ( .A(\dpath/a_reg/_029_ ), .X(\dpath/a_reg/_013_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_108_ ( .A(\dpath/a_lt_b$in0[8] ), .X(\dpath/a_reg/_064_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_109_ ( .A(\dpath/a_mux$out[8] ), .X(\dpath/a_reg/_047_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_110_ ( .A(\dpath/a_reg/_030_ ), .X(\dpath/a_reg/_014_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_111_ ( .A(\dpath/a_lt_b$in0[9] ), .X(\dpath/a_reg/_065_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_112_ ( .A(\dpath/a_mux$out[9] ), .X(\dpath/a_reg/_048_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_113_ ( .A(\dpath/a_reg/_031_ ), .X(\dpath/a_reg/_015_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_114_ ( .A(\dpath/a_lt_b$in0[10] ), .X(\dpath/a_reg/_051_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_115_ ( .A(\dpath/a_mux$out[10] ), .X(\dpath/a_reg/_034_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_116_ ( .A(\dpath/a_reg/_017_ ), .X(\dpath/a_reg/_001_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_117_ ( .A(\dpath/a_lt_b$in0[11] ), .X(\dpath/a_reg/_052_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_118_ ( .A(\dpath/a_mux$out[11] ), .X(\dpath/a_reg/_035_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_119_ ( .A(\dpath/a_reg/_018_ ), .X(\dpath/a_reg/_002_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_120_ ( .A(\dpath/a_lt_b$in0[12] ), .X(\dpath/a_reg/_053_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_121_ ( .A(\dpath/a_mux$out[12] ), .X(\dpath/a_reg/_036_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_122_ ( .A(\dpath/a_reg/_019_ ), .X(\dpath/a_reg/_003_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_123_ ( .A(\dpath/a_lt_b$in0[13] ), .X(\dpath/a_reg/_054_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_124_ ( .A(\dpath/a_mux$out[13] ), .X(\dpath/a_reg/_037_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_125_ ( .A(\dpath/a_reg/_020_ ), .X(\dpath/a_reg/_004_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_126_ ( .A(\dpath/a_lt_b$in0[14] ), .X(\dpath/a_reg/_055_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_127_ ( .A(\dpath/a_mux$out[14] ), .X(\dpath/a_reg/_038_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_128_ ( .A(\dpath/a_reg/_021_ ), .X(\dpath/a_reg/_005_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_129_ ( .A(\dpath/a_lt_b$in0[15] ), .X(\dpath/a_reg/_056_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_130_ ( .A(\dpath/a_mux$out[15] ), .X(\dpath/a_reg/_039_ ) );
sky130_fd_sc_hs__buf_1 \dpath/a_reg/_131_ ( .A(\dpath/a_reg/_022_ ), .X(\dpath/a_reg/_006_ ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_132_ ( .D(\dpath/a_reg/_000_ ), .Q(\dpath/a_lt_b$in0[0] ), .CLK(clk_66 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_133_ ( .D(\dpath/a_reg/_007_ ), .Q(\dpath/a_lt_b$in0[1] ), .CLK(clk_64 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_134_ ( .D(\dpath/a_reg/_008_ ), .Q(\dpath/a_lt_b$in0[2] ), .CLK(clk_63 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_135_ ( .D(\dpath/a_reg/_009_ ), .Q(\dpath/a_lt_b$in0[3] ), .CLK(clk_63 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_136_ ( .D(\dpath/a_reg/_010_ ), .Q(\dpath/a_lt_b$in0[4] ), .CLK(clk_86 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_137_ ( .D(\dpath/a_reg/_011_ ), .Q(\dpath/a_lt_b$in0[5] ), .CLK(clk_86 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_138_ ( .D(\dpath/a_reg/_012_ ), .Q(\dpath/a_lt_b$in0[6] ), .CLK(clk_70 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_139_ ( .D(\dpath/a_reg/_013_ ), .Q(\dpath/a_lt_b$in0[7] ), .CLK(clk_68 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_140_ ( .D(\dpath/a_reg/_014_ ), .Q(\dpath/a_lt_b$in0[8] ), .CLK(clk_69 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_141_ ( .D(\dpath/a_reg/_015_ ), .Q(\dpath/a_lt_b$in0[9] ), .CLK(clk_74 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_142_ ( .D(\dpath/a_reg/_001_ ), .Q(\dpath/a_lt_b$in0[10] ), .CLK(clk_76 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_143_ ( .D(\dpath/a_reg/_002_ ), .Q(\dpath/a_lt_b$in0[11] ), .CLK(clk_78 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_144_ ( .D(\dpath/a_reg/_003_ ), .Q(\dpath/a_lt_b$in0[12] ), .CLK(clk_80 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_145_ ( .D(\dpath/a_reg/_004_ ), .Q(\dpath/a_lt_b$in0[13] ), .CLK(clk_79 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_146_ ( .D(\dpath/a_reg/_005_ ), .Q(\dpath/a_lt_b$in0[14] ), .CLK(clk_58 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/a_reg/_147_ ( .D(\dpath/a_reg/_006_ ), .Q(\dpath/a_lt_b$in0[15] ), .CLK(clk_82 ) );
sky130_fd_sc_hs__buf_16 \dpath/b_mux/_050_ ( .A(\dpath/b_mux/_049_ ), .X(\dpath/b_mux/_032_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_051_ ( .A0(\dpath/b_mux/_000_ ), .A1(\dpath/b_mux/_016_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_033_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_052_ ( .A0(\dpath/b_mux/_007_ ), .A1(\dpath/b_mux/_023_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_040_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_053_ ( .A0(\dpath/b_mux/_008_ ), .A1(\dpath/b_mux/_024_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_041_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_054_ ( .A0(\dpath/b_mux/_009_ ), .A1(\dpath/b_mux/_025_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_042_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_055_ ( .A0(\dpath/b_mux/_010_ ), .A1(\dpath/b_mux/_026_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_043_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_056_ ( .A0(\dpath/b_mux/_011_ ), .A1(\dpath/b_mux/_027_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_044_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_057_ ( .A0(\dpath/b_mux/_012_ ), .A1(\dpath/b_mux/_028_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_045_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_058_ ( .A0(\dpath/b_mux/_013_ ), .A1(\dpath/b_mux/_029_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_046_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_059_ ( .A0(\dpath/b_mux/_014_ ), .A1(\dpath/b_mux/_030_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_047_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_060_ ( .A0(\dpath/b_mux/_015_ ), .A1(\dpath/b_mux/_031_ ), .S(\dpath/b_mux/_032_ ), .X(\dpath/b_mux/_048_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_061_ ( .A0(\dpath/b_mux/_001_ ), .A1(\dpath/b_mux/_017_ ), .S(\dpath/b_mux/_049_ ), .X(\dpath/b_mux/_034_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_062_ ( .A0(\dpath/b_mux/_002_ ), .A1(\dpath/b_mux/_018_ ), .S(\dpath/b_mux/_049_ ), .X(\dpath/b_mux/_035_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_063_ ( .A0(\dpath/b_mux/_003_ ), .A1(\dpath/b_mux/_019_ ), .S(\dpath/b_mux/_049_ ), .X(\dpath/b_mux/_036_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_064_ ( .A0(\dpath/b_mux/_004_ ), .A1(\dpath/b_mux/_020_ ), .S(\dpath/b_mux/_049_ ), .X(\dpath/b_mux/_037_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_065_ ( .A0(\dpath/b_mux/_005_ ), .A1(\dpath/b_mux/_021_ ), .S(\dpath/b_mux/_049_ ), .X(\dpath/b_mux/_038_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_mux/_066_ ( .A0(\dpath/b_mux/_006_ ), .A1(\dpath/b_mux/_022_ ), .S(\dpath/b_mux/_049_ ), .X(\dpath/b_mux/_039_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_067_ ( .A(\dpath/a_lt_b$in0[0] ), .X(\dpath/b_mux/_000_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_068_ ( .A(\req_msg[0] ), .X(\dpath/b_mux/_016_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_069_ ( .A(ctrl$b_mux_sel ), .X(\dpath/b_mux/_049_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_070_ ( .A(\dpath/b_mux/_033_ ), .X(\dpath/b_mux$out[0] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_071_ ( .A(\dpath/a_lt_b$in0[1] ), .X(\dpath/b_mux/_007_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_072_ ( .A(\req_msg[1] ), .X(\dpath/b_mux/_023_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_073_ ( .A(\dpath/b_mux/_040_ ), .X(\dpath/b_mux$out[1] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_074_ ( .A(\dpath/a_lt_b$in0[2] ), .X(\dpath/b_mux/_008_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_075_ ( .A(\req_msg[2] ), .X(\dpath/b_mux/_024_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_076_ ( .A(\dpath/b_mux/_041_ ), .X(\dpath/b_mux$out[2] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_077_ ( .A(\dpath/a_lt_b$in0[3] ), .X(\dpath/b_mux/_009_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_078_ ( .A(\req_msg[3] ), .X(\dpath/b_mux/_025_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_079_ ( .A(\dpath/b_mux/_042_ ), .X(\dpath/b_mux$out[3] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_080_ ( .A(\dpath/a_lt_b$in0[4] ), .X(\dpath/b_mux/_010_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_081_ ( .A(\req_msg[4] ), .X(\dpath/b_mux/_026_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_082_ ( .A(\dpath/b_mux/_043_ ), .X(\dpath/b_mux$out[4] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_083_ ( .A(\dpath/a_lt_b$in0[5] ), .X(\dpath/b_mux/_011_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_084_ ( .A(\req_msg[5] ), .X(\dpath/b_mux/_027_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_085_ ( .A(\dpath/b_mux/_044_ ), .X(\dpath/b_mux$out[5] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_086_ ( .A(\dpath/a_lt_b$in0[6] ), .X(\dpath/b_mux/_012_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_087_ ( .A(\req_msg[6] ), .X(\dpath/b_mux/_028_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_088_ ( .A(\dpath/b_mux/_045_ ), .X(\dpath/b_mux$out[6] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_089_ ( .A(\dpath/a_lt_b$in0[7] ), .X(\dpath/b_mux/_013_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_090_ ( .A(\req_msg[7] ), .X(\dpath/b_mux/_029_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_091_ ( .A(\dpath/b_mux/_046_ ), .X(\dpath/b_mux$out[7] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_092_ ( .A(\dpath/a_lt_b$in0[8] ), .X(\dpath/b_mux/_014_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_093_ ( .A(\req_msg[8] ), .X(\dpath/b_mux/_030_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_094_ ( .A(\dpath/b_mux/_047_ ), .X(\dpath/b_mux$out[8] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_095_ ( .A(\dpath/a_lt_b$in0[9] ), .X(\dpath/b_mux/_015_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_096_ ( .A(\req_msg[9] ), .X(\dpath/b_mux/_031_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_097_ ( .A(\dpath/b_mux/_048_ ), .X(\dpath/b_mux$out[9] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_098_ ( .A(\dpath/a_lt_b$in0[10] ), .X(\dpath/b_mux/_001_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_099_ ( .A(\req_msg[10] ), .X(\dpath/b_mux/_017_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_100_ ( .A(\dpath/b_mux/_034_ ), .X(\dpath/b_mux$out[10] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_101_ ( .A(\dpath/a_lt_b$in0[11] ), .X(\dpath/b_mux/_002_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_102_ ( .A(\req_msg[11] ), .X(\dpath/b_mux/_018_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_103_ ( .A(\dpath/b_mux/_035_ ), .X(\dpath/b_mux$out[11] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_104_ ( .A(\dpath/a_lt_b$in0[12] ), .X(\dpath/b_mux/_003_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_105_ ( .A(\req_msg[12] ), .X(\dpath/b_mux/_019_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_106_ ( .A(\dpath/b_mux/_036_ ), .X(\dpath/b_mux$out[12] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_107_ ( .A(\dpath/a_lt_b$in0[13] ), .X(\dpath/b_mux/_004_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_108_ ( .A(\req_msg[13] ), .X(\dpath/b_mux/_020_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_109_ ( .A(\dpath/b_mux/_037_ ), .X(\dpath/b_mux$out[13] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_110_ ( .A(\dpath/a_lt_b$in0[14] ), .X(\dpath/b_mux/_005_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_111_ ( .A(\req_msg[14] ), .X(\dpath/b_mux/_021_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_112_ ( .A(\dpath/b_mux/_038_ ), .X(\dpath/b_mux$out[14] ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_113_ ( .A(\dpath/a_lt_b$in0[15] ), .X(\dpath/b_mux/_006_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_114_ ( .A(\req_msg[15] ), .X(\dpath/b_mux/_022_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_mux/_115_ ( .A(\dpath/b_mux/_039_ ), .X(\dpath/b_mux$out[15] ) );
sky130_fd_sc_hs__buf_16 \dpath/b_reg/_066_ ( .A(\dpath/b_reg/_032_ ), .X(\dpath/b_reg/_049_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_067_ ( .A0(\dpath/b_reg/_050_ ), .A1(\dpath/b_reg/_033_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_016_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_068_ ( .A0(\dpath/b_reg/_057_ ), .A1(\dpath/b_reg/_040_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_023_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_069_ ( .A0(\dpath/b_reg/_058_ ), .A1(\dpath/b_reg/_041_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_024_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_070_ ( .A0(\dpath/b_reg/_059_ ), .A1(\dpath/b_reg/_042_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_025_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_071_ ( .A0(\dpath/b_reg/_060_ ), .A1(\dpath/b_reg/_043_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_026_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_072_ ( .A0(\dpath/b_reg/_061_ ), .A1(\dpath/b_reg/_044_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_027_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_073_ ( .A0(\dpath/b_reg/_062_ ), .A1(\dpath/b_reg/_045_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_028_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_074_ ( .A0(\dpath/b_reg/_063_ ), .A1(\dpath/b_reg/_046_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_029_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_075_ ( .A0(\dpath/b_reg/_064_ ), .A1(\dpath/b_reg/_047_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_030_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_076_ ( .A0(\dpath/b_reg/_065_ ), .A1(\dpath/b_reg/_048_ ), .S(\dpath/b_reg/_049_ ), .X(\dpath/b_reg/_031_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_077_ ( .A0(\dpath/b_reg/_051_ ), .A1(\dpath/b_reg/_034_ ), .S(\dpath/b_reg/_032_ ), .X(\dpath/b_reg/_017_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_078_ ( .A0(\dpath/b_reg/_052_ ), .A1(\dpath/b_reg/_035_ ), .S(\dpath/b_reg/_032_ ), .X(\dpath/b_reg/_018_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_079_ ( .A0(\dpath/b_reg/_053_ ), .A1(\dpath/b_reg/_036_ ), .S(\dpath/b_reg/_032_ ), .X(\dpath/b_reg/_019_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_080_ ( .A0(\dpath/b_reg/_054_ ), .A1(\dpath/b_reg/_037_ ), .S(\dpath/b_reg/_032_ ), .X(\dpath/b_reg/_020_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_081_ ( .A0(\dpath/b_reg/_055_ ), .A1(\dpath/b_reg/_038_ ), .S(\dpath/b_reg/_032_ ), .X(\dpath/b_reg/_021_ ) );
sky130_fd_sc_hs__mux2_1 \dpath/b_reg/_082_ ( .A0(\dpath/b_reg/_056_ ), .A1(\dpath/b_reg/_039_ ), .S(\dpath/b_reg/_032_ ), .X(\dpath/b_reg/_022_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_083_ ( .A(\dpath/a_lt_b$in1[0] ), .X(\dpath/b_reg/_050_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_084_ ( .A(\dpath/b_mux$out[0] ), .X(\dpath/b_reg/_033_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_085_ ( .A(ctrl$b_reg_en ), .X(\dpath/b_reg/_032_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_086_ ( .A(\dpath/b_reg/_016_ ), .X(\dpath/b_reg/_000_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_087_ ( .A(\dpath/a_lt_b$in1[1] ), .X(\dpath/b_reg/_057_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_088_ ( .A(\dpath/b_mux$out[1] ), .X(\dpath/b_reg/_040_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_089_ ( .A(\dpath/b_reg/_023_ ), .X(\dpath/b_reg/_007_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_090_ ( .A(\dpath/a_lt_b$in1[2] ), .X(\dpath/b_reg/_058_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_091_ ( .A(\dpath/b_mux$out[2] ), .X(\dpath/b_reg/_041_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_092_ ( .A(\dpath/b_reg/_024_ ), .X(\dpath/b_reg/_008_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_093_ ( .A(\dpath/a_lt_b$in1[3] ), .X(\dpath/b_reg/_059_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_094_ ( .A(\dpath/b_mux$out[3] ), .X(\dpath/b_reg/_042_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_095_ ( .A(\dpath/b_reg/_025_ ), .X(\dpath/b_reg/_009_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_096_ ( .A(\dpath/a_lt_b$in1[4] ), .X(\dpath/b_reg/_060_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_097_ ( .A(\dpath/b_mux$out[4] ), .X(\dpath/b_reg/_043_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_098_ ( .A(\dpath/b_reg/_026_ ), .X(\dpath/b_reg/_010_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_099_ ( .A(\dpath/a_lt_b$in1[5] ), .X(\dpath/b_reg/_061_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_100_ ( .A(\dpath/b_mux$out[5] ), .X(\dpath/b_reg/_044_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_101_ ( .A(\dpath/b_reg/_027_ ), .X(\dpath/b_reg/_011_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_102_ ( .A(\dpath/a_lt_b$in1[6] ), .X(\dpath/b_reg/_062_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_103_ ( .A(\dpath/b_mux$out[6] ), .X(\dpath/b_reg/_045_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_104_ ( .A(\dpath/b_reg/_028_ ), .X(\dpath/b_reg/_012_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_105_ ( .A(\dpath/a_lt_b$in1[7] ), .X(\dpath/b_reg/_063_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_106_ ( .A(\dpath/b_mux$out[7] ), .X(\dpath/b_reg/_046_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_107_ ( .A(\dpath/b_reg/_029_ ), .X(\dpath/b_reg/_013_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_108_ ( .A(\dpath/a_lt_b$in1[8] ), .X(\dpath/b_reg/_064_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_109_ ( .A(\dpath/b_mux$out[8] ), .X(\dpath/b_reg/_047_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_110_ ( .A(\dpath/b_reg/_030_ ), .X(\dpath/b_reg/_014_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_111_ ( .A(\dpath/a_lt_b$in1[9] ), .X(\dpath/b_reg/_065_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_112_ ( .A(\dpath/b_mux$out[9] ), .X(\dpath/b_reg/_048_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_113_ ( .A(\dpath/b_reg/_031_ ), .X(\dpath/b_reg/_015_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_114_ ( .A(\dpath/a_lt_b$in1[10] ), .X(\dpath/b_reg/_051_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_115_ ( .A(\dpath/b_mux$out[10] ), .X(\dpath/b_reg/_034_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_116_ ( .A(\dpath/b_reg/_017_ ), .X(\dpath/b_reg/_001_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_117_ ( .A(\dpath/a_lt_b$in1[11] ), .X(\dpath/b_reg/_052_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_118_ ( .A(\dpath/b_mux$out[11] ), .X(\dpath/b_reg/_035_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_119_ ( .A(\dpath/b_reg/_018_ ), .X(\dpath/b_reg/_002_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_120_ ( .A(\dpath/a_lt_b$in1[12] ), .X(\dpath/b_reg/_053_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_121_ ( .A(\dpath/b_mux$out[12] ), .X(\dpath/b_reg/_036_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_122_ ( .A(\dpath/b_reg/_019_ ), .X(\dpath/b_reg/_003_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_123_ ( .A(\dpath/a_lt_b$in1[13] ), .X(\dpath/b_reg/_054_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_124_ ( .A(\dpath/b_mux$out[13] ), .X(\dpath/b_reg/_037_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_125_ ( .A(\dpath/b_reg/_020_ ), .X(\dpath/b_reg/_004_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_126_ ( .A(\dpath/a_lt_b$in1[14] ), .X(\dpath/b_reg/_055_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_127_ ( .A(\dpath/b_mux$out[14] ), .X(\dpath/b_reg/_038_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_128_ ( .A(\dpath/b_reg/_021_ ), .X(\dpath/b_reg/_005_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_129_ ( .A(\dpath/a_lt_b$in1[15] ), .X(\dpath/b_reg/_056_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_130_ ( .A(\dpath/b_mux$out[15] ), .X(\dpath/b_reg/_039_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_reg/_131_ ( .A(\dpath/b_reg/_022_ ), .X(\dpath/b_reg/_006_ ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_132_ ( .D(\dpath/b_reg/_000_ ), .Q(\dpath/a_lt_b$in1[0] ), .CLK(clk_67 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_133_ ( .D(\dpath/b_reg/_007_ ), .Q(\dpath/a_lt_b$in1[1] ), .CLK(clk_65 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_134_ ( .D(\dpath/b_reg/_008_ ), .Q(\dpath/a_lt_b$in1[2] ), .CLK(clk_62 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_135_ ( .D(\dpath/b_reg/_009_ ), .Q(\dpath/a_lt_b$in1[3] ), .CLK(clk_62 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_136_ ( .D(\dpath/b_reg/_010_ ), .Q(\dpath/a_lt_b$in1[4] ), .CLK(clk_72 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_137_ ( .D(\dpath/b_reg/_011_ ), .Q(\dpath/a_lt_b$in1[5] ), .CLK(clk_73 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_138_ ( .D(\dpath/b_reg/_012_ ), .Q(\dpath/a_lt_b$in1[6] ), .CLK(clk_75 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_139_ ( .D(\dpath/b_reg/_013_ ), .Q(\dpath/a_lt_b$in1[7] ), .CLK(clk_71 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_140_ ( .D(\dpath/b_reg/_014_ ), .Q(\dpath/a_lt_b$in1[8] ), .CLK(clk_77 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_141_ ( .D(\dpath/b_reg/_015_ ), .Q(\dpath/a_lt_b$in1[9] ), .CLK(clk_77 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_142_ ( .D(\dpath/b_reg/_001_ ), .Q(\dpath/a_lt_b$in1[10] ), .CLK(clk_76 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_143_ ( .D(\dpath/b_reg/_002_ ), .Q(\dpath/a_lt_b$in1[11] ), .CLK(clk_83 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_144_ ( .D(\dpath/b_reg/_003_ ), .Q(\dpath/a_lt_b$in1[12] ), .CLK(clk_84 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_145_ ( .D(\dpath/b_reg/_004_ ), .Q(\dpath/a_lt_b$in1[13] ), .CLK(clk_57 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_146_ ( .D(\dpath/b_reg/_005_ ), .Q(\dpath/a_lt_b$in1[14] ), .CLK(clk_81 ) );
sky130_fd_sc_hs__dfxtp_1 \dpath/b_reg/_147_ ( .D(\dpath/b_reg/_006_ ), .Q(\dpath/a_lt_b$in1[15] ), .CLK(clk_58 ) );
sky130_fd_sc_hs__nor2_2 \dpath/b_zero/_25_ ( .A(\dpath/b_zero/_10_ ), .B(\dpath/b_zero/_13_ ), .Y(\dpath/b_zero/_16_ ) );
sky130_fd_sc_hs__nor3b_1 \dpath/b_zero/_26_ ( .A(\dpath/b_zero/_07_ ), .B(\dpath/b_zero/_08_ ), .C_N(\dpath/b_zero/_16_ ), .Y(\dpath/b_zero/_17_ ) );
sky130_fd_sc_hs__nor2_4 \dpath/b_zero/_27_ ( .A(\dpath/b_zero/_04_ ), .B(\dpath/b_zero/_05_ ), .Y(\dpath/b_zero/_18_ ) );
sky130_fd_sc_hs__nor3b_1 \dpath/b_zero/_28_ ( .A(\dpath/b_zero/_14_ ), .B(\dpath/b_zero/_02_ ), .C_N(\dpath/b_zero/_18_ ), .Y(\dpath/b_zero/_19_ ) );
sky130_fd_sc_hs__nor2_1 \dpath/b_zero/_29_ ( .A(\dpath/b_zero/_00_ ), .B(\dpath/b_zero/_09_ ), .Y(\dpath/b_zero/_20_ ) );
sky130_fd_sc_hs__nor3b_2 \dpath/b_zero/_30_ ( .A(\dpath/b_zero/_11_ ), .B(\dpath/b_zero/_12_ ), .C_N(\dpath/b_zero/_20_ ), .Y(\dpath/b_zero/_21_ ) );
sky130_fd_sc_hs__nor2_1 \dpath/b_zero/_31_ ( .A(\dpath/b_zero/_03_ ), .B(\dpath/b_zero/_06_ ), .Y(\dpath/b_zero/_22_ ) );
sky130_fd_sc_hs__nor3b_2 \dpath/b_zero/_32_ ( .A(\dpath/b_zero/_15_ ), .B(\dpath/b_zero/_01_ ), .C_N(\dpath/b_zero/_22_ ), .Y(\dpath/b_zero/_23_ ) );
sky130_fd_sc_hs__and4_1 \dpath/b_zero/_33_ ( .A(\dpath/b_zero/_17_ ), .B(\dpath/b_zero/_19_ ), .C(\dpath/b_zero/_21_ ), .D(\dpath/b_zero/_23_ ), .X(\dpath/b_zero/_24_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_34_ ( .A(\dpath/a_lt_b$in1[1] ), .X(\dpath/b_zero/_07_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_35_ ( .A(\dpath/a_lt_b$in1[0] ), .X(\dpath/b_zero/_00_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_36_ ( .A(\dpath/a_lt_b$in1[3] ), .X(\dpath/b_zero/_09_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_37_ ( .A(\dpath/a_lt_b$in1[2] ), .X(\dpath/b_zero/_08_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_38_ ( .A(\dpath/a_lt_b$in1[5] ), .X(\dpath/b_zero/_11_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_39_ ( .A(\dpath/a_lt_b$in1[4] ), .X(\dpath/b_zero/_10_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_40_ ( .A(\dpath/a_lt_b$in1[7] ), .X(\dpath/b_zero/_13_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_41_ ( .A(\dpath/a_lt_b$in1[6] ), .X(\dpath/b_zero/_12_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_42_ ( .A(\dpath/a_lt_b$in1[9] ), .X(\dpath/b_zero/_15_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_43_ ( .A(\dpath/a_lt_b$in1[8] ), .X(\dpath/b_zero/_14_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_44_ ( .A(\dpath/a_lt_b$in1[11] ), .X(\dpath/b_zero/_02_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_45_ ( .A(\dpath/a_lt_b$in1[10] ), .X(\dpath/b_zero/_01_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_46_ ( .A(\dpath/a_lt_b$in1[13] ), .X(\dpath/b_zero/_04_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_47_ ( .A(\dpath/a_lt_b$in1[12] ), .X(\dpath/b_zero/_03_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_48_ ( .A(\dpath/a_lt_b$in1[15] ), .X(\dpath/b_zero/_06_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_49_ ( .A(\dpath/a_lt_b$in1[14] ), .X(\dpath/b_zero/_05_ ) );
sky130_fd_sc_hs__buf_1 \dpath/b_zero/_50_ ( .A(\dpath/b_zero/_24_ ), .X(ctrl$is_b_zero ) );
sky130_fd_sc_hs__xor2_1 \dpath/sub/_121_ ( .A(\dpath/sub/_000_ ), .B(\dpath/sub/_016_ ), .X(\dpath/sub/_105_ ) );
sky130_fd_sc_hs__nand2b_4 \dpath/sub/_122_ ( .A_N(\dpath/sub/_000_ ), .B(\dpath/sub/_016_ ), .Y(\dpath/sub/_063_ ) );
sky130_fd_sc_hs__xnor3_4 \dpath/sub/_123_ ( .A(\dpath/sub/_007_ ), .B(\dpath/sub/_023_ ), .C(\dpath/sub/_063_ ), .X(\dpath/sub/_112_ ) );
sky130_fd_sc_hs__nand2b_4 \dpath/sub/_124_ ( .A_N(\dpath/sub/_023_ ), .B(\dpath/sub/_007_ ), .Y(\dpath/sub/_064_ ) );
sky130_fd_sc_hs__nand2b_4 \dpath/sub/_125_ ( .A_N(\dpath/sub/_007_ ), .B(\dpath/sub/_023_ ), .Y(\dpath/sub/_065_ ) );
sky130_fd_sc_hs__nand3_2 \dpath/sub/_126_ ( .A(\dpath/sub/_063_ ), .B(\dpath/sub/_064_ ), .C(\dpath/sub/_065_ ), .Y(\dpath/sub/_066_ ) );
sky130_fd_sc_hs__nand2_2 \dpath/sub/_127_ ( .A(\dpath/sub/_066_ ), .B(\dpath/sub/_064_ ), .Y(\dpath/sub/_067_ ) );
sky130_fd_sc_hs__xnor3_4 \dpath/sub/_128_ ( .A(\dpath/sub/_008_ ), .B(\dpath/sub/_024_ ), .C(\dpath/sub/_067_ ), .X(\dpath/sub/_113_ ) );
sky130_fd_sc_hs__xnor2_4 \dpath/sub/_129_ ( .A(\dpath/sub/_009_ ), .B(\dpath/sub/_025_ ), .Y(\dpath/sub/_068_ ) );
sky130_fd_sc_hs__and2b_4 \dpath/sub/_130_ ( .A_N(\dpath/sub/_024_ ), .B(\dpath/sub/_008_ ), .X(\dpath/sub/_069_ ) );
sky130_fd_sc_hs__xnor2_4 \dpath/sub/_131_ ( .A(\dpath/sub/_008_ ), .B(\dpath/sub/_024_ ), .Y(\dpath/sub/_070_ ) );
sky130_fd_sc_hs__a21boi_1 \dpath/sub/_132_ ( .A1(\dpath/sub/_066_ ), .A2(\dpath/sub/_064_ ), .B1_N(\dpath/sub/_070_ ), .Y(\dpath/sub/_071_ ) );
sky130_fd_sc_hs__nor2_1 \dpath/sub/_133_ ( .A(\dpath/sub/_069_ ), .B(\dpath/sub/_071_ ), .Y(\dpath/sub/_072_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_134_ ( .A(\dpath/sub/_068_ ), .B(\dpath/sub/_072_ ), .Y(\dpath/sub/_114_ ) );
sky130_fd_sc_hs__nand3_4 \dpath/sub/_135_ ( .A(\dpath/sub/_067_ ), .B(\dpath/sub/_070_ ), .C(\dpath/sub/_068_ ), .Y(\dpath/sub/_073_ ) );
sky130_fd_sc_hs__nor2b_2 \dpath/sub/_136_ ( .A(\dpath/sub/_025_ ), .B_N(\dpath/sub/_009_ ), .Y(\dpath/sub/_074_ ) );
sky130_fd_sc_hs__a21oi_2 \dpath/sub/_137_ ( .A1(\dpath/sub/_068_ ), .A2(\dpath/sub/_069_ ), .B1(\dpath/sub/_074_ ), .Y(\dpath/sub/_075_ ) );
sky130_fd_sc_hs__xnor2_2 \dpath/sub/_138_ ( .A(\dpath/sub/_010_ ), .B(\dpath/sub/_026_ ), .Y(\dpath/sub/_076_ ) );
sky130_fd_sc_hs__a21bo_1 \dpath/sub/_139_ ( .A1(\dpath/sub/_073_ ), .A2(\dpath/sub/_075_ ), .B1_N(\dpath/sub/_076_ ), .X(\dpath/sub/_077_ ) );
sky130_fd_sc_hs__nand3b_1 \dpath/sub/_140_ ( .A_N(\dpath/sub/_076_ ), .B(\dpath/sub/_073_ ), .C(\dpath/sub/_075_ ), .Y(\dpath/sub/_078_ ) );
sky130_fd_sc_hs__and2_1 \dpath/sub/_141_ ( .A(\dpath/sub/_077_ ), .B(\dpath/sub/_078_ ), .X(\dpath/sub/_115_ ) );
sky130_fd_sc_hs__xnor2_4 \dpath/sub/_142_ ( .A(\dpath/sub/_011_ ), .B(\dpath/sub/_027_ ), .Y(\dpath/sub/_079_ ) );
sky130_fd_sc_hs__nor2b_4 \dpath/sub/_143_ ( .A(\dpath/sub/_026_ ), .B_N(\dpath/sub/_010_ ), .Y(\dpath/sub/_080_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_144_ ( .A_N(\dpath/sub/_080_ ), .B(\dpath/sub/_077_ ), .X(\dpath/sub/_081_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_145_ ( .A(\dpath/sub/_079_ ), .B(\dpath/sub/_081_ ), .Y(\dpath/sub/_116_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_146_ ( .A_N(\dpath/sub/_027_ ), .B(\dpath/sub/_011_ ), .X(\dpath/sub/_082_ ) );
sky130_fd_sc_hs__a21oi_2 \dpath/sub/_147_ ( .A1(\dpath/sub/_079_ ), .A2(\dpath/sub/_080_ ), .B1(\dpath/sub/_082_ ), .Y(\dpath/sub/_083_ ) );
sky130_fd_sc_hs__inv_2 \dpath/sub/_148_ ( .A(\dpath/sub/_083_ ), .Y(\dpath/sub/_084_ ) );
sky130_fd_sc_hs__xnor2_4 \dpath/sub/_149_ ( .A(\dpath/sub/_012_ ), .B(\dpath/sub/_028_ ), .Y(\dpath/sub/_085_ ) );
sky130_fd_sc_hs__and2_1 \dpath/sub/_150_ ( .A(\dpath/sub/_076_ ), .B(\dpath/sub/_079_ ), .X(\dpath/sub/_086_ ) );
sky130_fd_sc_hs__a21boi_1 \dpath/sub/_151_ ( .A1(\dpath/sub/_073_ ), .A2(\dpath/sub/_075_ ), .B1_N(\dpath/sub/_086_ ), .Y(\dpath/sub/_087_ ) );
sky130_fd_sc_hs__or3_1 \dpath/sub/_152_ ( .A(\dpath/sub/_084_ ), .B(\dpath/sub/_085_ ), .C(\dpath/sub/_087_ ), .X(\dpath/sub/_088_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/sub/_153_ ( .A1(\dpath/sub/_084_ ), .A2(\dpath/sub/_087_ ), .B1(\dpath/sub/_085_ ), .Y(\dpath/sub/_089_ ) );
sky130_fd_sc_hs__and2_1 \dpath/sub/_154_ ( .A(\dpath/sub/_088_ ), .B(\dpath/sub/_089_ ), .X(\dpath/sub/_117_ ) );
sky130_fd_sc_hs__xnor2_2 \dpath/sub/_155_ ( .A(\dpath/sub/_013_ ), .B(\dpath/sub/_029_ ), .Y(\dpath/sub/_090_ ) );
sky130_fd_sc_hs__inv_1 \dpath/sub/_156_ ( .A(\dpath/sub/_090_ ), .Y(\dpath/sub/_091_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/sub/_157_ ( .A(\dpath/sub/_028_ ), .B_N(\dpath/sub/_012_ ), .X(\dpath/sub/_092_ ) );
sky130_fd_sc_hs__nand2_1 \dpath/sub/_158_ ( .A(\dpath/sub/_089_ ), .B(\dpath/sub/_092_ ), .Y(\dpath/sub/_093_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_159_ ( .A(\dpath/sub/_091_ ), .B(\dpath/sub/_093_ ), .Y(\dpath/sub/_118_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_160_ ( .A(\dpath/sub/_014_ ), .B(\dpath/sub/_030_ ), .Y(\dpath/sub/_094_ ) );
sky130_fd_sc_hs__and4_1 \dpath/sub/_161_ ( .A(\dpath/sub/_076_ ), .B(\dpath/sub/_079_ ), .C(\dpath/sub/_085_ ), .D(\dpath/sub/_090_ ), .X(\dpath/sub/_095_ ) );
sky130_fd_sc_hs__a21boi_4 \dpath/sub/_162_ ( .A1(\dpath/sub/_073_ ), .A2(\dpath/sub/_075_ ), .B1_N(\dpath/sub/_095_ ), .Y(\dpath/sub/_096_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_163_ ( .A_N(\dpath/sub/_029_ ), .B(\dpath/sub/_013_ ), .X(\dpath/sub/_097_ ) );
sky130_fd_sc_hs__o21bai_1 \dpath/sub/_164_ ( .A1(\dpath/sub/_092_ ), .A2(\dpath/sub/_091_ ), .B1_N(\dpath/sub/_097_ ), .Y(\dpath/sub/_098_ ) );
sky130_fd_sc_hs__a31oi_1 \dpath/sub/_165_ ( .A1(\dpath/sub/_084_ ), .A2(\dpath/sub/_085_ ), .A3(\dpath/sub/_090_ ), .B1(\dpath/sub/_098_ ), .Y(\dpath/sub/_099_ ) );
sky130_fd_sc_hs__nor2b_2 \dpath/sub/_166_ ( .A(\dpath/sub/_096_ ), .B_N(\dpath/sub/_099_ ), .Y(\dpath/sub/_100_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_167_ ( .A(\dpath/sub/_094_ ), .B(\dpath/sub/_100_ ), .Y(\dpath/sub/_119_ ) );
sky130_fd_sc_hs__xnor2_4 \dpath/sub/_168_ ( .A(\dpath/sub/_015_ ), .B(\dpath/sub/_031_ ), .Y(\dpath/sub/_101_ ) );
sky130_fd_sc_hs__nor2b_4 \dpath/sub/_169_ ( .A(\dpath/sub/_030_ ), .B_N(\dpath/sub/_014_ ), .Y(\dpath/sub/_102_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/sub/_170_ ( .A(\dpath/sub/_100_ ), .B_N(\dpath/sub/_094_ ), .X(\dpath/sub/_103_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_171_ ( .A_N(\dpath/sub/_102_ ), .B(\dpath/sub/_103_ ), .X(\dpath/sub/_104_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_172_ ( .A(\dpath/sub/_101_ ), .B(\dpath/sub/_104_ ), .Y(\dpath/sub/_120_ ) );
sky130_fd_sc_hs__nand3b_1 \dpath/sub/_173_ ( .A_N(\dpath/sub/_100_ ), .B(\dpath/sub/_094_ ), .C(\dpath/sub/_101_ ), .Y(\dpath/sub/_032_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_174_ ( .A_N(\dpath/sub/_031_ ), .B(\dpath/sub/_015_ ), .X(\dpath/sub/_033_ ) );
sky130_fd_sc_hs__a21oi_4 \dpath/sub/_175_ ( .A1(\dpath/sub/_101_ ), .A2(\dpath/sub/_102_ ), .B1(\dpath/sub/_033_ ), .Y(\dpath/sub/_034_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_176_ ( .A(\dpath/sub/_001_ ), .B(\dpath/sub/_017_ ), .Y(\dpath/sub/_035_ ) );
sky130_fd_sc_hs__inv_1 \dpath/sub/_177_ ( .A(\dpath/sub/_035_ ), .Y(\dpath/sub/_036_ ) );
sky130_fd_sc_hs__a21o_1 \dpath/sub/_178_ ( .A1(\dpath/sub/_032_ ), .A2(\dpath/sub/_034_ ), .B1(\dpath/sub/_036_ ), .X(\dpath/sub/_037_ ) );
sky130_fd_sc_hs__nand3_1 \dpath/sub/_179_ ( .A(\dpath/sub/_032_ ), .B(\dpath/sub/_034_ ), .C(\dpath/sub/_036_ ), .Y(\dpath/sub/_038_ ) );
sky130_fd_sc_hs__and2_1 \dpath/sub/_180_ ( .A(\dpath/sub/_037_ ), .B(\dpath/sub/_038_ ), .X(\dpath/sub/_106_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_181_ ( .A(\dpath/sub/_002_ ), .B(\dpath/sub/_018_ ), .Y(\dpath/sub/_039_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_182_ ( .A_N(\dpath/sub/_017_ ), .B(\dpath/sub/_001_ ), .X(\dpath/sub/_040_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_183_ ( .A_N(\dpath/sub/_040_ ), .B(\dpath/sub/_037_ ), .X(\dpath/sub/_041_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_184_ ( .A(\dpath/sub/_039_ ), .B(\dpath/sub/_041_ ), .Y(\dpath/sub/_107_ ) );
sky130_fd_sc_hs__and4_1 \dpath/sub/_185_ ( .A(\dpath/sub/_094_ ), .B(\dpath/sub/_101_ ), .C(\dpath/sub/_035_ ), .D(\dpath/sub/_039_ ), .X(\dpath/sub/_042_ ) );
sky130_fd_sc_hs__nand2b_2 \dpath/sub/_186_ ( .A_N(\dpath/sub/_100_ ), .B(\dpath/sub/_042_ ), .Y(\dpath/sub/_043_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_187_ ( .A_N(\dpath/sub/_018_ ), .B(\dpath/sub/_002_ ), .X(\dpath/sub/_044_ ) );
sky130_fd_sc_hs__nor3b_1 \dpath/sub/_188_ ( .A(\dpath/sub/_036_ ), .B(\dpath/sub/_034_ ), .C_N(\dpath/sub/_039_ ), .Y(\dpath/sub/_045_ ) );
sky130_fd_sc_hs__a211oi_1 \dpath/sub/_189_ ( .A1(\dpath/sub/_040_ ), .A2(\dpath/sub/_039_ ), .B1(\dpath/sub/_044_ ), .C1(\dpath/sub/_045_ ), .Y(\dpath/sub/_046_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_190_ ( .A(\dpath/sub/_003_ ), .B(\dpath/sub/_019_ ), .Y(\dpath/sub/_047_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/sub/_191_ ( .A(\dpath/sub/_047_ ), .Y(\dpath/sub/_048_ ) );
sky130_fd_sc_hs__a21o_1 \dpath/sub/_192_ ( .A1(\dpath/sub/_043_ ), .A2(\dpath/sub/_046_ ), .B1(\dpath/sub/_048_ ), .X(\dpath/sub/_049_ ) );
sky130_fd_sc_hs__nand3_1 \dpath/sub/_193_ ( .A(\dpath/sub/_043_ ), .B(\dpath/sub/_046_ ), .C(\dpath/sub/_048_ ), .Y(\dpath/sub/_050_ ) );
sky130_fd_sc_hs__and2_1 \dpath/sub/_194_ ( .A(\dpath/sub/_049_ ), .B(\dpath/sub/_050_ ), .X(\dpath/sub/_108_ ) );
sky130_fd_sc_hs__xor2_1 \dpath/sub/_195_ ( .A(\dpath/sub/_004_ ), .B(\dpath/sub/_020_ ), .X(\dpath/sub/_051_ ) );
sky130_fd_sc_hs__and2b_1 \dpath/sub/_196_ ( .A_N(\dpath/sub/_019_ ), .B(\dpath/sub/_003_ ), .X(\dpath/sub/_052_ ) );
sky130_fd_sc_hs__bufinv_8 \dpath/sub/_197_ ( .A(\dpath/sub/_052_ ), .Y(\dpath/sub/_053_ ) );
sky130_fd_sc_hs__nand2_1 \dpath/sub/_198_ ( .A(\dpath/sub/_049_ ), .B(\dpath/sub/_053_ ), .Y(\dpath/sub/_054_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_199_ ( .A(\dpath/sub/_051_ ), .B(\dpath/sub/_054_ ), .Y(\dpath/sub/_109_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/sub/_200_ ( .A(\dpath/sub/_020_ ), .B_N(\dpath/sub/_004_ ), .X(\dpath/sub/_055_ ) );
sky130_fd_sc_hs__o21ai_1 \dpath/sub/_201_ ( .A1(\dpath/sub/_053_ ), .A2(\dpath/sub/_051_ ), .B1(\dpath/sub/_055_ ), .Y(\dpath/sub/_056_ ) );
sky130_fd_sc_hs__xnor2_1 \dpath/sub/_202_ ( .A(\dpath/sub/_005_ ), .B(\dpath/sub/_021_ ), .Y(\dpath/sub/_057_ ) );
sky130_fd_sc_hs__a211oi_2 \dpath/sub/_203_ ( .A1(\dpath/sub/_043_ ), .A2(\dpath/sub/_046_ ), .B1(\dpath/sub/_048_ ), .C1(\dpath/sub/_051_ ), .Y(\dpath/sub/_058_ ) );
sky130_fd_sc_hs__or3_1 \dpath/sub/_204_ ( .A(\dpath/sub/_056_ ), .B(\dpath/sub/_057_ ), .C(\dpath/sub/_058_ ), .X(\dpath/sub/_059_ ) );
sky130_fd_sc_hs__o21ai_2 \dpath/sub/_205_ ( .A1(\dpath/sub/_056_ ), .A2(\dpath/sub/_058_ ), .B1(\dpath/sub/_057_ ), .Y(\dpath/sub/_060_ ) );
sky130_fd_sc_hs__and2_1 \dpath/sub/_206_ ( .A(\dpath/sub/_059_ ), .B(\dpath/sub/_060_ ), .X(\dpath/sub/_110_ ) );
sky130_fd_sc_hs__or2b_1 \dpath/sub/_207_ ( .A(\dpath/sub/_021_ ), .B_N(\dpath/sub/_005_ ), .X(\dpath/sub/_061_ ) );
sky130_fd_sc_hs__nand2_1 \dpath/sub/_208_ ( .A(\dpath/sub/_060_ ), .B(\dpath/sub/_061_ ), .Y(\dpath/sub/_062_ ) );
sky130_fd_sc_hs__xnor3_1 \dpath/sub/_209_ ( .A(\dpath/sub/_006_ ), .B(\dpath/sub/_022_ ), .C(\dpath/sub/_062_ ), .X(\dpath/sub/_111_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_210_ ( .A(\dpath/a_lt_b$in0[0] ), .X(\dpath/sub/_000_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_211_ ( .A(\dpath/a_lt_b$in1[0] ), .X(\dpath/sub/_016_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_212_ ( .A(\dpath/sub/_105_ ), .X(\resp_msg[0] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_213_ ( .A(\dpath/a_lt_b$in0[1] ), .X(\dpath/sub/_007_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_214_ ( .A(\dpath/a_lt_b$in1[1] ), .X(\dpath/sub/_023_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_215_ ( .A(\dpath/sub/_112_ ), .X(\resp_msg[1] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_216_ ( .A(\dpath/a_lt_b$in0[2] ), .X(\dpath/sub/_008_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_217_ ( .A(\dpath/a_lt_b$in1[2] ), .X(\dpath/sub/_024_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_218_ ( .A(\dpath/sub/_113_ ), .X(\resp_msg[2] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_219_ ( .A(\dpath/a_lt_b$in0[3] ), .X(\dpath/sub/_009_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_220_ ( .A(\dpath/a_lt_b$in1[3] ), .X(\dpath/sub/_025_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_221_ ( .A(\dpath/sub/_114_ ), .X(\resp_msg[3] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_222_ ( .A(\dpath/a_lt_b$in0[4] ), .X(\dpath/sub/_010_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_223_ ( .A(\dpath/a_lt_b$in1[4] ), .X(\dpath/sub/_026_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_224_ ( .A(\dpath/sub/_115_ ), .X(\resp_msg[4] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_225_ ( .A(\dpath/a_lt_b$in0[5] ), .X(\dpath/sub/_011_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_226_ ( .A(\dpath/a_lt_b$in1[5] ), .X(\dpath/sub/_027_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_227_ ( .A(\dpath/sub/_116_ ), .X(\resp_msg[5] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_228_ ( .A(\dpath/a_lt_b$in0[6] ), .X(\dpath/sub/_012_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_229_ ( .A(\dpath/a_lt_b$in1[6] ), .X(\dpath/sub/_028_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_230_ ( .A(\dpath/sub/_117_ ), .X(\resp_msg[6] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_231_ ( .A(\dpath/a_lt_b$in0[7] ), .X(\dpath/sub/_013_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_232_ ( .A(\dpath/a_lt_b$in1[7] ), .X(\dpath/sub/_029_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_233_ ( .A(\dpath/sub/_118_ ), .X(\resp_msg[7] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_234_ ( .A(\dpath/a_lt_b$in0[8] ), .X(\dpath/sub/_014_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_235_ ( .A(\dpath/a_lt_b$in1[8] ), .X(\dpath/sub/_030_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_236_ ( .A(\dpath/sub/_119_ ), .X(\resp_msg[8] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_237_ ( .A(\dpath/a_lt_b$in0[9] ), .X(\dpath/sub/_015_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_238_ ( .A(\dpath/a_lt_b$in1[9] ), .X(\dpath/sub/_031_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_239_ ( .A(\dpath/sub/_120_ ), .X(\resp_msg[9] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_240_ ( .A(\dpath/a_lt_b$in0[10] ), .X(\dpath/sub/_001_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_241_ ( .A(\dpath/a_lt_b$in1[10] ), .X(\dpath/sub/_017_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_242_ ( .A(\dpath/sub/_106_ ), .X(\resp_msg[10] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_243_ ( .A(\dpath/a_lt_b$in0[11] ), .X(\dpath/sub/_002_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_244_ ( .A(\dpath/a_lt_b$in1[11] ), .X(\dpath/sub/_018_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_245_ ( .A(\dpath/sub/_107_ ), .X(\resp_msg[11] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_246_ ( .A(\dpath/a_lt_b$in0[12] ), .X(\dpath/sub/_003_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_247_ ( .A(\dpath/a_lt_b$in1[12] ), .X(\dpath/sub/_019_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_248_ ( .A(\dpath/sub/_108_ ), .X(\resp_msg[12] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_249_ ( .A(\dpath/a_lt_b$in0[13] ), .X(\dpath/sub/_004_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_250_ ( .A(\dpath/a_lt_b$in1[13] ), .X(\dpath/sub/_020_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_251_ ( .A(\dpath/sub/_109_ ), .X(\resp_msg[13] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_252_ ( .A(\dpath/a_lt_b$in0[14] ), .X(\dpath/sub/_005_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_253_ ( .A(\dpath/a_lt_b$in1[14] ), .X(\dpath/sub/_021_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_254_ ( .A(\dpath/sub/_110_ ), .X(\resp_msg[14] ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_255_ ( .A(\dpath/a_lt_b$in0[15] ), .X(\dpath/sub/_006_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_256_ ( .A(\dpath/a_lt_b$in1[15] ), .X(\dpath/sub/_022_ ) );
sky130_fd_sc_hs__buf_1 \dpath/sub/_257_ ( .A(\dpath/sub/_111_ ), .X(\resp_msg[15] ) );
sky130_fd_sc_hs__buf_1 clk_86_buf ( .A(clk_61 ), .X(clk_86 ) );
sky130_fd_sc_hs__buf_1 clk_85_buf ( .A(clk_60 ), .X(clk_85 ) );
sky130_fd_sc_hs__buf_1 clk_84_buf ( .A(clk_59 ), .X(clk_84 ) );
sky130_fd_sc_hs__buf_1 clk_83_buf ( .A(clk_59 ), .X(clk_83 ) );
sky130_fd_sc_hs__buf_1 clk_82_buf ( .A(clk_56 ), .X(clk_82 ) );
sky130_fd_sc_hs__buf_1 clk_81_buf ( .A(clk_55 ), .X(clk_81 ) );
sky130_fd_sc_hs__buf_1 clk_80_buf ( .A(clk_55 ), .X(clk_80 ) );
sky130_fd_sc_hs__buf_1 clk_79_buf ( .A(clk_54 ), .X(clk_79 ) );
sky130_fd_sc_hs__buf_1 clk_78_buf ( .A(clk_54 ), .X(clk_78 ) );
sky130_fd_sc_hs__buf_1 clk_77_buf ( .A(clk_53 ), .X(clk_77 ) );
sky130_fd_sc_hs__buf_1 clk_76_buf ( .A(clk_52 ), .X(clk_76 ) );
sky130_fd_sc_hs__buf_1 clk_75_buf ( .A(clk_51 ), .X(clk_75 ) );
sky130_fd_sc_hs__buf_1 clk_74_buf ( .A(clk_51 ), .X(clk_74 ) );
sky130_fd_sc_hs__buf_1 clk_73_buf ( .A(clk_50 ), .X(clk_73 ) );
sky130_fd_sc_hs__buf_1 clk_72_buf ( .A(clk_50 ), .X(clk_72 ) );
sky130_fd_sc_hs__buf_1 clk_71_buf ( .A(clk_49 ), .X(clk_71 ) );
sky130_fd_sc_hs__buf_1 clk_70_buf ( .A(clk_49 ), .X(clk_70 ) );
sky130_fd_sc_hs__buf_1 clk_69_buf ( .A(clk_48 ), .X(clk_69 ) );
sky130_fd_sc_hs__buf_1 clk_68_buf ( .A(clk_48 ), .X(clk_68 ) );
sky130_fd_sc_hs__buf_1 clk_67_buf ( .A(clk_47 ), .X(clk_67 ) );
sky130_fd_sc_hs__buf_1 clk_66_buf ( .A(clk_47 ), .X(clk_66 ) );
sky130_fd_sc_hs__buf_1 clk_65_buf ( .A(clk_46 ), .X(clk_65 ) );
sky130_fd_sc_hs__buf_1 clk_64_buf ( .A(clk_46 ), .X(clk_64 ) );
sky130_fd_sc_hs__buf_1 clk_63_buf ( .A(clk_45 ), .X(clk_63 ) );
sky130_fd_sc_hs__buf_1 clk_62_buf ( .A(clk_44 ), .X(clk_62 ) );
sky130_fd_sc_hs__buf_1 clk_61_buf ( .A(clk_43 ), .X(clk_61 ) );
sky130_fd_sc_hs__buf_1 clk_60_buf ( .A(clk_43 ), .X(clk_60 ) );
sky130_fd_sc_hs__buf_1 clk_59_buf ( .A(clk_42 ), .X(clk_59 ) );
sky130_fd_sc_hs__buf_1 clk_58_buf ( .A(clk_41 ), .X(clk_58 ) );
sky130_fd_sc_hs__buf_1 clk_57_buf ( .A(clk_40 ), .X(clk_57 ) );
sky130_fd_sc_hs__buf_1 clk_56_buf ( .A(clk_39 ), .X(clk_56 ) );
sky130_fd_sc_hs__buf_1 clk_55_buf ( .A(clk_38 ), .X(clk_55 ) );
sky130_fd_sc_hs__buf_1 clk_54_buf ( .A(clk_37 ), .X(clk_54 ) );
sky130_fd_sc_hs__buf_1 clk_53_buf ( .A(clk_36 ), .X(clk_53 ) );
sky130_fd_sc_hs__buf_1 clk_52_buf ( .A(clk_36 ), .X(clk_52 ) );
sky130_fd_sc_hs__buf_1 clk_51_buf ( .A(clk_35 ), .X(clk_51 ) );
sky130_fd_sc_hs__buf_1 clk_50_buf ( .A(clk_35 ), .X(clk_50 ) );
sky130_fd_sc_hs__buf_1 clk_49_buf ( .A(clk_34 ), .X(clk_49 ) );
sky130_fd_sc_hs__buf_1 clk_48_buf ( .A(clk_34 ), .X(clk_48 ) );
sky130_fd_sc_hs__buf_1 clk_47_buf ( .A(clk_33 ), .X(clk_47 ) );
sky130_fd_sc_hs__buf_1 clk_46_buf ( .A(clk_33 ), .X(clk_46 ) );
sky130_fd_sc_hs__buf_1 clk_45_buf ( .A(clk_32 ), .X(clk_45 ) );
sky130_fd_sc_hs__buf_1 clk_44_buf ( .A(clk_32 ), .X(clk_44 ) );
sky130_fd_sc_hs__buf_1 clk_43_buf ( .A(clk_31 ), .X(clk_43 ) );
sky130_fd_sc_hs__buf_1 clk_42_buf ( .A(clk_30 ), .X(clk_42 ) );
sky130_fd_sc_hs__buf_1 clk_41_buf ( .A(clk_29 ), .X(clk_41 ) );
sky130_fd_sc_hs__buf_1 clk_40_buf ( .A(clk_29 ), .X(clk_40 ) );
sky130_fd_sc_hs__buf_1 clk_39_buf ( .A(clk_28 ), .X(clk_39 ) );
sky130_fd_sc_hs__buf_1 clk_38_buf ( .A(clk_27 ), .X(clk_38 ) );
sky130_fd_sc_hs__buf_1 clk_37_buf ( .A(clk_27 ), .X(clk_37 ) );
sky130_fd_sc_hs__buf_1 clk_36_buf ( .A(clk_26 ), .X(clk_36 ) );
sky130_fd_sc_hs__buf_1 clk_35_buf ( .A(clk_25 ), .X(clk_35 ) );
sky130_fd_sc_hs__buf_1 clk_34_buf ( .A(clk_24 ), .X(clk_34 ) );
sky130_fd_sc_hs__buf_1 clk_33_buf ( .A(clk_23 ), .X(clk_33 ) );
sky130_fd_sc_hs__buf_1 clk_32_buf ( .A(clk_22 ), .X(clk_32 ) );
sky130_fd_sc_hs__buf_1 clk_31_buf ( .A(clk_21 ), .X(clk_31 ) );
sky130_fd_sc_hs__buf_1 clk_30_buf ( .A(clk_20 ), .X(clk_30 ) );
sky130_fd_sc_hs__buf_1 clk_29_buf ( .A(clk_19 ), .X(clk_29 ) );
sky130_fd_sc_hs__buf_1 clk_28_buf ( .A(clk_18 ), .X(clk_28 ) );
sky130_fd_sc_hs__buf_1 clk_27_buf ( .A(clk_17 ), .X(clk_27 ) );
sky130_fd_sc_hs__buf_1 clk_26_buf ( .A(clk_17 ), .X(clk_26 ) );
sky130_fd_sc_hs__buf_1 clk_25_buf ( .A(clk_16 ), .X(clk_25 ) );
sky130_fd_sc_hs__buf_1 clk_24_buf ( .A(clk_16 ), .X(clk_24 ) );
sky130_fd_sc_hs__buf_1 clk_23_buf ( .A(clk_15 ), .X(clk_23 ) );
sky130_fd_sc_hs__buf_1 clk_22_buf ( .A(clk_15 ), .X(clk_22 ) );
sky130_fd_sc_hs__buf_1 clk_21_buf ( .A(clk_14 ), .X(clk_21 ) );
sky130_fd_sc_hs__buf_1 clk_20_buf ( .A(clk_14 ), .X(clk_20 ) );
sky130_fd_sc_hs__buf_1 clk_19_buf ( .A(clk_13 ), .X(clk_19 ) );
sky130_fd_sc_hs__buf_1 clk_18_buf ( .A(clk_13 ), .X(clk_18 ) );
sky130_fd_sc_hs__buf_1 clk_17_buf ( .A(clk_12 ), .X(clk_17 ) );
sky130_fd_sc_hs__buf_1 clk_16_buf ( .A(clk_11 ), .X(clk_16 ) );
sky130_fd_sc_hs__buf_1 clk_15_buf ( .A(clk_10 ), .X(clk_15 ) );
sky130_fd_sc_hs__buf_1 clk_14_buf ( .A(clk_9 ), .X(clk_14 ) );
sky130_fd_sc_hs__buf_1 clk_13_buf ( .A(clk_8 ), .X(clk_13 ) );
sky130_fd_sc_hs__buf_1 clk_12_buf ( .A(clk_7 ), .X(clk_12 ) );
sky130_fd_sc_hs__buf_1 clk_11_buf ( .A(clk_6 ), .X(clk_11 ) );
sky130_fd_sc_hs__buf_1 clk_10_buf ( .A(clk_6 ), .X(clk_10 ) );
sky130_fd_sc_hs__buf_1 clk_9_buf ( .A(clk_5 ), .X(clk_9 ) );
sky130_fd_sc_hs__buf_1 clk_8_buf ( .A(clk_5 ), .X(clk_8 ) );
sky130_fd_sc_hs__buf_1 clk_7_buf ( .A(clk_4 ), .X(clk_7 ) );
sky130_fd_sc_hs__buf_1 clk_6_buf ( .A(clk_3 ), .X(clk_6 ) );
sky130_fd_sc_hs__buf_1 clk_5_buf ( .A(clk_2 ), .X(clk_5 ) );
sky130_fd_sc_hs__buf_1 clk_4_buf ( .A(clk_2 ), .X(clk_4 ) );
sky130_fd_sc_hs__buf_1 clk_3_buf ( .A(clk_1 ), .X(clk_3 ) );
sky130_fd_sc_hs__buf_1 clk_2_buf ( .A(clk_0 ), .X(clk_2 ) );
sky130_fd_sc_hs__buf_1 clk_1_buf ( .A(clk_0 ), .X(clk_1 ) );
sky130_fd_sc_hs__buf_1 clk_0_buf ( .A(clk ), .X(clk_0 ) );

endmodule
