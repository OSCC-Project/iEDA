module aes_cipher_top (
clk,
done,
ld,
rst,
key,
text_in,
text_out
);

input clk ;
output done ;
input ld ;
input rst ;
input [127:0] key ;
input [127:0] text_in ;
output [127:0] text_out ;

wire FE_OFN0_text_out_80 ;
wire CTS_23 ;
wire CTS_22 ;
wire CTS_19 ;
wire CTS_18 ;
wire CTS_21 ;
wire CTS_20 ;
wire CTS_15 ;
wire CTS_14 ;
wire CTS_17 ;
wire CTS_16 ;
wire CTS_13 ;
wire CTS_10 ;
wire CTS_9 ;
wire CTS_12 ;
wire CTS_11 ;
wire CTS_6 ;
wire CTS_5 ;
wire CTS_8 ;
wire CTS_7 ;
wire CTS_2 ;
wire CTS_1 ;
wire CTS_4 ;
wire CTS_3 ;
wire clk ;
wire done ;
wire ld ;
wire rst ;
wire _0164_ ;
wire _0261_ ;
wire _0262_ ;
wire _0263_ ;
wire _0264_ ;
wire _0265_ ;
wire _0266_ ;
wire _0267_ ;
wire _0268_ ;
wire _0269_ ;
wire _0270_ ;
wire _0271_ ;
wire _0272_ ;
wire _0273_ ;
wire _0274_ ;
wire _0275_ ;
wire _0276_ ;
wire _0277_ ;
wire _0278_ ;
wire _0279_ ;
wire _0280_ ;
wire _0281_ ;
wire _0282_ ;
wire _0283_ ;
wire _0284_ ;
wire _0285_ ;
wire _0286_ ;
wire _0287_ ;
wire _0288_ ;
wire _0289_ ;
wire _0290_ ;
wire _0291_ ;
wire _0292_ ;
wire _0293_ ;
wire _0294_ ;
wire _0295_ ;
wire _0296_ ;
wire _0297_ ;
wire _0298_ ;
wire _0299_ ;
wire _0300_ ;
wire _0301_ ;
wire _0302_ ;
wire _0303_ ;
wire _0304_ ;
wire _0305_ ;
wire _0306_ ;
wire _0307_ ;
wire _0308_ ;
wire _0309_ ;
wire _0310_ ;
wire _0311_ ;
wire _0312_ ;
wire _0313_ ;
wire _0314_ ;
wire _0315_ ;
wire _0316_ ;
wire _0317_ ;
wire _0318_ ;
wire _0319_ ;
wire _0320_ ;
wire _0321_ ;
wire _0322_ ;
wire _0323_ ;
wire _0324_ ;
wire _0325_ ;
wire _0326_ ;
wire _0327_ ;
wire _0328_ ;
wire _0329_ ;
wire _0330_ ;
wire _0331_ ;
wire _0332_ ;
wire _0333_ ;
wire _0334_ ;
wire _0335_ ;
wire _0336_ ;
wire _0337_ ;
wire _0338_ ;
wire _0339_ ;
wire _0340_ ;
wire _0341_ ;
wire _0342_ ;
wire _0343_ ;
wire _0344_ ;
wire _0345_ ;
wire _0346_ ;
wire _0347_ ;
wire _0348_ ;
wire _0349_ ;
wire _0350_ ;
wire _0351_ ;
wire _0352_ ;
wire _0353_ ;
wire _0354_ ;
wire _0355_ ;
wire _0356_ ;
wire _0357_ ;
wire _0358_ ;
wire _0359_ ;
wire _0360_ ;
wire _0361_ ;
wire _0362_ ;
wire _0363_ ;
wire _0364_ ;
wire _0365_ ;
wire _0366_ ;
wire _0367_ ;
wire _0368_ ;
wire _0369_ ;
wire _0370_ ;
wire _0371_ ;
wire _0372_ ;
wire _0373_ ;
wire _0374_ ;
wire _0375_ ;
wire _0376_ ;
wire _0377_ ;
wire _0378_ ;
wire _0379_ ;
wire _0380_ ;
wire _0381_ ;
wire _0382_ ;
wire _0383_ ;
wire _0384_ ;
wire _0385_ ;
wire _0386_ ;
wire _0387_ ;
wire _0388_ ;
wire _0389_ ;
wire _0390_ ;
wire _0391_ ;
wire _0392_ ;
wire _0393_ ;
wire _0394_ ;
wire _0395_ ;
wire _0396_ ;
wire _0397_ ;
wire _0398_ ;
wire _0399_ ;
wire _0400_ ;
wire _0401_ ;
wire _0402_ ;
wire _0403_ ;
wire _0404_ ;
wire _0405_ ;
wire _0406_ ;
wire _0407_ ;
wire _0408_ ;
wire _0409_ ;
wire _0410_ ;
wire _0411_ ;
wire _0412_ ;
wire _0413_ ;
wire _0414_ ;
wire _0415_ ;
wire _0416_ ;
wire _0417_ ;
wire _0418_ ;
wire _0419_ ;
wire _0420_ ;
wire _0421_ ;
wire _0422_ ;
wire _0423_ ;
wire _0424_ ;
wire _0425_ ;
wire _0426_ ;
wire _0427_ ;
wire _0428_ ;
wire _0429_ ;
wire _0430_ ;
wire _0431_ ;
wire _0432_ ;
wire _0433_ ;
wire _0434_ ;
wire _0435_ ;
wire _0436_ ;
wire _0437_ ;
wire _0438_ ;
wire _0439_ ;
wire _0440_ ;
wire _0441_ ;
wire _0442_ ;
wire _0443_ ;
wire _0444_ ;
wire _0445_ ;
wire _0446_ ;
wire _0447_ ;
wire _0448_ ;
wire _0449_ ;
wire _0450_ ;
wire _0451_ ;
wire _0452_ ;
wire _0453_ ;
wire _0454_ ;
wire _0455_ ;
wire _0456_ ;
wire _0457_ ;
wire _0458_ ;
wire _0459_ ;
wire _0460_ ;
wire _0461_ ;
wire _0462_ ;
wire _0463_ ;
wire _0464_ ;
wire _0465_ ;
wire _0466_ ;
wire _0467_ ;
wire _0468_ ;
wire _0469_ ;
wire _0470_ ;
wire _0471_ ;
wire _0472_ ;
wire _0473_ ;
wire _0474_ ;
wire _0475_ ;
wire _0476_ ;
wire _0477_ ;
wire _0478_ ;
wire _0479_ ;
wire _0480_ ;
wire _0481_ ;
wire _0482_ ;
wire _0483_ ;
wire _0484_ ;
wire _0485_ ;
wire _0486_ ;
wire _0487_ ;
wire _0488_ ;
wire _0489_ ;
wire _0490_ ;
wire _0491_ ;
wire _0492_ ;
wire _0493_ ;
wire _0494_ ;
wire _0495_ ;
wire _0496_ ;
wire _0497_ ;
wire _0498_ ;
wire _0499_ ;
wire _0500_ ;
wire _0501_ ;
wire _0502_ ;
wire _0503_ ;
wire _0504_ ;
wire _0505_ ;
wire _0506_ ;
wire _0507_ ;
wire _0508_ ;
wire _0509_ ;
wire _0510_ ;
wire _0511_ ;
wire _0512_ ;
wire _0513_ ;
wire _0514_ ;
wire _0515_ ;
wire _0516_ ;
wire _0517_ ;
wire _0518_ ;
wire _0519_ ;
wire _0520_ ;
wire _0521_ ;
wire _0529_ ;
wire _0530_ ;
wire _0531_ ;
wire _0532_ ;
wire _0533_ ;
wire _0534_ ;
wire _0535_ ;
wire _0536_ ;
wire _0537_ ;
wire _0538_ ;
wire _0539_ ;
wire _0541_ ;
wire _0542_ ;
wire _0543_ ;
wire _0544_ ;
wire _0545_ ;
wire _0546_ ;
wire _0547_ ;
wire _0548_ ;
wire _0549_ ;
wire _0550_ ;
wire _0551_ ;
wire _0552_ ;
wire _0554_ ;
wire _0555_ ;
wire _0556_ ;
wire _0557_ ;
wire _0558_ ;
wire _0559_ ;
wire _0560_ ;
wire _0561_ ;
wire _0562_ ;
wire _0563_ ;
wire _0564_ ;
wire _0565_ ;
wire _0566_ ;
wire _0567_ ;
wire _0568_ ;
wire _0569_ ;
wire _0570_ ;
wire _0571_ ;
wire _0572_ ;
wire _0573_ ;
wire _0574_ ;
wire _0575_ ;
wire _0576_ ;
wire _0577_ ;
wire _0578_ ;
wire _0579_ ;
wire _0580_ ;
wire _0581_ ;
wire _0582_ ;
wire _0583_ ;
wire _0584_ ;
wire _0585_ ;
wire _0586_ ;
wire _0587_ ;
wire _0588_ ;
wire _0589_ ;
wire _0591_ ;
wire _0592_ ;
wire _0593_ ;
wire _0594_ ;
wire _0595_ ;
wire _0596_ ;
wire _0597_ ;
wire _0598_ ;
wire _0599_ ;
wire _0600_ ;
wire _0601_ ;
wire _0602_ ;
wire _0603_ ;
wire _0604_ ;
wire _0605_ ;
wire _0606_ ;
wire _0607_ ;
wire _0608_ ;
wire _0609_ ;
wire _0610_ ;
wire _0611_ ;
wire _0612_ ;
wire _0613_ ;
wire _0614_ ;
wire _0615_ ;
wire _0616_ ;
wire _0617_ ;
wire _0618_ ;
wire _0619_ ;
wire _0620_ ;
wire _0621_ ;
wire _0622_ ;
wire _0623_ ;
wire _0624_ ;
wire _0625_ ;
wire _0626_ ;
wire _0627_ ;
wire _0628_ ;
wire _0629_ ;
wire _0630_ ;
wire _0631_ ;
wire _0632_ ;
wire _0633_ ;
wire _0634_ ;
wire _0635_ ;
wire _0636_ ;
wire _0637_ ;
wire _0638_ ;
wire _0639_ ;
wire _0640_ ;
wire _0641_ ;
wire _0643_ ;
wire _0644_ ;
wire _0645_ ;
wire _0646_ ;
wire _0647_ ;
wire _0648_ ;
wire _0649_ ;
wire _0650_ ;
wire _0651_ ;
wire _0652_ ;
wire _0653_ ;
wire _0654_ ;
wire _0655_ ;
wire _0656_ ;
wire _0657_ ;
wire _0658_ ;
wire _0659_ ;
wire _0660_ ;
wire _0661_ ;
wire _0662_ ;
wire _0663_ ;
wire _0664_ ;
wire _0665_ ;
wire _0666_ ;
wire _0667_ ;
wire _0668_ ;
wire _0669_ ;
wire _0670_ ;
wire _0671_ ;
wire _0672_ ;
wire _0673_ ;
wire _0674_ ;
wire _0675_ ;
wire _0676_ ;
wire _0677_ ;
wire _0678_ ;
wire _0679_ ;
wire _0680_ ;
wire _0681_ ;
wire _0682_ ;
wire _0683_ ;
wire _0684_ ;
wire _0685_ ;
wire _0686_ ;
wire _0687_ ;
wire _0688_ ;
wire _0689_ ;
wire _0690_ ;
wire _0691_ ;
wire _0692_ ;
wire _0693_ ;
wire _0694_ ;
wire _0695_ ;
wire _0696_ ;
wire _0697_ ;
wire _0698_ ;
wire _0699_ ;
wire _0700_ ;
wire _0701_ ;
wire _0702_ ;
wire _0704_ ;
wire _0705_ ;
wire _0706_ ;
wire _0707_ ;
wire _0708_ ;
wire _0709_ ;
wire _0710_ ;
wire _0711_ ;
wire _0712_ ;
wire _0713_ ;
wire _0714_ ;
wire _0715_ ;
wire _0716_ ;
wire _0717_ ;
wire _0718_ ;
wire _0719_ ;
wire _0720_ ;
wire _0721_ ;
wire _0722_ ;
wire _0723_ ;
wire _0724_ ;
wire _0725_ ;
wire _0726_ ;
wire _0727_ ;
wire _0728_ ;
wire _0729_ ;
wire _0730_ ;
wire _0731_ ;
wire _0732_ ;
wire _0733_ ;
wire _0734_ ;
wire _0735_ ;
wire _0736_ ;
wire _0737_ ;
wire _0738_ ;
wire _0739_ ;
wire _0740_ ;
wire _0741_ ;
wire _0742_ ;
wire _0743_ ;
wire _0744_ ;
wire _0745_ ;
wire _0746_ ;
wire _0747_ ;
wire _0748_ ;
wire _0749_ ;
wire _0750_ ;
wire _0751_ ;
wire _0752_ ;
wire _0753_ ;
wire _0754_ ;
wire _0755_ ;
wire _0756_ ;
wire _0758_ ;
wire _0759_ ;
wire _0760_ ;
wire _0761_ ;
wire _0762_ ;
wire _0763_ ;
wire _0764_ ;
wire _0765_ ;
wire _0766_ ;
wire _0767_ ;
wire _0768_ ;
wire _0769_ ;
wire _0770_ ;
wire _0771_ ;
wire _0772_ ;
wire _0773_ ;
wire _0774_ ;
wire _0775_ ;
wire _0776_ ;
wire _0777_ ;
wire _0778_ ;
wire _0779_ ;
wire _0780_ ;
wire _0781_ ;
wire _0782_ ;
wire _0783_ ;
wire _0784_ ;
wire _0785_ ;
wire _0786_ ;
wire _0787_ ;
wire _0788_ ;
wire _0789_ ;
wire _0790_ ;
wire _0791_ ;
wire _0792_ ;
wire _0793_ ;
wire _0794_ ;
wire _0795_ ;
wire _0796_ ;
wire _0797_ ;
wire _0798_ ;
wire _0799_ ;
wire _0800_ ;
wire _0801_ ;
wire _0802_ ;
wire _0803_ ;
wire _0805_ ;
wire _0806_ ;
wire _0807_ ;
wire _0808_ ;
wire _0809_ ;
wire _0810_ ;
wire _0811_ ;
wire _0812_ ;
wire _0813_ ;
wire _0814_ ;
wire _0815_ ;
wire _0816_ ;
wire _0817_ ;
wire _0818_ ;
wire _0819_ ;
wire _0820_ ;
wire _0821_ ;
wire _0822_ ;
wire _0823_ ;
wire _0824_ ;
wire _0825_ ;
wire _0826_ ;
wire _0827_ ;
wire _0828_ ;
wire _0829_ ;
wire _0830_ ;
wire _0831_ ;
wire _0832_ ;
wire _0833_ ;
wire _0834_ ;
wire _0835_ ;
wire _0836_ ;
wire _0837_ ;
wire _0838_ ;
wire _0839_ ;
wire _0840_ ;
wire _0841_ ;
wire _0842_ ;
wire _0843_ ;
wire _0844_ ;
wire _0845_ ;
wire _0846_ ;
wire _0847_ ;
wire _0848_ ;
wire _0849_ ;
wire _0850_ ;
wire _0851_ ;
wire _0852_ ;
wire _0853_ ;
wire _0854_ ;
wire _0855_ ;
wire _0856_ ;
wire _0857_ ;
wire _0858_ ;
wire _0859_ ;
wire _0860_ ;
wire _0861_ ;
wire _0862_ ;
wire _0863_ ;
wire _0864_ ;
wire _0865_ ;
wire _0866_ ;
wire _0867_ ;
wire _0868_ ;
wire _0869_ ;
wire _0870_ ;
wire _0871_ ;
wire _0872_ ;
wire _0873_ ;
wire _0874_ ;
wire _0875_ ;
wire _0876_ ;
wire _0877_ ;
wire _0878_ ;
wire _0879_ ;
wire _0880_ ;
wire _0881_ ;
wire _0882_ ;
wire _0883_ ;
wire _0884_ ;
wire _0885_ ;
wire _0886_ ;
wire _0887_ ;
wire _0888_ ;
wire _0889_ ;
wire _0890_ ;
wire _0891_ ;
wire _0892_ ;
wire _0893_ ;
wire _0894_ ;
wire _0895_ ;
wire _0896_ ;
wire _0897_ ;
wire _0898_ ;
wire _0899_ ;
wire _0900_ ;
wire _0901_ ;
wire _0902_ ;
wire _0903_ ;
wire _0904_ ;
wire _0905_ ;
wire _0906_ ;
wire _0907_ ;
wire _0908_ ;
wire _0909_ ;
wire _0910_ ;
wire _0911_ ;
wire _0912_ ;
wire _0913_ ;
wire _0914_ ;
wire _0915_ ;
wire _0916_ ;
wire _0917_ ;
wire _0918_ ;
wire _0919_ ;
wire _0920_ ;
wire _0921_ ;
wire _0922_ ;
wire _0923_ ;
wire _0924_ ;
wire _0925_ ;
wire _0926_ ;
wire _0927_ ;
wire _0928_ ;
wire _0929_ ;
wire _0930_ ;
wire _0931_ ;
wire _0932_ ;
wire _0933_ ;
wire _0934_ ;
wire _0935_ ;
wire _0936_ ;
wire _0937_ ;
wire _0938_ ;
wire _0939_ ;
wire _0940_ ;
wire _0941_ ;
wire _0942_ ;
wire _0943_ ;
wire _0944_ ;
wire _0945_ ;
wire _0946_ ;
wire _0947_ ;
wire _0948_ ;
wire _0949_ ;
wire _0950_ ;
wire _0951_ ;
wire _0952_ ;
wire _0953_ ;
wire _0954_ ;
wire _0955_ ;
wire _0956_ ;
wire _0957_ ;
wire _0958_ ;
wire _0959_ ;
wire _0960_ ;
wire _0961_ ;
wire _0962_ ;
wire _0963_ ;
wire _0964_ ;
wire _0965_ ;
wire _0966_ ;
wire _0967_ ;
wire _0968_ ;
wire _0969_ ;
wire _0970_ ;
wire _0971_ ;
wire _0972_ ;
wire _0973_ ;
wire _0974_ ;
wire _0975_ ;
wire _0976_ ;
wire _0977_ ;
wire _0978_ ;
wire _0979_ ;
wire _0980_ ;
wire _0981_ ;
wire _0982_ ;
wire _0983_ ;
wire _0984_ ;
wire _0985_ ;
wire _0986_ ;
wire _0987_ ;
wire _0988_ ;
wire _0989_ ;
wire _0990_ ;
wire _0991_ ;
wire _0992_ ;
wire _0993_ ;
wire _0994_ ;
wire _0995_ ;
wire _0996_ ;
wire _0997_ ;
wire _0998_ ;
wire _0999_ ;
wire _1000_ ;
wire _1001_ ;
wire _1002_ ;
wire _1003_ ;
wire _1004_ ;
wire _1005_ ;
wire _1006_ ;
wire _1007_ ;
wire _1008_ ;
wire _1009_ ;
wire _1010_ ;
wire _1011_ ;
wire _1012_ ;
wire _1013_ ;
wire _1014_ ;
wire _1015_ ;
wire _1016_ ;
wire _1017_ ;
wire _1018_ ;
wire _1019_ ;
wire _1020_ ;
wire _1021_ ;
wire _1022_ ;
wire _1023_ ;
wire _1024_ ;
wire _1025_ ;
wire _1026_ ;
wire _1027_ ;
wire _1028_ ;
wire _1029_ ;
wire _1030_ ;
wire _1031_ ;
wire _1032_ ;
wire _1033_ ;
wire _1034_ ;
wire _1035_ ;
wire _1036_ ;
wire _1037_ ;
wire _1038_ ;
wire _1039_ ;
wire _1040_ ;
wire _1041_ ;
wire _1042_ ;
wire _1043_ ;
wire _1044_ ;
wire _1045_ ;
wire _1046_ ;
wire _1047_ ;
wire _1048_ ;
wire _1049_ ;
wire _1050_ ;
wire _1051_ ;
wire _1052_ ;
wire _1053_ ;
wire _1054_ ;
wire _1055_ ;
wire _1056_ ;
wire _1057_ ;
wire _1058_ ;
wire _1059_ ;
wire _1060_ ;
wire _1061_ ;
wire _1062_ ;
wire _1063_ ;
wire _1064_ ;
wire _1065_ ;
wire _1066_ ;
wire _1067_ ;
wire _1068_ ;
wire _1069_ ;
wire _1070_ ;
wire _1071_ ;
wire _1072_ ;
wire _1073_ ;
wire _1074_ ;
wire _1075_ ;
wire _1076_ ;
wire _1077_ ;
wire _1078_ ;
wire _1079_ ;
wire _1080_ ;
wire _1081_ ;
wire _1082_ ;
wire _1083_ ;
wire _1084_ ;
wire _1085_ ;
wire _1086_ ;
wire _1087_ ;
wire _1088_ ;
wire _1089_ ;
wire _1090_ ;
wire _1091_ ;
wire _1092_ ;
wire _1093_ ;
wire _1094_ ;
wire _1095_ ;
wire _1096_ ;
wire _1097_ ;
wire _1098_ ;
wire _1099_ ;
wire _1100_ ;
wire _1101_ ;
wire _1102_ ;
wire _1103_ ;
wire _1104_ ;
wire _1105_ ;
wire _1106_ ;
wire _1107_ ;
wire _1108_ ;
wire _1109_ ;
wire _1110_ ;
wire _1111_ ;
wire _1112_ ;
wire _1113_ ;
wire _1114_ ;
wire _1115_ ;
wire _1116_ ;
wire _1117_ ;
wire _1118_ ;
wire _1119_ ;
wire _1120_ ;
wire _1121_ ;
wire _1122_ ;
wire _1123_ ;
wire _1124_ ;
wire _1125_ ;
wire _1126_ ;
wire _1127_ ;
wire _1128_ ;
wire _1129_ ;
wire _1130_ ;
wire _1131_ ;
wire _1132_ ;
wire _1133_ ;
wire _1134_ ;
wire _1135_ ;
wire _1136_ ;
wire _1137_ ;
wire _1138_ ;
wire _1139_ ;
wire _1140_ ;
wire _1141_ ;
wire _1142_ ;
wire _1143_ ;
wire _1144_ ;
wire _1145_ ;
wire _1146_ ;
wire _1147_ ;
wire _1148_ ;
wire _1149_ ;
wire _1150_ ;
wire _1151_ ;
wire _1152_ ;
wire _1153_ ;
wire _1154_ ;
wire _1155_ ;
wire _1156_ ;
wire _1157_ ;
wire _1158_ ;
wire _1159_ ;
wire _1160_ ;
wire _1161_ ;
wire _1162_ ;
wire _1163_ ;
wire _1164_ ;
wire _1165_ ;
wire _1166_ ;
wire _1167_ ;
wire _1168_ ;
wire _1169_ ;
wire _1170_ ;
wire _1171_ ;
wire _1172_ ;
wire _1173_ ;
wire _1174_ ;
wire _1175_ ;
wire _1176_ ;
wire _1177_ ;
wire _1178_ ;
wire _1179_ ;
wire _1180_ ;
wire _1181_ ;
wire _1182_ ;
wire _1183_ ;
wire _1184_ ;
wire _1185_ ;
wire _1186_ ;
wire _1187_ ;
wire _1188_ ;
wire _1189_ ;
wire _1190_ ;
wire _1191_ ;
wire _1192_ ;
wire _1193_ ;
wire _1194_ ;
wire _1195_ ;
wire _1196_ ;
wire _1197_ ;
wire _1198_ ;
wire _1199_ ;
wire _1200_ ;
wire _1201_ ;
wire _1202_ ;
wire _1203_ ;
wire _1204_ ;
wire _1205_ ;
wire _1206_ ;
wire _1207_ ;
wire _1208_ ;
wire _1209_ ;
wire _1210_ ;
wire _1211_ ;
wire _1212_ ;
wire _1213_ ;
wire _1214_ ;
wire _1215_ ;
wire _1216_ ;
wire _1217_ ;
wire _1218_ ;
wire _1219_ ;
wire _1220_ ;
wire _1221_ ;
wire _1222_ ;
wire _1223_ ;
wire _1224_ ;
wire _1225_ ;
wire _1226_ ;
wire _1227_ ;
wire _1228_ ;
wire _1229_ ;
wire _1230_ ;
wire _1231_ ;
wire _1232_ ;
wire _1233_ ;
wire _1234_ ;
wire _1235_ ;
wire _1236_ ;
wire _1237_ ;
wire _1238_ ;
wire _1239_ ;
wire _1240_ ;
wire _1241_ ;
wire _1242_ ;
wire _1243_ ;
wire _1244_ ;
wire _1245_ ;
wire _1246_ ;
wire _1247_ ;
wire _1248_ ;
wire _1249_ ;
wire _1250_ ;
wire _1251_ ;
wire _1252_ ;
wire _1253_ ;
wire _1254_ ;
wire _1255_ ;
wire _1256_ ;
wire _1257_ ;
wire _1258_ ;
wire _1259_ ;
wire _1260_ ;
wire _1261_ ;
wire _1262_ ;
wire _1263_ ;
wire _1264_ ;
wire _1265_ ;
wire _1266_ ;
wire _1267_ ;
wire _1268_ ;
wire _1269_ ;
wire _1270_ ;
wire _1271_ ;
wire _1272_ ;
wire _1273_ ;
wire _1274_ ;
wire _1275_ ;
wire _1276_ ;
wire _1277_ ;
wire _1278_ ;
wire _1279_ ;
wire _1280_ ;
wire _1281_ ;
wire _1282_ ;
wire _1283_ ;
wire _1284_ ;
wire _1285_ ;
wire _1286_ ;
wire _1287_ ;
wire _1288_ ;
wire _1289_ ;
wire _1290_ ;
wire _1291_ ;
wire _1292_ ;
wire _1293_ ;
wire _1294_ ;
wire _1295_ ;
wire _1296_ ;
wire _1297_ ;
wire _1298_ ;
wire _1300_ ;
wire _1301_ ;
wire _1302_ ;
wire _1303_ ;
wire _1304_ ;
wire _1305_ ;
wire _1306_ ;
wire _1307_ ;
wire _1316_ ;
wire _1317_ ;
wire _1318_ ;
wire _1319_ ;
wire _1320_ ;
wire _1321_ ;
wire _1322_ ;
wire _1323_ ;
wire _1332_ ;
wire _1333_ ;
wire _1334_ ;
wire _1335_ ;
wire _1336_ ;
wire _1337_ ;
wire _1338_ ;
wire _1339_ ;
wire _1348_ ;
wire _1349_ ;
wire _1350_ ;
wire _1351_ ;
wire _1352_ ;
wire _1353_ ;
wire _1354_ ;
wire _1355_ ;
wire _1364_ ;
wire _1365_ ;
wire _1366_ ;
wire _1367_ ;
wire _1368_ ;
wire _1369_ ;
wire _1370_ ;
wire _1371_ ;
wire _1373_ ;
wire _1377_ ;
wire _1379_ ;
wire _1387_ ;
wire _1388_ ;
wire _1389_ ;
wire _1390_ ;
wire _1391_ ;
wire _1392_ ;
wire _1393_ ;
wire _1394_ ;
wire _1395_ ;
wire _1404_ ;
wire _1405_ ;
wire _1406_ ;
wire _1407_ ;
wire _1408_ ;
wire _1409_ ;
wire _1410_ ;
wire _1411_ ;
wire _1419_ ;
wire _1420_ ;
wire _1421_ ;
wire _1422_ ;
wire _1423_ ;
wire _1424_ ;
wire _1425_ ;
wire _1426_ ;
wire _1427_ ;
wire _1428_ ;
wire _1429_ ;
wire _1430_ ;
wire _1431_ ;
wire _1432_ ;
wire _1433_ ;
wire _1434_ ;
wire _1435_ ;
wire _1451_ ;
wire _1452_ ;
wire _1453_ ;
wire _1454_ ;
wire _1455_ ;
wire _1456_ ;
wire _1457_ ;
wire _1458_ ;
wire _1459_ ;
wire _1476_ ;
wire _1477_ ;
wire _1478_ ;
wire _1479_ ;
wire _1480_ ;
wire _1481_ ;
wire _1482_ ;
wire _1483_ ;
wire _1484_ ;
wire _1485_ ;
wire _1486_ ;
wire _1487_ ;
wire _1488_ ;
wire _1489_ ;
wire _1490_ ;
wire _1491_ ;
wire _1492_ ;
wire _1493_ ;
wire _1494_ ;
wire _1495_ ;
wire _1496_ ;
wire _1497_ ;
wire _1498_ ;
wire _1499_ ;
wire _1516_ ;
wire _1517_ ;
wire _1518_ ;
wire _1519_ ;
wire _1520_ ;
wire _1521_ ;
wire _1522_ ;
wire _1523_ ;
wire _1532_ ;
wire _1533_ ;
wire _1534_ ;
wire _1535_ ;
wire _1536_ ;
wire _1537_ ;
wire _1538_ ;
wire _1539_ ;
wire _1548_ ;
wire _1549_ ;
wire _1550_ ;
wire _1551_ ;
wire _1552_ ;
wire _1553_ ;
wire _1554_ ;
wire _1555_ ;
wire \dcnt[0] ;
wire \dcnt[1] ;
wire \dcnt[2] ;
wire \dcnt[3] ;
wire ld_r ;
wire net1 ;
wire net10 ;
wire net11 ;
wire net12 ;
wire net13 ;
wire net14 ;
wire net15 ;
wire net16 ;
wire net17 ;
wire net18 ;
wire net19 ;
wire net2 ;
wire net20 ;
wire net21 ;
wire net22 ;
wire net23 ;
wire net24 ;
wire net25 ;
wire net26 ;
wire net27 ;
wire net28 ;
wire net29 ;
wire net3 ;
wire net30 ;
wire net31 ;
wire net32 ;
wire net33 ;
wire net34 ;
wire net35 ;
wire net36 ;
wire net37 ;
wire net38 ;
wire net39 ;
wire net4 ;
wire net40 ;
wire net41 ;
wire net42 ;
wire net43 ;
wire net44 ;
wire net45 ;
wire net46 ;
wire net47 ;
wire net48 ;
wire net5 ;
wire net6 ;
wire net7 ;
wire net8 ;
wire net9 ;
wire \sa00[0] ;
wire \sa00[1] ;
wire \sa00[2] ;
wire \sa00[3] ;
wire \sa00[4] ;
wire \sa00[5] ;
wire \sa00[6] ;
wire \sa00[7] ;
wire \sa01[0] ;
wire \sa01[1] ;
wire \sa01[2] ;
wire \sa01[3] ;
wire \sa01[4] ;
wire \sa01[5] ;
wire \sa01[6] ;
wire \sa01[7] ;
wire \sa02[0] ;
wire \sa02[1] ;
wire \sa02[2] ;
wire \sa02[3] ;
wire \sa02[4] ;
wire \sa02[5] ;
wire \sa02[6] ;
wire \sa02[7] ;
wire \sa03[0] ;
wire \sa03[1] ;
wire \sa03[2] ;
wire \sa03[3] ;
wire \sa03[4] ;
wire \sa03[5] ;
wire \sa03[6] ;
wire \sa03[7] ;
wire \sa10[0] ;
wire \sa10[1] ;
wire \sa10[2] ;
wire \sa10[3] ;
wire \sa10[4] ;
wire \sa10[5] ;
wire \sa10[6] ;
wire \sa10[7] ;
wire \sa11[0] ;
wire \sa11[1] ;
wire \sa11[2] ;
wire \sa11[3] ;
wire \sa11[4] ;
wire \sa11[5] ;
wire \sa11[6] ;
wire \sa11[7] ;
wire \sa12[0] ;
wire \sa12[1] ;
wire \sa12[2] ;
wire \sa12[3] ;
wire \sa12[4] ;
wire \sa12[5] ;
wire \sa12[6] ;
wire \sa12[7] ;
wire \sa13[0] ;
wire \sa13[1] ;
wire \sa13[2] ;
wire \sa13[3] ;
wire \sa13[4] ;
wire \sa13[5] ;
wire \sa13[6] ;
wire \sa13[7] ;
wire \sa20[0] ;
wire \sa20[1] ;
wire \sa20[2] ;
wire \sa20[3] ;
wire \sa20[4] ;
wire \sa20[5] ;
wire \sa20[6] ;
wire \sa20[7] ;
wire \sa21[0] ;
wire \sa21[1] ;
wire \sa21[2] ;
wire \sa21[3] ;
wire \sa21[4] ;
wire \sa21[5] ;
wire \sa21[6] ;
wire \sa21[7] ;
wire \sa22[0] ;
wire \sa22[1] ;
wire \sa22[2] ;
wire \sa22[3] ;
wire \sa22[4] ;
wire \sa22[5] ;
wire \sa22[6] ;
wire \sa22[7] ;
wire \sa23[0] ;
wire \sa23[1] ;
wire \sa23[2] ;
wire \sa23[3] ;
wire \sa23[4] ;
wire \sa23[5] ;
wire \sa23[6] ;
wire \sa23[7] ;
wire \sa30[0] ;
wire \sa30[1] ;
wire \sa30[2] ;
wire \sa30[3] ;
wire \sa30[4] ;
wire \sa30[5] ;
wire \sa30[6] ;
wire \sa30[7] ;
wire \sa31[0] ;
wire \sa31[1] ;
wire \sa31[2] ;
wire \sa31[3] ;
wire \sa31[4] ;
wire \sa31[5] ;
wire \sa31[6] ;
wire \sa31[7] ;
wire \sa32[0] ;
wire \sa32[1] ;
wire \sa32[2] ;
wire \sa32[3] ;
wire \sa32[4] ;
wire \sa32[5] ;
wire \sa32[6] ;
wire \sa32[7] ;
wire \sa33[0] ;
wire \sa33[1] ;
wire \sa33[2] ;
wire \sa33[3] ;
wire \sa33[4] ;
wire \sa33[5] ;
wire \sa33[6] ;
wire \sa33[7] ;
wire \text_in_r[0] ;
wire \text_in_r[100] ;
wire \text_in_r[101] ;
wire \text_in_r[102] ;
wire \text_in_r[103] ;
wire \text_in_r[104] ;
wire \text_in_r[105] ;
wire \text_in_r[106] ;
wire \text_in_r[107] ;
wire \text_in_r[108] ;
wire \text_in_r[109] ;
wire \text_in_r[10] ;
wire \text_in_r[110] ;
wire \text_in_r[111] ;
wire \text_in_r[112] ;
wire \text_in_r[113] ;
wire \text_in_r[114] ;
wire \text_in_r[115] ;
wire \text_in_r[116] ;
wire \text_in_r[117] ;
wire \text_in_r[118] ;
wire \text_in_r[119] ;
wire \text_in_r[11] ;
wire \text_in_r[120] ;
wire \text_in_r[121] ;
wire \text_in_r[122] ;
wire \text_in_r[123] ;
wire \text_in_r[124] ;
wire \text_in_r[125] ;
wire \text_in_r[126] ;
wire \text_in_r[127] ;
wire \text_in_r[12] ;
wire \text_in_r[13] ;
wire \text_in_r[14] ;
wire \text_in_r[15] ;
wire \text_in_r[16] ;
wire \text_in_r[17] ;
wire \text_in_r[18] ;
wire \text_in_r[19] ;
wire \text_in_r[1] ;
wire \text_in_r[20] ;
wire \text_in_r[21] ;
wire \text_in_r[22] ;
wire \text_in_r[23] ;
wire \text_in_r[24] ;
wire \text_in_r[25] ;
wire \text_in_r[26] ;
wire \text_in_r[27] ;
wire \text_in_r[28] ;
wire \text_in_r[29] ;
wire \text_in_r[2] ;
wire \text_in_r[30] ;
wire \text_in_r[31] ;
wire \text_in_r[32] ;
wire \text_in_r[33] ;
wire \text_in_r[34] ;
wire \text_in_r[35] ;
wire \text_in_r[36] ;
wire \text_in_r[37] ;
wire \text_in_r[38] ;
wire \text_in_r[39] ;
wire \text_in_r[3] ;
wire \text_in_r[40] ;
wire \text_in_r[41] ;
wire \text_in_r[42] ;
wire \text_in_r[43] ;
wire \text_in_r[44] ;
wire \text_in_r[45] ;
wire \text_in_r[46] ;
wire \text_in_r[47] ;
wire \text_in_r[48] ;
wire \text_in_r[49] ;
wire \text_in_r[4] ;
wire \text_in_r[50] ;
wire \text_in_r[51] ;
wire \text_in_r[52] ;
wire \text_in_r[53] ;
wire \text_in_r[54] ;
wire \text_in_r[55] ;
wire \text_in_r[56] ;
wire \text_in_r[57] ;
wire \text_in_r[58] ;
wire \text_in_r[59] ;
wire \text_in_r[5] ;
wire \text_in_r[60] ;
wire \text_in_r[61] ;
wire \text_in_r[62] ;
wire \text_in_r[63] ;
wire \text_in_r[64] ;
wire \text_in_r[65] ;
wire \text_in_r[66] ;
wire \text_in_r[67] ;
wire \text_in_r[68] ;
wire \text_in_r[69] ;
wire \text_in_r[6] ;
wire \text_in_r[70] ;
wire \text_in_r[71] ;
wire \text_in_r[72] ;
wire \text_in_r[73] ;
wire \text_in_r[74] ;
wire \text_in_r[75] ;
wire \text_in_r[76] ;
wire \text_in_r[77] ;
wire \text_in_r[78] ;
wire \text_in_r[79] ;
wire \text_in_r[7] ;
wire \text_in_r[80] ;
wire \text_in_r[81] ;
wire \text_in_r[82] ;
wire \text_in_r[83] ;
wire \text_in_r[84] ;
wire \text_in_r[85] ;
wire \text_in_r[86] ;
wire \text_in_r[87] ;
wire \text_in_r[88] ;
wire \text_in_r[89] ;
wire \text_in_r[8] ;
wire \text_in_r[90] ;
wire \text_in_r[91] ;
wire \text_in_r[92] ;
wire \text_in_r[93] ;
wire \text_in_r[94] ;
wire \text_in_r[95] ;
wire \text_in_r[96] ;
wire \text_in_r[97] ;
wire \text_in_r[98] ;
wire \text_in_r[99] ;
wire \text_in_r[9] ;
wire \u0/_0128_ ;
wire \u0/_0129_ ;
wire \u0/_0130_ ;
wire \u0/_0131_ ;
wire \u0/_0132_ ;
wire \u0/_0133_ ;
wire \u0/_0134_ ;
wire \u0/_0135_ ;
wire \u0/_0136_ ;
wire \u0/_0137_ ;
wire \u0/_0138_ ;
wire \u0/_0139_ ;
wire \u0/_0140_ ;
wire \u0/_0141_ ;
wire \u0/_0142_ ;
wire \u0/_0143_ ;
wire \u0/_0144_ ;
wire \u0/_0145_ ;
wire \u0/_0146_ ;
wire \u0/_0147_ ;
wire \u0/_0148_ ;
wire \u0/_0149_ ;
wire \u0/_0150_ ;
wire \u0/_0151_ ;
wire \u0/_0152_ ;
wire \u0/_0153_ ;
wire \u0/_0154_ ;
wire \u0/_0155_ ;
wire \u0/_0156_ ;
wire \u0/_0157_ ;
wire \u0/_0158_ ;
wire \u0/_0159_ ;
wire \u0/_0160_ ;
wire \u0/_0161_ ;
wire \u0/_0162_ ;
wire \u0/_0163_ ;
wire \u0/_0164_ ;
wire \u0/_0165_ ;
wire \u0/_0166_ ;
wire \u0/_0167_ ;
wire \u0/_0168_ ;
wire \u0/_0169_ ;
wire \u0/_0170_ ;
wire \u0/_0171_ ;
wire \u0/_0172_ ;
wire \u0/_0173_ ;
wire \u0/_0174_ ;
wire \u0/_0175_ ;
wire \u0/_0176_ ;
wire \u0/_0177_ ;
wire \u0/_0178_ ;
wire \u0/_0179_ ;
wire \u0/_0180_ ;
wire \u0/_0181_ ;
wire \u0/_0182_ ;
wire \u0/_0183_ ;
wire \u0/_0184_ ;
wire \u0/_0185_ ;
wire \u0/_0186_ ;
wire \u0/_0187_ ;
wire \u0/_0188_ ;
wire \u0/_0189_ ;
wire \u0/_0190_ ;
wire \u0/_0191_ ;
wire \u0/_0192_ ;
wire \u0/_0193_ ;
wire \u0/_0194_ ;
wire \u0/_0195_ ;
wire \u0/_0196_ ;
wire \u0/_0197_ ;
wire \u0/_0198_ ;
wire \u0/_0199_ ;
wire \u0/_0200_ ;
wire \u0/_0201_ ;
wire \u0/_0202_ ;
wire \u0/_0203_ ;
wire \u0/_0204_ ;
wire \u0/_0205_ ;
wire \u0/_0206_ ;
wire \u0/_0207_ ;
wire \u0/_0208_ ;
wire \u0/_0209_ ;
wire \u0/_0210_ ;
wire \u0/_0211_ ;
wire \u0/_0212_ ;
wire \u0/_0213_ ;
wire \u0/_0214_ ;
wire \u0/_0215_ ;
wire \u0/_0216_ ;
wire \u0/_0217_ ;
wire \u0/_0218_ ;
wire \u0/_0219_ ;
wire \u0/_0220_ ;
wire \u0/_0221_ ;
wire \u0/_0222_ ;
wire \u0/_0223_ ;
wire \u0/_0224_ ;
wire \u0/_0225_ ;
wire \u0/_0226_ ;
wire \u0/_0227_ ;
wire \u0/_0228_ ;
wire \u0/_0229_ ;
wire \u0/_0230_ ;
wire \u0/_0231_ ;
wire \u0/_0232_ ;
wire \u0/_0233_ ;
wire \u0/_0234_ ;
wire \u0/_0235_ ;
wire \u0/_0236_ ;
wire \u0/_0237_ ;
wire \u0/_0238_ ;
wire \u0/_0239_ ;
wire \u0/_0240_ ;
wire \u0/_0241_ ;
wire \u0/_0242_ ;
wire \u0/_0243_ ;
wire \u0/_0244_ ;
wire \u0/_0245_ ;
wire \u0/_0246_ ;
wire \u0/_0247_ ;
wire \u0/_0248_ ;
wire \u0/_0249_ ;
wire \u0/_0250_ ;
wire \u0/_0251_ ;
wire \u0/_0252_ ;
wire \u0/_0253_ ;
wire \u0/_0254_ ;
wire \u0/_0255_ ;
wire \u0/_0385_ ;
wire \u0/_0386_ ;
wire \u0/_0387_ ;
wire \u0/_0388_ ;
wire \u0/_0389_ ;
wire \u0/_0390_ ;
wire \u0/_0391_ ;
wire \u0/_0392_ ;
wire \u0/_0393_ ;
wire \u0/_0394_ ;
wire \u0/_0395_ ;
wire \u0/_0396_ ;
wire \u0/_0397_ ;
wire \u0/_0398_ ;
wire \u0/_0399_ ;
wire \u0/_0400_ ;
wire \u0/_0401_ ;
wire \u0/_0402_ ;
wire \u0/_0403_ ;
wire \u0/_0404_ ;
wire \u0/_0405_ ;
wire \u0/_0406_ ;
wire \u0/_0407_ ;
wire \u0/_0408_ ;
wire \u0/_0409_ ;
wire \u0/_0410_ ;
wire \u0/_0411_ ;
wire \u0/_0412_ ;
wire \u0/_0413_ ;
wire \u0/_0414_ ;
wire \u0/_0415_ ;
wire \u0/_0416_ ;
wire \u0/_0417_ ;
wire \u0/_0418_ ;
wire \u0/_0419_ ;
wire \u0/_0420_ ;
wire \u0/_0421_ ;
wire \u0/_0422_ ;
wire \u0/_0423_ ;
wire \u0/_0424_ ;
wire \u0/_0425_ ;
wire \u0/_0426_ ;
wire \u0/_0427_ ;
wire \u0/_0428_ ;
wire \u0/_0429_ ;
wire \u0/_0430_ ;
wire \u0/_0431_ ;
wire \u0/_0432_ ;
wire \u0/_0433_ ;
wire \u0/_0434_ ;
wire \u0/_0435_ ;
wire \u0/_0436_ ;
wire \u0/_0437_ ;
wire \u0/_0438_ ;
wire \u0/_0439_ ;
wire \u0/_0440_ ;
wire \u0/_0441_ ;
wire \u0/_0442_ ;
wire \u0/_0443_ ;
wire \u0/_0444_ ;
wire \u0/_0445_ ;
wire \u0/_0446_ ;
wire \u0/_0447_ ;
wire \u0/_0448_ ;
wire \u0/_0449_ ;
wire \u0/_0450_ ;
wire \u0/_0451_ ;
wire \u0/_0452_ ;
wire \u0/_0453_ ;
wire \u0/_0454_ ;
wire \u0/_0455_ ;
wire \u0/_0456_ ;
wire \u0/_0457_ ;
wire \u0/_0458_ ;
wire \u0/_0459_ ;
wire \u0/_0460_ ;
wire \u0/_0461_ ;
wire \u0/_0462_ ;
wire \u0/_0463_ ;
wire \u0/_0464_ ;
wire \u0/_0465_ ;
wire \u0/_0466_ ;
wire \u0/_0467_ ;
wire \u0/_0468_ ;
wire \u0/_0469_ ;
wire \u0/_0470_ ;
wire \u0/_0471_ ;
wire \u0/_0472_ ;
wire \u0/_0473_ ;
wire \u0/_0474_ ;
wire \u0/_0475_ ;
wire \u0/_0476_ ;
wire \u0/_0478_ ;
wire \u0/_0479_ ;
wire \u0/_0480_ ;
wire \u0/_0481_ ;
wire \u0/_0482_ ;
wire \u0/_0483_ ;
wire \u0/_0484_ ;
wire \u0/_0485_ ;
wire \u0/_0486_ ;
wire \u0/_0487_ ;
wire \u0/_0488_ ;
wire \u0/_0489_ ;
wire \u0/_0490_ ;
wire \u0/_0491_ ;
wire \u0/_0492_ ;
wire \u0/_0493_ ;
wire \u0/_0494_ ;
wire \u0/_0495_ ;
wire \u0/_0496_ ;
wire \u0/_0497_ ;
wire \u0/_0498_ ;
wire \u0/_0499_ ;
wire \u0/_0500_ ;
wire \u0/_0501_ ;
wire \u0/_0502_ ;
wire \u0/_0503_ ;
wire \u0/_0504_ ;
wire \u0/_0505_ ;
wire \u0/_0506_ ;
wire \u0/_0507_ ;
wire \u0/_0508_ ;
wire \u0/_0509_ ;
wire \u0/_0510_ ;
wire \u0/_0511_ ;
wire \u0/_0512_ ;
wire \u0/_0513_ ;
wire \u0/_0514_ ;
wire \u0/_0515_ ;
wire \u0/_0516_ ;
wire \u0/_0517_ ;
wire \u0/_0518_ ;
wire \u0/_0519_ ;
wire \u0/_0520_ ;
wire \u0/_0521_ ;
wire \u0/_0522_ ;
wire \u0/_0523_ ;
wire \u0/_0524_ ;
wire \u0/_0525_ ;
wire \u0/_0526_ ;
wire \u0/_0527_ ;
wire \u0/_0528_ ;
wire \u0/_0529_ ;
wire \u0/_0530_ ;
wire \u0/_0531_ ;
wire \u0/_0532_ ;
wire \u0/_0533_ ;
wire \u0/_0534_ ;
wire \u0/_0535_ ;
wire \u0/_0536_ ;
wire \u0/_0537_ ;
wire \u0/_0538_ ;
wire \u0/_0539_ ;
wire \u0/_0540_ ;
wire \u0/_0541_ ;
wire \u0/_0542_ ;
wire \u0/_0543_ ;
wire \u0/_0544_ ;
wire \u0/_0545_ ;
wire \u0/_0546_ ;
wire \u0/_0547_ ;
wire \u0/_0548_ ;
wire \u0/_0549_ ;
wire \u0/_0550_ ;
wire \u0/_0551_ ;
wire \u0/_0552_ ;
wire \u0/_0553_ ;
wire \u0/_0554_ ;
wire \u0/_0555_ ;
wire \u0/_0556_ ;
wire \u0/_0557_ ;
wire \u0/_0558_ ;
wire \u0/_0559_ ;
wire \u0/_0560_ ;
wire \u0/_0561_ ;
wire \u0/_0562_ ;
wire \u0/_0563_ ;
wire \u0/_0564_ ;
wire \u0/_0565_ ;
wire \u0/_0566_ ;
wire \u0/_0567_ ;
wire \u0/_0568_ ;
wire \u0/_0569_ ;
wire \u0/_0570_ ;
wire \u0/_0571_ ;
wire \u0/_0572_ ;
wire \u0/_0573_ ;
wire \u0/_0574_ ;
wire \u0/_0576_ ;
wire \u0/_0577_ ;
wire \u0/_0578_ ;
wire \u0/_0579_ ;
wire \u0/_0580_ ;
wire \u0/_0581_ ;
wire \u0/_0582_ ;
wire \u0/_0583_ ;
wire \u0/_0584_ ;
wire \u0/_0585_ ;
wire \u0/_0586_ ;
wire \u0/_0587_ ;
wire \u0/_0588_ ;
wire \u0/_0589_ ;
wire \u0/_0590_ ;
wire \u0/_0591_ ;
wire \u0/_0592_ ;
wire \u0/_0593_ ;
wire \u0/_0594_ ;
wire \u0/_0595_ ;
wire \u0/_0596_ ;
wire \u0/_0597_ ;
wire \u0/_0598_ ;
wire \u0/_0599_ ;
wire \u0/_0600_ ;
wire \u0/_0601_ ;
wire \u0/_0602_ ;
wire \u0/_0603_ ;
wire \u0/_0604_ ;
wire \u0/_0605_ ;
wire \u0/_0606_ ;
wire \u0/_0607_ ;
wire \u0/_0608_ ;
wire \u0/_0609_ ;
wire \u0/_0610_ ;
wire \u0/_0611_ ;
wire \u0/_0612_ ;
wire \u0/_0613_ ;
wire \u0/_0614_ ;
wire \u0/_0615_ ;
wire \u0/_0616_ ;
wire \u0/_0617_ ;
wire \u0/_0618_ ;
wire \u0/_0619_ ;
wire \u0/_0620_ ;
wire \u0/_0621_ ;
wire \u0/_0622_ ;
wire \u0/_0623_ ;
wire \u0/_0624_ ;
wire \u0/_0625_ ;
wire \u0/_0626_ ;
wire \u0/_0627_ ;
wire \u0/_0628_ ;
wire \u0/_0629_ ;
wire \u0/_0630_ ;
wire \u0/_0631_ ;
wire \u0/_0632_ ;
wire \u0/_0633_ ;
wire \u0/_0634_ ;
wire \u0/_0635_ ;
wire \u0/_0636_ ;
wire \u0/_0637_ ;
wire \u0/_0638_ ;
wire \u0/_0639_ ;
wire \u0/_0640_ ;
wire \u0/_0641_ ;
wire \u0/_0642_ ;
wire \u0/_0643_ ;
wire \u0/_0644_ ;
wire \u0/_0645_ ;
wire \u0/_0646_ ;
wire \u0/_0647_ ;
wire \u0/_0648_ ;
wire \u0/_0649_ ;
wire \u0/_0650_ ;
wire \u0/_0651_ ;
wire \u0/_0652_ ;
wire \u0/_0653_ ;
wire \u0/_0654_ ;
wire \u0/_0655_ ;
wire \u0/_0656_ ;
wire \u0/_0657_ ;
wire \u0/_0842_ ;
wire \u0/r0/_036_ ;
wire \u0/r0/_037_ ;
wire \u0/r0/_038_ ;
wire \u0/r0/_039_ ;
wire \u0/r0/_040_ ;
wire \u0/r0/_041_ ;
wire \u0/r0/_042_ ;
wire \u0/r0/_043_ ;
wire \u0/r0/_044_ ;
wire \u0/r0/_045_ ;
wire \u0/r0/_046_ ;
wire \u0/r0/_047_ ;
wire \u0/r0/_049_ ;
wire \u0/r0/_050_ ;
wire \u0/r0/_051_ ;
wire \u0/r0/_052_ ;
wire \u0/r0/_053_ ;
wire \u0/r0/_054_ ;
wire \u0/r0/_055_ ;
wire \u0/r0/_056_ ;
wire \u0/r0/_057_ ;
wire \u0/r0/_058_ ;
wire \u0/r0/_059_ ;
wire \u0/r0/_060_ ;
wire \u0/r0/_061_ ;
wire \u0/r0/_062_ ;
wire \u0/r0/_063_ ;
wire \u0/r0/_064_ ;
wire \u0/r0/_065_ ;
wire \u0/r0/_066_ ;
wire \u0/r0/rcnt[0] ;
wire \u0/r0/rcnt[1] ;
wire \u0/r0/rcnt[2] ;
wire \u0/r0/rcnt[3] ;
wire \u0/rcon[0] ;
wire \u0/rcon[10] ;
wire \u0/rcon[11] ;
wire \u0/rcon[12] ;
wire \u0/rcon[13] ;
wire \u0/rcon[14] ;
wire \u0/rcon[15] ;
wire \u0/rcon[16] ;
wire \u0/rcon[17] ;
wire \u0/rcon[18] ;
wire \u0/rcon[19] ;
wire \u0/rcon[1] ;
wire \u0/rcon[20] ;
wire \u0/rcon[21] ;
wire \u0/rcon[22] ;
wire \u0/rcon[23] ;
wire \u0/rcon[24] ;
wire \u0/rcon[25] ;
wire \u0/rcon[26] ;
wire \u0/rcon[27] ;
wire \u0/rcon[28] ;
wire \u0/rcon[29] ;
wire \u0/rcon[2] ;
wire \u0/rcon[30] ;
wire \u0/rcon[31] ;
wire \u0/rcon[3] ;
wire \u0/rcon[4] ;
wire \u0/rcon[5] ;
wire \u0/rcon[6] ;
wire \u0/rcon[7] ;
wire \u0/rcon[8] ;
wire \u0/rcon[9] ;
wire \u0/u0/_0001_ ;
wire \u0/u0/_0008_ ;
wire \u0/u0/_0009_ ;
wire \u0/u0/_0010_ ;
wire \u0/u0/_0011_ ;
wire \u0/u0/_0012_ ;
wire \u0/u0/_0013_ ;
wire \u0/u0/_0014_ ;
wire \u0/u0/_0015_ ;
wire \u0/u0/_0016_ ;
wire \u0/u0/_0017_ ;
wire \u0/u0/_0018_ ;
wire \u0/u0/_0019_ ;
wire \u0/u0/_0020_ ;
wire \u0/u0/_0022_ ;
wire \u0/u0/_0023_ ;
wire \u0/u0/_0024_ ;
wire \u0/u0/_0025_ ;
wire \u0/u0/_0026_ ;
wire \u0/u0/_0027_ ;
wire \u0/u0/_0030_ ;
wire \u0/u0/_0032_ ;
wire \u0/u0/_0033_ ;
wire \u0/u0/_0034_ ;
wire \u0/u0/_0035_ ;
wire \u0/u0/_0036_ ;
wire \u0/u0/_0037_ ;
wire \u0/u0/_0038_ ;
wire \u0/u0/_0039_ ;
wire \u0/u0/_0040_ ;
wire \u0/u0/_0041_ ;
wire \u0/u0/_0042_ ;
wire \u0/u0/_0043_ ;
wire \u0/u0/_0045_ ;
wire \u0/u0/_0046_ ;
wire \u0/u0/_0047_ ;
wire \u0/u0/_0049_ ;
wire \u0/u0/_0050_ ;
wire \u0/u0/_0051_ ;
wire \u0/u0/_0052_ ;
wire \u0/u0/_0053_ ;
wire \u0/u0/_0054_ ;
wire \u0/u0/_0056_ ;
wire \u0/u0/_0057_ ;
wire \u0/u0/_0058_ ;
wire \u0/u0/_0060_ ;
wire \u0/u0/_0061_ ;
wire \u0/u0/_0062_ ;
wire \u0/u0/_0064_ ;
wire \u0/u0/_0065_ ;
wire \u0/u0/_0066_ ;
wire \u0/u0/_0067_ ;
wire \u0/u0/_0069_ ;
wire \u0/u0/_0070_ ;
wire \u0/u0/_0072_ ;
wire \u0/u0/_0073_ ;
wire \u0/u0/_0074_ ;
wire \u0/u0/_0075_ ;
wire \u0/u0/_0076_ ;
wire \u0/u0/_0077_ ;
wire \u0/u0/_0078_ ;
wire \u0/u0/_0079_ ;
wire \u0/u0/_0081_ ;
wire \u0/u0/_0082_ ;
wire \u0/u0/_0084_ ;
wire \u0/u0/_0085_ ;
wire \u0/u0/_0086_ ;
wire \u0/u0/_0087_ ;
wire \u0/u0/_0088_ ;
wire \u0/u0/_0089_ ;
wire \u0/u0/_0090_ ;
wire \u0/u0/_0091_ ;
wire \u0/u0/_0092_ ;
wire \u0/u0/_0093_ ;
wire \u0/u0/_0094_ ;
wire \u0/u0/_0095_ ;
wire \u0/u0/_0096_ ;
wire \u0/u0/_0097_ ;
wire \u0/u0/_0098_ ;
wire \u0/u0/_0099_ ;
wire \u0/u0/_0100_ ;
wire \u0/u0/_0101_ ;
wire \u0/u0/_0102_ ;
wire \u0/u0/_0103_ ;
wire \u0/u0/_0104_ ;
wire \u0/u0/_0105_ ;
wire \u0/u0/_0106_ ;
wire \u0/u0/_0108_ ;
wire \u0/u0/_0109_ ;
wire \u0/u0/_0110_ ;
wire \u0/u0/_0111_ ;
wire \u0/u0/_0113_ ;
wire \u0/u0/_0114_ ;
wire \u0/u0/_0115_ ;
wire \u0/u0/_0116_ ;
wire \u0/u0/_0117_ ;
wire \u0/u0/_0118_ ;
wire \u0/u0/_0119_ ;
wire \u0/u0/_0120_ ;
wire \u0/u0/_0121_ ;
wire \u0/u0/_0122_ ;
wire \u0/u0/_0123_ ;
wire \u0/u0/_0124_ ;
wire \u0/u0/_0126_ ;
wire \u0/u0/_0127_ ;
wire \u0/u0/_0128_ ;
wire \u0/u0/_0129_ ;
wire \u0/u0/_0130_ ;
wire \u0/u0/_0132_ ;
wire \u0/u0/_0133_ ;
wire \u0/u0/_0134_ ;
wire \u0/u0/_0135_ ;
wire \u0/u0/_0136_ ;
wire \u0/u0/_0137_ ;
wire \u0/u0/_0139_ ;
wire \u0/u0/_0140_ ;
wire \u0/u0/_0141_ ;
wire \u0/u0/_0142_ ;
wire \u0/u0/_0144_ ;
wire \u0/u0/_0145_ ;
wire \u0/u0/_0146_ ;
wire \u0/u0/_0147_ ;
wire \u0/u0/_0148_ ;
wire \u0/u0/_0149_ ;
wire \u0/u0/_0150_ ;
wire \u0/u0/_0151_ ;
wire \u0/u0/_0153_ ;
wire \u0/u0/_0154_ ;
wire \u0/u0/_0155_ ;
wire \u0/u0/_0156_ ;
wire \u0/u0/_0157_ ;
wire \u0/u0/_0158_ ;
wire \u0/u0/_0159_ ;
wire \u0/u0/_0161_ ;
wire \u0/u0/_0162_ ;
wire \u0/u0/_0163_ ;
wire \u0/u0/_0164_ ;
wire \u0/u0/_0165_ ;
wire \u0/u0/_0166_ ;
wire \u0/u0/_0167_ ;
wire \u0/u0/_0168_ ;
wire \u0/u0/_0169_ ;
wire \u0/u0/_0170_ ;
wire \u0/u0/_0171_ ;
wire \u0/u0/_0172_ ;
wire \u0/u0/_0174_ ;
wire \u0/u0/_0175_ ;
wire \u0/u0/_0176_ ;
wire \u0/u0/_0177_ ;
wire \u0/u0/_0178_ ;
wire \u0/u0/_0179_ ;
wire \u0/u0/_0180_ ;
wire \u0/u0/_0181_ ;
wire \u0/u0/_0182_ ;
wire \u0/u0/_0183_ ;
wire \u0/u0/_0184_ ;
wire \u0/u0/_0185_ ;
wire \u0/u0/_0186_ ;
wire \u0/u0/_0187_ ;
wire \u0/u0/_0188_ ;
wire \u0/u0/_0189_ ;
wire \u0/u0/_0190_ ;
wire \u0/u0/_0191_ ;
wire \u0/u0/_0192_ ;
wire \u0/u0/_0193_ ;
wire \u0/u0/_0194_ ;
wire \u0/u0/_0195_ ;
wire \u0/u0/_0196_ ;
wire \u0/u0/_0197_ ;
wire \u0/u0/_0198_ ;
wire \u0/u0/_0199_ ;
wire \u0/u0/_0200_ ;
wire \u0/u0/_0201_ ;
wire \u0/u0/_0202_ ;
wire \u0/u0/_0203_ ;
wire \u0/u0/_0204_ ;
wire \u0/u0/_0205_ ;
wire \u0/u0/_0206_ ;
wire \u0/u0/_0207_ ;
wire \u0/u0/_0208_ ;
wire \u0/u0/_0209_ ;
wire \u0/u0/_0210_ ;
wire \u0/u0/_0211_ ;
wire \u0/u0/_0212_ ;
wire \u0/u0/_0213_ ;
wire \u0/u0/_0214_ ;
wire \u0/u0/_0215_ ;
wire \u0/u0/_0216_ ;
wire \u0/u0/_0217_ ;
wire \u0/u0/_0218_ ;
wire \u0/u0/_0219_ ;
wire \u0/u0/_0220_ ;
wire \u0/u0/_0221_ ;
wire \u0/u0/_0222_ ;
wire \u0/u0/_0223_ ;
wire \u0/u0/_0224_ ;
wire \u0/u0/_0225_ ;
wire \u0/u0/_0226_ ;
wire \u0/u0/_0227_ ;
wire \u0/u0/_0228_ ;
wire \u0/u0/_0229_ ;
wire \u0/u0/_0230_ ;
wire \u0/u0/_0231_ ;
wire \u0/u0/_0232_ ;
wire \u0/u0/_0233_ ;
wire \u0/u0/_0234_ ;
wire \u0/u0/_0235_ ;
wire \u0/u0/_0236_ ;
wire \u0/u0/_0237_ ;
wire \u0/u0/_0238_ ;
wire \u0/u0/_0239_ ;
wire \u0/u0/_0240_ ;
wire \u0/u0/_0241_ ;
wire \u0/u0/_0242_ ;
wire \u0/u0/_0243_ ;
wire \u0/u0/_0244_ ;
wire \u0/u0/_0245_ ;
wire \u0/u0/_0246_ ;
wire \u0/u0/_0247_ ;
wire \u0/u0/_0248_ ;
wire \u0/u0/_0249_ ;
wire \u0/u0/_0250_ ;
wire \u0/u0/_0251_ ;
wire \u0/u0/_0252_ ;
wire \u0/u0/_0253_ ;
wire \u0/u0/_0254_ ;
wire \u0/u0/_0255_ ;
wire \u0/u0/_0256_ ;
wire \u0/u0/_0257_ ;
wire \u0/u0/_0258_ ;
wire \u0/u0/_0259_ ;
wire \u0/u0/_0260_ ;
wire \u0/u0/_0261_ ;
wire \u0/u0/_0263_ ;
wire \u0/u0/_0264_ ;
wire \u0/u0/_0265_ ;
wire \u0/u0/_0266_ ;
wire \u0/u0/_0267_ ;
wire \u0/u0/_0268_ ;
wire \u0/u0/_0269_ ;
wire \u0/u0/_0270_ ;
wire \u0/u0/_0271_ ;
wire \u0/u0/_0272_ ;
wire \u0/u0/_0273_ ;
wire \u0/u0/_0274_ ;
wire \u0/u0/_0275_ ;
wire \u0/u0/_0276_ ;
wire \u0/u0/_0277_ ;
wire \u0/u0/_0278_ ;
wire \u0/u0/_0279_ ;
wire \u0/u0/_0281_ ;
wire \u0/u0/_0283_ ;
wire \u0/u0/_0284_ ;
wire \u0/u0/_0285_ ;
wire \u0/u0/_0286_ ;
wire \u0/u0/_0287_ ;
wire \u0/u0/_0288_ ;
wire \u0/u0/_0289_ ;
wire \u0/u0/_0290_ ;
wire \u0/u0/_0291_ ;
wire \u0/u0/_0293_ ;
wire \u0/u0/_0294_ ;
wire \u0/u0/_0295_ ;
wire \u0/u0/_0296_ ;
wire \u0/u0/_0297_ ;
wire \u0/u0/_0298_ ;
wire \u0/u0/_0299_ ;
wire \u0/u0/_0300_ ;
wire \u0/u0/_0301_ ;
wire \u0/u0/_0302_ ;
wire \u0/u0/_0303_ ;
wire \u0/u0/_0304_ ;
wire \u0/u0/_0305_ ;
wire \u0/u0/_0306_ ;
wire \u0/u0/_0307_ ;
wire \u0/u0/_0308_ ;
wire \u0/u0/_0309_ ;
wire \u0/u0/_0310_ ;
wire \u0/u0/_0311_ ;
wire \u0/u0/_0312_ ;
wire \u0/u0/_0313_ ;
wire \u0/u0/_0314_ ;
wire \u0/u0/_0315_ ;
wire \u0/u0/_0316_ ;
wire \u0/u0/_0317_ ;
wire \u0/u0/_0318_ ;
wire \u0/u0/_0319_ ;
wire \u0/u0/_0320_ ;
wire \u0/u0/_0321_ ;
wire \u0/u0/_0322_ ;
wire \u0/u0/_0323_ ;
wire \u0/u0/_0324_ ;
wire \u0/u0/_0325_ ;
wire \u0/u0/_0326_ ;
wire \u0/u0/_0327_ ;
wire \u0/u0/_0328_ ;
wire \u0/u0/_0329_ ;
wire \u0/u0/_0330_ ;
wire \u0/u0/_0331_ ;
wire \u0/u0/_0332_ ;
wire \u0/u0/_0333_ ;
wire \u0/u0/_0334_ ;
wire \u0/u0/_0335_ ;
wire \u0/u0/_0337_ ;
wire \u0/u0/_0338_ ;
wire \u0/u0/_0339_ ;
wire \u0/u0/_0340_ ;
wire \u0/u0/_0341_ ;
wire \u0/u0/_0342_ ;
wire \u0/u0/_0343_ ;
wire \u0/u0/_0344_ ;
wire \u0/u0/_0345_ ;
wire \u0/u0/_0347_ ;
wire \u0/u0/_0348_ ;
wire \u0/u0/_0349_ ;
wire \u0/u0/_0350_ ;
wire \u0/u0/_0351_ ;
wire \u0/u0/_0352_ ;
wire \u0/u0/_0353_ ;
wire \u0/u0/_0354_ ;
wire \u0/u0/_0355_ ;
wire \u0/u0/_0356_ ;
wire \u0/u0/_0357_ ;
wire \u0/u0/_0358_ ;
wire \u0/u0/_0359_ ;
wire \u0/u0/_0360_ ;
wire \u0/u0/_0361_ ;
wire \u0/u0/_0362_ ;
wire \u0/u0/_0363_ ;
wire \u0/u0/_0365_ ;
wire \u0/u0/_0366_ ;
wire \u0/u0/_0367_ ;
wire \u0/u0/_0368_ ;
wire \u0/u0/_0370_ ;
wire \u0/u0/_0371_ ;
wire \u0/u0/_0372_ ;
wire \u0/u0/_0373_ ;
wire \u0/u0/_0374_ ;
wire \u0/u0/_0375_ ;
wire \u0/u0/_0376_ ;
wire \u0/u0/_0377_ ;
wire \u0/u0/_0378_ ;
wire \u0/u0/_0379_ ;
wire \u0/u0/_0380_ ;
wire \u0/u0/_0381_ ;
wire \u0/u0/_0382_ ;
wire \u0/u0/_0383_ ;
wire \u0/u0/_0384_ ;
wire \u0/u0/_0385_ ;
wire \u0/u0/_0386_ ;
wire \u0/u0/_0387_ ;
wire \u0/u0/_0388_ ;
wire \u0/u0/_0389_ ;
wire \u0/u0/_0390_ ;
wire \u0/u0/_0391_ ;
wire \u0/u0/_0392_ ;
wire \u0/u0/_0393_ ;
wire \u0/u0/_0394_ ;
wire \u0/u0/_0395_ ;
wire \u0/u0/_0396_ ;
wire \u0/u0/_0397_ ;
wire \u0/u0/_0398_ ;
wire \u0/u0/_0399_ ;
wire \u0/u0/_0400_ ;
wire \u0/u0/_0401_ ;
wire \u0/u0/_0402_ ;
wire \u0/u0/_0403_ ;
wire \u0/u0/_0404_ ;
wire \u0/u0/_0405_ ;
wire \u0/u0/_0406_ ;
wire \u0/u0/_0407_ ;
wire \u0/u0/_0408_ ;
wire \u0/u0/_0409_ ;
wire \u0/u0/_0410_ ;
wire \u0/u0/_0411_ ;
wire \u0/u0/_0412_ ;
wire \u0/u0/_0413_ ;
wire \u0/u0/_0414_ ;
wire \u0/u0/_0415_ ;
wire \u0/u0/_0416_ ;
wire \u0/u0/_0417_ ;
wire \u0/u0/_0418_ ;
wire \u0/u0/_0419_ ;
wire \u0/u0/_0420_ ;
wire \u0/u0/_0421_ ;
wire \u0/u0/_0422_ ;
wire \u0/u0/_0423_ ;
wire \u0/u0/_0424_ ;
wire \u0/u0/_0425_ ;
wire \u0/u0/_0426_ ;
wire \u0/u0/_0427_ ;
wire \u0/u0/_0428_ ;
wire \u0/u0/_0429_ ;
wire \u0/u0/_0430_ ;
wire \u0/u0/_0431_ ;
wire \u0/u0/_0432_ ;
wire \u0/u0/_0433_ ;
wire \u0/u0/_0434_ ;
wire \u0/u0/_0435_ ;
wire \u0/u0/_0436_ ;
wire \u0/u0/_0437_ ;
wire \u0/u0/_0438_ ;
wire \u0/u0/_0439_ ;
wire \u0/u0/_0440_ ;
wire \u0/u0/_0441_ ;
wire \u0/u0/_0442_ ;
wire \u0/u0/_0443_ ;
wire \u0/u0/_0444_ ;
wire \u0/u0/_0446_ ;
wire \u0/u0/_0447_ ;
wire \u0/u0/_0448_ ;
wire \u0/u0/_0449_ ;
wire \u0/u0/_0450_ ;
wire \u0/u0/_0451_ ;
wire \u0/u0/_0452_ ;
wire \u0/u0/_0453_ ;
wire \u0/u0/_0454_ ;
wire \u0/u0/_0455_ ;
wire \u0/u0/_0457_ ;
wire \u0/u0/_0458_ ;
wire \u0/u0/_0459_ ;
wire \u0/u0/_0460_ ;
wire \u0/u0/_0461_ ;
wire \u0/u0/_0462_ ;
wire \u0/u0/_0463_ ;
wire \u0/u0/_0464_ ;
wire \u0/u0/_0465_ ;
wire \u0/u0/_0466_ ;
wire \u0/u0/_0467_ ;
wire \u0/u0/_0468_ ;
wire \u0/u0/_0469_ ;
wire \u0/u0/_0470_ ;
wire \u0/u0/_0471_ ;
wire \u0/u0/_0472_ ;
wire \u0/u0/_0473_ ;
wire \u0/u0/_0474_ ;
wire \u0/u0/_0475_ ;
wire \u0/u0/_0476_ ;
wire \u0/u0/_0477_ ;
wire \u0/u0/_0478_ ;
wire \u0/u0/_0479_ ;
wire \u0/u0/_0480_ ;
wire \u0/u0/_0481_ ;
wire \u0/u0/_0482_ ;
wire \u0/u0/_0483_ ;
wire \u0/u0/_0484_ ;
wire \u0/u0/_0485_ ;
wire \u0/u0/_0486_ ;
wire \u0/u0/_0487_ ;
wire \u0/u0/_0488_ ;
wire \u0/u0/_0490_ ;
wire \u0/u0/_0491_ ;
wire \u0/u0/_0492_ ;
wire \u0/u0/_0493_ ;
wire \u0/u0/_0494_ ;
wire \u0/u0/_0495_ ;
wire \u0/u0/_0496_ ;
wire \u0/u0/_0497_ ;
wire \u0/u0/_0498_ ;
wire \u0/u0/_0500_ ;
wire \u0/u0/_0501_ ;
wire \u0/u0/_0502_ ;
wire \u0/u0/_0503_ ;
wire \u0/u0/_0504_ ;
wire \u0/u0/_0505_ ;
wire \u0/u0/_0506_ ;
wire \u0/u0/_0507_ ;
wire \u0/u0/_0508_ ;
wire \u0/u0/_0509_ ;
wire \u0/u0/_0510_ ;
wire \u0/u0/_0511_ ;
wire \u0/u0/_0512_ ;
wire \u0/u0/_0513_ ;
wire \u0/u0/_0514_ ;
wire \u0/u0/_0515_ ;
wire \u0/u0/_0516_ ;
wire \u0/u0/_0517_ ;
wire \u0/u0/_0518_ ;
wire \u0/u0/_0519_ ;
wire \u0/u0/_0520_ ;
wire \u0/u0/_0521_ ;
wire \u0/u0/_0522_ ;
wire \u0/u0/_0523_ ;
wire \u0/u0/_0524_ ;
wire \u0/u0/_0525_ ;
wire \u0/u0/_0526_ ;
wire \u0/u0/_0527_ ;
wire \u0/u0/_0528_ ;
wire \u0/u0/_0529_ ;
wire \u0/u0/_0530_ ;
wire \u0/u0/_0531_ ;
wire \u0/u0/_0532_ ;
wire \u0/u0/_0533_ ;
wire \u0/u0/_0534_ ;
wire \u0/u0/_0535_ ;
wire \u0/u0/_0536_ ;
wire \u0/u0/_0537_ ;
wire \u0/u0/_0538_ ;
wire \u0/u0/_0539_ ;
wire \u0/u0/_0540_ ;
wire \u0/u0/_0541_ ;
wire \u0/u0/_0542_ ;
wire \u0/u0/_0543_ ;
wire \u0/u0/_0544_ ;
wire \u0/u0/_0545_ ;
wire \u0/u0/_0546_ ;
wire \u0/u0/_0547_ ;
wire \u0/u0/_0548_ ;
wire \u0/u0/_0549_ ;
wire \u0/u0/_0550_ ;
wire \u0/u0/_0551_ ;
wire \u0/u0/_0552_ ;
wire \u0/u0/_0553_ ;
wire \u0/u0/_0554_ ;
wire \u0/u0/_0555_ ;
wire \u0/u0/_0556_ ;
wire \u0/u0/_0557_ ;
wire \u0/u0/_0558_ ;
wire \u0/u0/_0559_ ;
wire \u0/u0/_0560_ ;
wire \u0/u0/_0561_ ;
wire \u0/u0/_0562_ ;
wire \u0/u0/_0563_ ;
wire \u0/u0/_0565_ ;
wire \u0/u0/_0566_ ;
wire \u0/u0/_0567_ ;
wire \u0/u0/_0568_ ;
wire \u0/u0/_0569_ ;
wire \u0/u0/_0570_ ;
wire \u0/u0/_0571_ ;
wire \u0/u0/_0572_ ;
wire \u0/u0/_0573_ ;
wire \u0/u0/_0574_ ;
wire \u0/u0/_0575_ ;
wire \u0/u0/_0576_ ;
wire \u0/u0/_0577_ ;
wire \u0/u0/_0578_ ;
wire \u0/u0/_0579_ ;
wire \u0/u0/_0580_ ;
wire \u0/u0/_0581_ ;
wire \u0/u0/_0582_ ;
wire \u0/u0/_0583_ ;
wire \u0/u0/_0584_ ;
wire \u0/u0/_0585_ ;
wire \u0/u0/_0586_ ;
wire \u0/u0/_0587_ ;
wire \u0/u0/_0588_ ;
wire \u0/u0/_0589_ ;
wire \u0/u0/_0590_ ;
wire \u0/u0/_0591_ ;
wire \u0/u0/_0592_ ;
wire \u0/u0/_0593_ ;
wire \u0/u0/_0594_ ;
wire \u0/u0/_0595_ ;
wire \u0/u0/_0596_ ;
wire \u0/u0/_0598_ ;
wire \u0/u0/_0599_ ;
wire \u0/u0/_0600_ ;
wire \u0/u0/_0601_ ;
wire \u0/u0/_0602_ ;
wire \u0/u0/_0603_ ;
wire \u0/u0/_0604_ ;
wire \u0/u0/_0605_ ;
wire \u0/u0/_0606_ ;
wire \u0/u0/_0607_ ;
wire \u0/u0/_0608_ ;
wire \u0/u0/_0609_ ;
wire \u0/u0/_0610_ ;
wire \u0/u0/_0611_ ;
wire \u0/u0/_0612_ ;
wire \u0/u0/_0613_ ;
wire \u0/u0/_0614_ ;
wire \u0/u0/_0615_ ;
wire \u0/u0/_0616_ ;
wire \u0/u0/_0617_ ;
wire \u0/u0/_0618_ ;
wire \u0/u0/_0619_ ;
wire \u0/u0/_0620_ ;
wire \u0/u0/_0621_ ;
wire \u0/u0/_0622_ ;
wire \u0/u0/_0623_ ;
wire \u0/u0/_0624_ ;
wire \u0/u0/_0625_ ;
wire \u0/u0/_0626_ ;
wire \u0/u0/_0627_ ;
wire \u0/u0/_0628_ ;
wire \u0/u0/_0629_ ;
wire \u0/u0/_0630_ ;
wire \u0/u0/_0631_ ;
wire \u0/u0/_0632_ ;
wire \u0/u0/_0633_ ;
wire \u0/u0/_0634_ ;
wire \u0/u0/_0635_ ;
wire \u0/u0/_0636_ ;
wire \u0/u0/_0637_ ;
wire \u0/u0/_0638_ ;
wire \u0/u0/_0639_ ;
wire \u0/u0/_0640_ ;
wire \u0/u0/_0641_ ;
wire \u0/u0/_0642_ ;
wire \u0/u0/_0643_ ;
wire \u0/u0/_0644_ ;
wire \u0/u0/_0645_ ;
wire \u0/u0/_0646_ ;
wire \u0/u0/_0647_ ;
wire \u0/u0/_0648_ ;
wire \u0/u0/_0649_ ;
wire \u0/u0/_0650_ ;
wire \u0/u0/_0651_ ;
wire \u0/u0/_0652_ ;
wire \u0/u0/_0653_ ;
wire \u0/u0/_0654_ ;
wire \u0/u0/_0655_ ;
wire \u0/u0/_0656_ ;
wire \u0/u0/_0657_ ;
wire \u0/u0/_0658_ ;
wire \u0/u0/_0659_ ;
wire \u0/u0/_0660_ ;
wire \u0/u0/_0661_ ;
wire \u0/u0/_0662_ ;
wire \u0/u0/_0663_ ;
wire \u0/u0/_0664_ ;
wire \u0/u0/_0665_ ;
wire \u0/u0/_0666_ ;
wire \u0/u0/_0667_ ;
wire \u0/u0/_0668_ ;
wire \u0/u0/_0669_ ;
wire \u0/u0/_0670_ ;
wire \u0/u0/_0671_ ;
wire \u0/u0/_0672_ ;
wire \u0/u0/_0673_ ;
wire \u0/u0/_0674_ ;
wire \u0/u0/_0675_ ;
wire \u0/u0/_0676_ ;
wire \u0/u0/_0677_ ;
wire \u0/u0/_0678_ ;
wire \u0/u0/_0679_ ;
wire \u0/u0/_0680_ ;
wire \u0/u0/_0681_ ;
wire \u0/u0/_0682_ ;
wire \u0/u0/_0683_ ;
wire \u0/u0/_0684_ ;
wire \u0/u0/_0685_ ;
wire \u0/u0/_0686_ ;
wire \u0/u0/_0687_ ;
wire \u0/u0/_0688_ ;
wire \u0/u0/_0689_ ;
wire \u0/u0/_0690_ ;
wire \u0/u0/_0691_ ;
wire \u0/u0/_0692_ ;
wire \u0/u0/_0693_ ;
wire \u0/u0/_0694_ ;
wire \u0/u0/_0695_ ;
wire \u0/u0/_0696_ ;
wire \u0/u0/_0697_ ;
wire \u0/u0/_0698_ ;
wire \u0/u0/_0699_ ;
wire \u0/u0/_0700_ ;
wire \u0/u0/_0701_ ;
wire \u0/u0/_0702_ ;
wire \u0/u0/_0703_ ;
wire \u0/u0/_0704_ ;
wire \u0/u0/_0705_ ;
wire \u0/u0/_0706_ ;
wire \u0/u0/_0707_ ;
wire \u0/u0/_0708_ ;
wire \u0/u0/_0709_ ;
wire \u0/u0/_0710_ ;
wire \u0/u0/_0711_ ;
wire \u0/u0/_0712_ ;
wire \u0/u0/_0713_ ;
wire \u0/u0/_0714_ ;
wire \u0/u0/_0715_ ;
wire \u0/u0/_0717_ ;
wire \u0/u0/_0718_ ;
wire \u0/u0/_0719_ ;
wire \u0/u0/_0720_ ;
wire \u0/u0/_0721_ ;
wire \u0/u0/_0722_ ;
wire \u0/u0/_0723_ ;
wire \u0/u0/_0724_ ;
wire \u0/u0/_0725_ ;
wire \u0/u0/_0726_ ;
wire \u0/u0/_0727_ ;
wire \u0/u0/_0728_ ;
wire \u0/u0/_0729_ ;
wire \u0/u0/_0730_ ;
wire \u0/u0/_0731_ ;
wire \u0/u0/_0732_ ;
wire \u0/u0/_0733_ ;
wire \u0/u0/_0734_ ;
wire \u0/u0/_0735_ ;
wire \u0/u0/_0736_ ;
wire \u0/u0/_0738_ ;
wire \u0/u0/_0739_ ;
wire \u0/u0/_0740_ ;
wire \u0/u0/_0741_ ;
wire \u0/u0/_0742_ ;
wire \u0/u0/_0743_ ;
wire \u0/u0/_0744_ ;
wire \u0/u0/_0745_ ;
wire \u0/u0/_0746_ ;
wire \u0/u0/_0747_ ;
wire \u0/u0/_0748_ ;
wire \u0/u0/_0749_ ;
wire \u0/u0/_0750_ ;
wire \u0/u0/_0752_ ;
wire \u0/u1/_0008_ ;
wire \u0/u1/_0009_ ;
wire \u0/u1/_0010_ ;
wire \u0/u1/_0011_ ;
wire \u0/u1/_0012_ ;
wire \u0/u1/_0013_ ;
wire \u0/u1/_0014_ ;
wire \u0/u1/_0015_ ;
wire \u0/u1/_0016_ ;
wire \u0/u1/_0017_ ;
wire \u0/u1/_0019_ ;
wire \u0/u1/_0020_ ;
wire \u0/u1/_0022_ ;
wire \u0/u1/_0024_ ;
wire \u0/u1/_0025_ ;
wire \u0/u1/_0026_ ;
wire \u0/u1/_0027_ ;
wire \u0/u1/_0029_ ;
wire \u0/u1/_0030_ ;
wire \u0/u1/_0032_ ;
wire \u0/u1/_0033_ ;
wire \u0/u1/_0034_ ;
wire \u0/u1/_0035_ ;
wire \u0/u1/_0037_ ;
wire \u0/u1/_0038_ ;
wire \u0/u1/_0039_ ;
wire \u0/u1/_0040_ ;
wire \u0/u1/_0041_ ;
wire \u0/u1/_0042_ ;
wire \u0/u1/_0043_ ;
wire \u0/u1/_0045_ ;
wire \u0/u1/_0046_ ;
wire \u0/u1/_0047_ ;
wire \u0/u1/_0049_ ;
wire \u0/u1/_0050_ ;
wire \u0/u1/_0051_ ;
wire \u0/u1/_0052_ ;
wire \u0/u1/_0053_ ;
wire \u0/u1/_0054_ ;
wire \u0/u1/_0056_ ;
wire \u0/u1/_0057_ ;
wire \u0/u1/_0058_ ;
wire \u0/u1/_0060_ ;
wire \u0/u1/_0061_ ;
wire \u0/u1/_0062_ ;
wire \u0/u1/_0064_ ;
wire \u0/u1/_0065_ ;
wire \u0/u1/_0066_ ;
wire \u0/u1/_0067_ ;
wire \u0/u1/_0069_ ;
wire \u0/u1/_0070_ ;
wire \u0/u1/_0072_ ;
wire \u0/u1/_0073_ ;
wire \u0/u1/_0074_ ;
wire \u0/u1/_0075_ ;
wire \u0/u1/_0076_ ;
wire \u0/u1/_0077_ ;
wire \u0/u1/_0078_ ;
wire \u0/u1/_0079_ ;
wire \u0/u1/_0081_ ;
wire \u0/u1/_0082_ ;
wire \u0/u1/_0084_ ;
wire \u0/u1/_0085_ ;
wire \u0/u1/_0086_ ;
wire \u0/u1/_0087_ ;
wire \u0/u1/_0088_ ;
wire \u0/u1/_0089_ ;
wire \u0/u1/_0090_ ;
wire \u0/u1/_0091_ ;
wire \u0/u1/_0092_ ;
wire \u0/u1/_0093_ ;
wire \u0/u1/_0094_ ;
wire \u0/u1/_0095_ ;
wire \u0/u1/_0096_ ;
wire \u0/u1/_0097_ ;
wire \u0/u1/_0098_ ;
wire \u0/u1/_0099_ ;
wire \u0/u1/_0100_ ;
wire \u0/u1/_0101_ ;
wire \u0/u1/_0102_ ;
wire \u0/u1/_0103_ ;
wire \u0/u1/_0104_ ;
wire \u0/u1/_0105_ ;
wire \u0/u1/_0106_ ;
wire \u0/u1/_0108_ ;
wire \u0/u1/_0109_ ;
wire \u0/u1/_0110_ ;
wire \u0/u1/_0111_ ;
wire \u0/u1/_0113_ ;
wire \u0/u1/_0114_ ;
wire \u0/u1/_0115_ ;
wire \u0/u1/_0116_ ;
wire \u0/u1/_0117_ ;
wire \u0/u1/_0118_ ;
wire \u0/u1/_0119_ ;
wire \u0/u1/_0120_ ;
wire \u0/u1/_0121_ ;
wire \u0/u1/_0122_ ;
wire \u0/u1/_0123_ ;
wire \u0/u1/_0124_ ;
wire \u0/u1/_0126_ ;
wire \u0/u1/_0127_ ;
wire \u0/u1/_0128_ ;
wire \u0/u1/_0129_ ;
wire \u0/u1/_0130_ ;
wire \u0/u1/_0132_ ;
wire \u0/u1/_0133_ ;
wire \u0/u1/_0135_ ;
wire \u0/u1/_0136_ ;
wire \u0/u1/_0137_ ;
wire \u0/u1/_0139_ ;
wire \u0/u1/_0140_ ;
wire \u0/u1/_0141_ ;
wire \u0/u1/_0142_ ;
wire \u0/u1/_0144_ ;
wire \u0/u1/_0145_ ;
wire \u0/u1/_0146_ ;
wire \u0/u1/_0147_ ;
wire \u0/u1/_0148_ ;
wire \u0/u1/_0149_ ;
wire \u0/u1/_0150_ ;
wire \u0/u1/_0151_ ;
wire \u0/u1/_0153_ ;
wire \u0/u1/_0154_ ;
wire \u0/u1/_0155_ ;
wire \u0/u1/_0156_ ;
wire \u0/u1/_0157_ ;
wire \u0/u1/_0158_ ;
wire \u0/u1/_0159_ ;
wire \u0/u1/_0161_ ;
wire \u0/u1/_0162_ ;
wire \u0/u1/_0163_ ;
wire \u0/u1/_0164_ ;
wire \u0/u1/_0165_ ;
wire \u0/u1/_0166_ ;
wire \u0/u1/_0167_ ;
wire \u0/u1/_0168_ ;
wire \u0/u1/_0169_ ;
wire \u0/u1/_0170_ ;
wire \u0/u1/_0171_ ;
wire \u0/u1/_0172_ ;
wire \u0/u1/_0174_ ;
wire \u0/u1/_0175_ ;
wire \u0/u1/_0176_ ;
wire \u0/u1/_0177_ ;
wire \u0/u1/_0178_ ;
wire \u0/u1/_0179_ ;
wire \u0/u1/_0180_ ;
wire \u0/u1/_0181_ ;
wire \u0/u1/_0182_ ;
wire \u0/u1/_0183_ ;
wire \u0/u1/_0184_ ;
wire \u0/u1/_0185_ ;
wire \u0/u1/_0186_ ;
wire \u0/u1/_0187_ ;
wire \u0/u1/_0188_ ;
wire \u0/u1/_0189_ ;
wire \u0/u1/_0190_ ;
wire \u0/u1/_0191_ ;
wire \u0/u1/_0192_ ;
wire \u0/u1/_0193_ ;
wire \u0/u1/_0194_ ;
wire \u0/u1/_0195_ ;
wire \u0/u1/_0196_ ;
wire \u0/u1/_0197_ ;
wire \u0/u1/_0198_ ;
wire \u0/u1/_0199_ ;
wire \u0/u1/_0200_ ;
wire \u0/u1/_0201_ ;
wire \u0/u1/_0202_ ;
wire \u0/u1/_0203_ ;
wire \u0/u1/_0204_ ;
wire \u0/u1/_0205_ ;
wire \u0/u1/_0206_ ;
wire \u0/u1/_0207_ ;
wire \u0/u1/_0208_ ;
wire \u0/u1/_0209_ ;
wire \u0/u1/_0210_ ;
wire \u0/u1/_0211_ ;
wire \u0/u1/_0212_ ;
wire \u0/u1/_0213_ ;
wire \u0/u1/_0214_ ;
wire \u0/u1/_0215_ ;
wire \u0/u1/_0216_ ;
wire \u0/u1/_0217_ ;
wire \u0/u1/_0218_ ;
wire \u0/u1/_0219_ ;
wire \u0/u1/_0220_ ;
wire \u0/u1/_0221_ ;
wire \u0/u1/_0222_ ;
wire \u0/u1/_0223_ ;
wire \u0/u1/_0224_ ;
wire \u0/u1/_0225_ ;
wire \u0/u1/_0226_ ;
wire \u0/u1/_0227_ ;
wire \u0/u1/_0228_ ;
wire \u0/u1/_0229_ ;
wire \u0/u1/_0230_ ;
wire \u0/u1/_0231_ ;
wire \u0/u1/_0232_ ;
wire \u0/u1/_0233_ ;
wire \u0/u1/_0234_ ;
wire \u0/u1/_0235_ ;
wire \u0/u1/_0236_ ;
wire \u0/u1/_0237_ ;
wire \u0/u1/_0238_ ;
wire \u0/u1/_0239_ ;
wire \u0/u1/_0240_ ;
wire \u0/u1/_0241_ ;
wire \u0/u1/_0242_ ;
wire \u0/u1/_0243_ ;
wire \u0/u1/_0244_ ;
wire \u0/u1/_0245_ ;
wire \u0/u1/_0246_ ;
wire \u0/u1/_0248_ ;
wire \u0/u1/_0249_ ;
wire \u0/u1/_0250_ ;
wire \u0/u1/_0251_ ;
wire \u0/u1/_0252_ ;
wire \u0/u1/_0253_ ;
wire \u0/u1/_0254_ ;
wire \u0/u1/_0255_ ;
wire \u0/u1/_0256_ ;
wire \u0/u1/_0257_ ;
wire \u0/u1/_0258_ ;
wire \u0/u1/_0259_ ;
wire \u0/u1/_0260_ ;
wire \u0/u1/_0261_ ;
wire \u0/u1/_0263_ ;
wire \u0/u1/_0264_ ;
wire \u0/u1/_0265_ ;
wire \u0/u1/_0266_ ;
wire \u0/u1/_0267_ ;
wire \u0/u1/_0268_ ;
wire \u0/u1/_0269_ ;
wire \u0/u1/_0270_ ;
wire \u0/u1/_0271_ ;
wire \u0/u1/_0272_ ;
wire \u0/u1/_0273_ ;
wire \u0/u1/_0274_ ;
wire \u0/u1/_0275_ ;
wire \u0/u1/_0276_ ;
wire \u0/u1/_0277_ ;
wire \u0/u1/_0278_ ;
wire \u0/u1/_0279_ ;
wire \u0/u1/_0281_ ;
wire \u0/u1/_0283_ ;
wire \u0/u1/_0284_ ;
wire \u0/u1/_0285_ ;
wire \u0/u1/_0286_ ;
wire \u0/u1/_0287_ ;
wire \u0/u1/_0288_ ;
wire \u0/u1/_0289_ ;
wire \u0/u1/_0290_ ;
wire \u0/u1/_0291_ ;
wire \u0/u1/_0293_ ;
wire \u0/u1/_0294_ ;
wire \u0/u1/_0295_ ;
wire \u0/u1/_0296_ ;
wire \u0/u1/_0297_ ;
wire \u0/u1/_0298_ ;
wire \u0/u1/_0299_ ;
wire \u0/u1/_0300_ ;
wire \u0/u1/_0301_ ;
wire \u0/u1/_0302_ ;
wire \u0/u1/_0303_ ;
wire \u0/u1/_0304_ ;
wire \u0/u1/_0305_ ;
wire \u0/u1/_0306_ ;
wire \u0/u1/_0307_ ;
wire \u0/u1/_0308_ ;
wire \u0/u1/_0309_ ;
wire \u0/u1/_0310_ ;
wire \u0/u1/_0311_ ;
wire \u0/u1/_0312_ ;
wire \u0/u1/_0313_ ;
wire \u0/u1/_0314_ ;
wire \u0/u1/_0315_ ;
wire \u0/u1/_0316_ ;
wire \u0/u1/_0317_ ;
wire \u0/u1/_0318_ ;
wire \u0/u1/_0319_ ;
wire \u0/u1/_0320_ ;
wire \u0/u1/_0321_ ;
wire \u0/u1/_0322_ ;
wire \u0/u1/_0323_ ;
wire \u0/u1/_0324_ ;
wire \u0/u1/_0325_ ;
wire \u0/u1/_0326_ ;
wire \u0/u1/_0327_ ;
wire \u0/u1/_0328_ ;
wire \u0/u1/_0329_ ;
wire \u0/u1/_0330_ ;
wire \u0/u1/_0331_ ;
wire \u0/u1/_0332_ ;
wire \u0/u1/_0333_ ;
wire \u0/u1/_0334_ ;
wire \u0/u1/_0335_ ;
wire \u0/u1/_0337_ ;
wire \u0/u1/_0338_ ;
wire \u0/u1/_0339_ ;
wire \u0/u1/_0340_ ;
wire \u0/u1/_0341_ ;
wire \u0/u1/_0342_ ;
wire \u0/u1/_0343_ ;
wire \u0/u1/_0344_ ;
wire \u0/u1/_0345_ ;
wire \u0/u1/_0347_ ;
wire \u0/u1/_0348_ ;
wire \u0/u1/_0349_ ;
wire \u0/u1/_0350_ ;
wire \u0/u1/_0351_ ;
wire \u0/u1/_0352_ ;
wire \u0/u1/_0353_ ;
wire \u0/u1/_0354_ ;
wire \u0/u1/_0355_ ;
wire \u0/u1/_0356_ ;
wire \u0/u1/_0357_ ;
wire \u0/u1/_0358_ ;
wire \u0/u1/_0359_ ;
wire \u0/u1/_0360_ ;
wire \u0/u1/_0361_ ;
wire \u0/u1/_0362_ ;
wire \u0/u1/_0363_ ;
wire \u0/u1/_0365_ ;
wire \u0/u1/_0366_ ;
wire \u0/u1/_0367_ ;
wire \u0/u1/_0368_ ;
wire \u0/u1/_0370_ ;
wire \u0/u1/_0371_ ;
wire \u0/u1/_0372_ ;
wire \u0/u1/_0373_ ;
wire \u0/u1/_0374_ ;
wire \u0/u1/_0375_ ;
wire \u0/u1/_0376_ ;
wire \u0/u1/_0377_ ;
wire \u0/u1/_0378_ ;
wire \u0/u1/_0379_ ;
wire \u0/u1/_0380_ ;
wire \u0/u1/_0381_ ;
wire \u0/u1/_0382_ ;
wire \u0/u1/_0383_ ;
wire \u0/u1/_0384_ ;
wire \u0/u1/_0385_ ;
wire \u0/u1/_0386_ ;
wire \u0/u1/_0387_ ;
wire \u0/u1/_0388_ ;
wire \u0/u1/_0389_ ;
wire \u0/u1/_0390_ ;
wire \u0/u1/_0391_ ;
wire \u0/u1/_0392_ ;
wire \u0/u1/_0393_ ;
wire \u0/u1/_0394_ ;
wire \u0/u1/_0395_ ;
wire \u0/u1/_0396_ ;
wire \u0/u1/_0397_ ;
wire \u0/u1/_0398_ ;
wire \u0/u1/_0399_ ;
wire \u0/u1/_0400_ ;
wire \u0/u1/_0401_ ;
wire \u0/u1/_0402_ ;
wire \u0/u1/_0403_ ;
wire \u0/u1/_0404_ ;
wire \u0/u1/_0405_ ;
wire \u0/u1/_0406_ ;
wire \u0/u1/_0407_ ;
wire \u0/u1/_0408_ ;
wire \u0/u1/_0409_ ;
wire \u0/u1/_0410_ ;
wire \u0/u1/_0411_ ;
wire \u0/u1/_0412_ ;
wire \u0/u1/_0413_ ;
wire \u0/u1/_0414_ ;
wire \u0/u1/_0415_ ;
wire \u0/u1/_0416_ ;
wire \u0/u1/_0417_ ;
wire \u0/u1/_0418_ ;
wire \u0/u1/_0419_ ;
wire \u0/u1/_0420_ ;
wire \u0/u1/_0421_ ;
wire \u0/u1/_0422_ ;
wire \u0/u1/_0424_ ;
wire \u0/u1/_0425_ ;
wire \u0/u1/_0426_ ;
wire \u0/u1/_0427_ ;
wire \u0/u1/_0428_ ;
wire \u0/u1/_0429_ ;
wire \u0/u1/_0430_ ;
wire \u0/u1/_0431_ ;
wire \u0/u1/_0432_ ;
wire \u0/u1/_0433_ ;
wire \u0/u1/_0434_ ;
wire \u0/u1/_0435_ ;
wire \u0/u1/_0436_ ;
wire \u0/u1/_0437_ ;
wire \u0/u1/_0438_ ;
wire \u0/u1/_0439_ ;
wire \u0/u1/_0440_ ;
wire \u0/u1/_0441_ ;
wire \u0/u1/_0442_ ;
wire \u0/u1/_0443_ ;
wire \u0/u1/_0444_ ;
wire \u0/u1/_0446_ ;
wire \u0/u1/_0447_ ;
wire \u0/u1/_0448_ ;
wire \u0/u1/_0449_ ;
wire \u0/u1/_0450_ ;
wire \u0/u1/_0451_ ;
wire \u0/u1/_0452_ ;
wire \u0/u1/_0453_ ;
wire \u0/u1/_0454_ ;
wire \u0/u1/_0455_ ;
wire \u0/u1/_0456_ ;
wire \u0/u1/_0457_ ;
wire \u0/u1/_0458_ ;
wire \u0/u1/_0459_ ;
wire \u0/u1/_0460_ ;
wire \u0/u1/_0461_ ;
wire \u0/u1/_0462_ ;
wire \u0/u1/_0463_ ;
wire \u0/u1/_0464_ ;
wire \u0/u1/_0465_ ;
wire \u0/u1/_0466_ ;
wire \u0/u1/_0467_ ;
wire \u0/u1/_0468_ ;
wire \u0/u1/_0469_ ;
wire \u0/u1/_0470_ ;
wire \u0/u1/_0471_ ;
wire \u0/u1/_0472_ ;
wire \u0/u1/_0473_ ;
wire \u0/u1/_0474_ ;
wire \u0/u1/_0475_ ;
wire \u0/u1/_0476_ ;
wire \u0/u1/_0477_ ;
wire \u0/u1/_0478_ ;
wire \u0/u1/_0479_ ;
wire \u0/u1/_0480_ ;
wire \u0/u1/_0481_ ;
wire \u0/u1/_0482_ ;
wire \u0/u1/_0483_ ;
wire \u0/u1/_0484_ ;
wire \u0/u1/_0485_ ;
wire \u0/u1/_0486_ ;
wire \u0/u1/_0487_ ;
wire \u0/u1/_0488_ ;
wire \u0/u1/_0490_ ;
wire \u0/u1/_0491_ ;
wire \u0/u1/_0492_ ;
wire \u0/u1/_0493_ ;
wire \u0/u1/_0494_ ;
wire \u0/u1/_0495_ ;
wire \u0/u1/_0496_ ;
wire \u0/u1/_0497_ ;
wire \u0/u1/_0498_ ;
wire \u0/u1/_0500_ ;
wire \u0/u1/_0501_ ;
wire \u0/u1/_0502_ ;
wire \u0/u1/_0503_ ;
wire \u0/u1/_0504_ ;
wire \u0/u1/_0505_ ;
wire \u0/u1/_0506_ ;
wire \u0/u1/_0507_ ;
wire \u0/u1/_0508_ ;
wire \u0/u1/_0509_ ;
wire \u0/u1/_0510_ ;
wire \u0/u1/_0511_ ;
wire \u0/u1/_0512_ ;
wire \u0/u1/_0513_ ;
wire \u0/u1/_0514_ ;
wire \u0/u1/_0515_ ;
wire \u0/u1/_0516_ ;
wire \u0/u1/_0517_ ;
wire \u0/u1/_0518_ ;
wire \u0/u1/_0519_ ;
wire \u0/u1/_0520_ ;
wire \u0/u1/_0521_ ;
wire \u0/u1/_0522_ ;
wire \u0/u1/_0523_ ;
wire \u0/u1/_0524_ ;
wire \u0/u1/_0525_ ;
wire \u0/u1/_0526_ ;
wire \u0/u1/_0527_ ;
wire \u0/u1/_0528_ ;
wire \u0/u1/_0529_ ;
wire \u0/u1/_0530_ ;
wire \u0/u1/_0531_ ;
wire \u0/u1/_0532_ ;
wire \u0/u1/_0533_ ;
wire \u0/u1/_0534_ ;
wire \u0/u1/_0535_ ;
wire \u0/u1/_0536_ ;
wire \u0/u1/_0537_ ;
wire \u0/u1/_0538_ ;
wire \u0/u1/_0539_ ;
wire \u0/u1/_0540_ ;
wire \u0/u1/_0541_ ;
wire \u0/u1/_0542_ ;
wire \u0/u1/_0543_ ;
wire \u0/u1/_0544_ ;
wire \u0/u1/_0545_ ;
wire \u0/u1/_0546_ ;
wire \u0/u1/_0547_ ;
wire \u0/u1/_0548_ ;
wire \u0/u1/_0549_ ;
wire \u0/u1/_0550_ ;
wire \u0/u1/_0551_ ;
wire \u0/u1/_0552_ ;
wire \u0/u1/_0553_ ;
wire \u0/u1/_0554_ ;
wire \u0/u1/_0555_ ;
wire \u0/u1/_0556_ ;
wire \u0/u1/_0557_ ;
wire \u0/u1/_0558_ ;
wire \u0/u1/_0559_ ;
wire \u0/u1/_0560_ ;
wire \u0/u1/_0561_ ;
wire \u0/u1/_0562_ ;
wire \u0/u1/_0563_ ;
wire \u0/u1/_0565_ ;
wire \u0/u1/_0566_ ;
wire \u0/u1/_0567_ ;
wire \u0/u1/_0568_ ;
wire \u0/u1/_0569_ ;
wire \u0/u1/_0570_ ;
wire \u0/u1/_0571_ ;
wire \u0/u1/_0572_ ;
wire \u0/u1/_0573_ ;
wire \u0/u1/_0574_ ;
wire \u0/u1/_0575_ ;
wire \u0/u1/_0576_ ;
wire \u0/u1/_0577_ ;
wire \u0/u1/_0578_ ;
wire \u0/u1/_0579_ ;
wire \u0/u1/_0580_ ;
wire \u0/u1/_0581_ ;
wire \u0/u1/_0582_ ;
wire \u0/u1/_0583_ ;
wire \u0/u1/_0584_ ;
wire \u0/u1/_0585_ ;
wire \u0/u1/_0586_ ;
wire \u0/u1/_0587_ ;
wire \u0/u1/_0588_ ;
wire \u0/u1/_0589_ ;
wire \u0/u1/_0590_ ;
wire \u0/u1/_0591_ ;
wire \u0/u1/_0592_ ;
wire \u0/u1/_0593_ ;
wire \u0/u1/_0594_ ;
wire \u0/u1/_0595_ ;
wire \u0/u1/_0596_ ;
wire \u0/u1/_0598_ ;
wire \u0/u1/_0599_ ;
wire \u0/u1/_0600_ ;
wire \u0/u1/_0601_ ;
wire \u0/u1/_0602_ ;
wire \u0/u1/_0603_ ;
wire \u0/u1/_0604_ ;
wire \u0/u1/_0605_ ;
wire \u0/u1/_0606_ ;
wire \u0/u1/_0607_ ;
wire \u0/u1/_0608_ ;
wire \u0/u1/_0609_ ;
wire \u0/u1/_0610_ ;
wire \u0/u1/_0611_ ;
wire \u0/u1/_0612_ ;
wire \u0/u1/_0613_ ;
wire \u0/u1/_0614_ ;
wire \u0/u1/_0615_ ;
wire \u0/u1/_0616_ ;
wire \u0/u1/_0617_ ;
wire \u0/u1/_0618_ ;
wire \u0/u1/_0619_ ;
wire \u0/u1/_0620_ ;
wire \u0/u1/_0621_ ;
wire \u0/u1/_0622_ ;
wire \u0/u1/_0623_ ;
wire \u0/u1/_0624_ ;
wire \u0/u1/_0625_ ;
wire \u0/u1/_0626_ ;
wire \u0/u1/_0627_ ;
wire \u0/u1/_0628_ ;
wire \u0/u1/_0629_ ;
wire \u0/u1/_0630_ ;
wire \u0/u1/_0631_ ;
wire \u0/u1/_0632_ ;
wire \u0/u1/_0633_ ;
wire \u0/u1/_0634_ ;
wire \u0/u1/_0635_ ;
wire \u0/u1/_0636_ ;
wire \u0/u1/_0637_ ;
wire \u0/u1/_0638_ ;
wire \u0/u1/_0639_ ;
wire \u0/u1/_0640_ ;
wire \u0/u1/_0641_ ;
wire \u0/u1/_0642_ ;
wire \u0/u1/_0643_ ;
wire \u0/u1/_0644_ ;
wire \u0/u1/_0645_ ;
wire \u0/u1/_0646_ ;
wire \u0/u1/_0647_ ;
wire \u0/u1/_0648_ ;
wire \u0/u1/_0649_ ;
wire \u0/u1/_0650_ ;
wire \u0/u1/_0652_ ;
wire \u0/u1/_0653_ ;
wire \u0/u1/_0654_ ;
wire \u0/u1/_0655_ ;
wire \u0/u1/_0656_ ;
wire \u0/u1/_0657_ ;
wire \u0/u1/_0658_ ;
wire \u0/u1/_0659_ ;
wire \u0/u1/_0660_ ;
wire \u0/u1/_0661_ ;
wire \u0/u1/_0662_ ;
wire \u0/u1/_0663_ ;
wire \u0/u1/_0664_ ;
wire \u0/u1/_0665_ ;
wire \u0/u1/_0666_ ;
wire \u0/u1/_0667_ ;
wire \u0/u1/_0668_ ;
wire \u0/u1/_0669_ ;
wire \u0/u1/_0670_ ;
wire \u0/u1/_0671_ ;
wire \u0/u1/_0673_ ;
wire \u0/u1/_0674_ ;
wire \u0/u1/_0675_ ;
wire \u0/u1/_0676_ ;
wire \u0/u1/_0677_ ;
wire \u0/u1/_0678_ ;
wire \u0/u1/_0679_ ;
wire \u0/u1/_0680_ ;
wire \u0/u1/_0681_ ;
wire \u0/u1/_0682_ ;
wire \u0/u1/_0683_ ;
wire \u0/u1/_0684_ ;
wire \u0/u1/_0685_ ;
wire \u0/u1/_0686_ ;
wire \u0/u1/_0687_ ;
wire \u0/u1/_0688_ ;
wire \u0/u1/_0689_ ;
wire \u0/u1/_0690_ ;
wire \u0/u1/_0691_ ;
wire \u0/u1/_0692_ ;
wire \u0/u1/_0693_ ;
wire \u0/u1/_0694_ ;
wire \u0/u1/_0695_ ;
wire \u0/u1/_0696_ ;
wire \u0/u1/_0697_ ;
wire \u0/u1/_0698_ ;
wire \u0/u1/_0699_ ;
wire \u0/u1/_0700_ ;
wire \u0/u1/_0701_ ;
wire \u0/u1/_0702_ ;
wire \u0/u1/_0703_ ;
wire \u0/u1/_0704_ ;
wire \u0/u1/_0705_ ;
wire \u0/u1/_0706_ ;
wire \u0/u1/_0707_ ;
wire \u0/u1/_0708_ ;
wire \u0/u1/_0709_ ;
wire \u0/u1/_0710_ ;
wire \u0/u1/_0711_ ;
wire \u0/u1/_0712_ ;
wire \u0/u1/_0713_ ;
wire \u0/u1/_0714_ ;
wire \u0/u1/_0715_ ;
wire \u0/u1/_0717_ ;
wire \u0/u1/_0718_ ;
wire \u0/u1/_0719_ ;
wire \u0/u1/_0720_ ;
wire \u0/u1/_0721_ ;
wire \u0/u1/_0722_ ;
wire \u0/u1/_0723_ ;
wire \u0/u1/_0724_ ;
wire \u0/u1/_0725_ ;
wire \u0/u1/_0726_ ;
wire \u0/u1/_0727_ ;
wire \u0/u1/_0728_ ;
wire \u0/u1/_0729_ ;
wire \u0/u1/_0730_ ;
wire \u0/u1/_0731_ ;
wire \u0/u1/_0733_ ;
wire \u0/u1/_0734_ ;
wire \u0/u1/_0735_ ;
wire \u0/u1/_0736_ ;
wire \u0/u1/_0738_ ;
wire \u0/u1/_0739_ ;
wire \u0/u1/_0740_ ;
wire \u0/u1/_0741_ ;
wire \u0/u1/_0742_ ;
wire \u0/u1/_0744_ ;
wire \u0/u1/_0745_ ;
wire \u0/u1/_0746_ ;
wire \u0/u1/_0748_ ;
wire \u0/u1/_0749_ ;
wire \u0/u1/_0750_ ;
wire \u0/u1/_0752_ ;
wire \u0/u2/_0008_ ;
wire \u0/u2/_0009_ ;
wire \u0/u2/_0010_ ;
wire \u0/u2/_0011_ ;
wire \u0/u2/_0012_ ;
wire \u0/u2/_0013_ ;
wire \u0/u2/_0014_ ;
wire \u0/u2/_0015_ ;
wire \u0/u2/_0016_ ;
wire \u0/u2/_0017_ ;
wire \u0/u2/_0019_ ;
wire \u0/u2/_0020_ ;
wire \u0/u2/_0022_ ;
wire \u0/u2/_0024_ ;
wire \u0/u2/_0025_ ;
wire \u0/u2/_0026_ ;
wire \u0/u2/_0027_ ;
wire \u0/u2/_0030_ ;
wire \u0/u2/_0032_ ;
wire \u0/u2/_0033_ ;
wire \u0/u2/_0034_ ;
wire \u0/u2/_0035_ ;
wire \u0/u2/_0037_ ;
wire \u0/u2/_0038_ ;
wire \u0/u2/_0039_ ;
wire \u0/u2/_0040_ ;
wire \u0/u2/_0041_ ;
wire \u0/u2/_0042_ ;
wire \u0/u2/_0043_ ;
wire \u0/u2/_0045_ ;
wire \u0/u2/_0046_ ;
wire \u0/u2/_0047_ ;
wire \u0/u2/_0049_ ;
wire \u0/u2/_0050_ ;
wire \u0/u2/_0051_ ;
wire \u0/u2/_0052_ ;
wire \u0/u2/_0053_ ;
wire \u0/u2/_0054_ ;
wire \u0/u2/_0056_ ;
wire \u0/u2/_0057_ ;
wire \u0/u2/_0058_ ;
wire \u0/u2/_0060_ ;
wire \u0/u2/_0061_ ;
wire \u0/u2/_0062_ ;
wire \u0/u2/_0064_ ;
wire \u0/u2/_0065_ ;
wire \u0/u2/_0066_ ;
wire \u0/u2/_0067_ ;
wire \u0/u2/_0069_ ;
wire \u0/u2/_0070_ ;
wire \u0/u2/_0072_ ;
wire \u0/u2/_0073_ ;
wire \u0/u2/_0074_ ;
wire \u0/u2/_0075_ ;
wire \u0/u2/_0076_ ;
wire \u0/u2/_0077_ ;
wire \u0/u2/_0078_ ;
wire \u0/u2/_0079_ ;
wire \u0/u2/_0081_ ;
wire \u0/u2/_0082_ ;
wire \u0/u2/_0085_ ;
wire \u0/u2/_0086_ ;
wire \u0/u2/_0087_ ;
wire \u0/u2/_0088_ ;
wire \u0/u2/_0089_ ;
wire \u0/u2/_0090_ ;
wire \u0/u2/_0091_ ;
wire \u0/u2/_0092_ ;
wire \u0/u2/_0093_ ;
wire \u0/u2/_0094_ ;
wire \u0/u2/_0095_ ;
wire \u0/u2/_0096_ ;
wire \u0/u2/_0097_ ;
wire \u0/u2/_0098_ ;
wire \u0/u2/_0099_ ;
wire \u0/u2/_0100_ ;
wire \u0/u2/_0101_ ;
wire \u0/u2/_0102_ ;
wire \u0/u2/_0103_ ;
wire \u0/u2/_0104_ ;
wire \u0/u2/_0105_ ;
wire \u0/u2/_0106_ ;
wire \u0/u2/_0108_ ;
wire \u0/u2/_0109_ ;
wire \u0/u2/_0110_ ;
wire \u0/u2/_0111_ ;
wire \u0/u2/_0113_ ;
wire \u0/u2/_0114_ ;
wire \u0/u2/_0115_ ;
wire \u0/u2/_0116_ ;
wire \u0/u2/_0117_ ;
wire \u0/u2/_0118_ ;
wire \u0/u2/_0119_ ;
wire \u0/u2/_0120_ ;
wire \u0/u2/_0121_ ;
wire \u0/u2/_0122_ ;
wire \u0/u2/_0123_ ;
wire \u0/u2/_0124_ ;
wire \u0/u2/_0126_ ;
wire \u0/u2/_0127_ ;
wire \u0/u2/_0128_ ;
wire \u0/u2/_0129_ ;
wire \u0/u2/_0130_ ;
wire \u0/u2/_0132_ ;
wire \u0/u2/_0133_ ;
wire \u0/u2/_0135_ ;
wire \u0/u2/_0136_ ;
wire \u0/u2/_0137_ ;
wire \u0/u2/_0139_ ;
wire \u0/u2/_0140_ ;
wire \u0/u2/_0141_ ;
wire \u0/u2/_0142_ ;
wire \u0/u2/_0144_ ;
wire \u0/u2/_0145_ ;
wire \u0/u2/_0146_ ;
wire \u0/u2/_0147_ ;
wire \u0/u2/_0148_ ;
wire \u0/u2/_0149_ ;
wire \u0/u2/_0150_ ;
wire \u0/u2/_0151_ ;
wire \u0/u2/_0153_ ;
wire \u0/u2/_0154_ ;
wire \u0/u2/_0155_ ;
wire \u0/u2/_0156_ ;
wire \u0/u2/_0157_ ;
wire \u0/u2/_0158_ ;
wire \u0/u2/_0159_ ;
wire \u0/u2/_0161_ ;
wire \u0/u2/_0162_ ;
wire \u0/u2/_0163_ ;
wire \u0/u2/_0164_ ;
wire \u0/u2/_0165_ ;
wire \u0/u2/_0166_ ;
wire \u0/u2/_0167_ ;
wire \u0/u2/_0168_ ;
wire \u0/u2/_0169_ ;
wire \u0/u2/_0170_ ;
wire \u0/u2/_0171_ ;
wire \u0/u2/_0172_ ;
wire \u0/u2/_0174_ ;
wire \u0/u2/_0175_ ;
wire \u0/u2/_0176_ ;
wire \u0/u2/_0177_ ;
wire \u0/u2/_0178_ ;
wire \u0/u2/_0179_ ;
wire \u0/u2/_0180_ ;
wire \u0/u2/_0181_ ;
wire \u0/u2/_0182_ ;
wire \u0/u2/_0183_ ;
wire \u0/u2/_0184_ ;
wire \u0/u2/_0185_ ;
wire \u0/u2/_0186_ ;
wire \u0/u2/_0187_ ;
wire \u0/u2/_0188_ ;
wire \u0/u2/_0189_ ;
wire \u0/u2/_0190_ ;
wire \u0/u2/_0191_ ;
wire \u0/u2/_0192_ ;
wire \u0/u2/_0193_ ;
wire \u0/u2/_0194_ ;
wire \u0/u2/_0195_ ;
wire \u0/u2/_0196_ ;
wire \u0/u2/_0197_ ;
wire \u0/u2/_0198_ ;
wire \u0/u2/_0199_ ;
wire \u0/u2/_0200_ ;
wire \u0/u2/_0201_ ;
wire \u0/u2/_0202_ ;
wire \u0/u2/_0203_ ;
wire \u0/u2/_0204_ ;
wire \u0/u2/_0205_ ;
wire \u0/u2/_0206_ ;
wire \u0/u2/_0207_ ;
wire \u0/u2/_0208_ ;
wire \u0/u2/_0209_ ;
wire \u0/u2/_0210_ ;
wire \u0/u2/_0211_ ;
wire \u0/u2/_0212_ ;
wire \u0/u2/_0213_ ;
wire \u0/u2/_0214_ ;
wire \u0/u2/_0215_ ;
wire \u0/u2/_0216_ ;
wire \u0/u2/_0217_ ;
wire \u0/u2/_0219_ ;
wire \u0/u2/_0220_ ;
wire \u0/u2/_0221_ ;
wire \u0/u2/_0222_ ;
wire \u0/u2/_0223_ ;
wire \u0/u2/_0224_ ;
wire \u0/u2/_0225_ ;
wire \u0/u2/_0226_ ;
wire \u0/u2/_0227_ ;
wire \u0/u2/_0228_ ;
wire \u0/u2/_0229_ ;
wire \u0/u2/_0230_ ;
wire \u0/u2/_0231_ ;
wire \u0/u2/_0232_ ;
wire \u0/u2/_0233_ ;
wire \u0/u2/_0234_ ;
wire \u0/u2/_0235_ ;
wire \u0/u2/_0236_ ;
wire \u0/u2/_0237_ ;
wire \u0/u2/_0238_ ;
wire \u0/u2/_0239_ ;
wire \u0/u2/_0240_ ;
wire \u0/u2/_0241_ ;
wire \u0/u2/_0242_ ;
wire \u0/u2/_0243_ ;
wire \u0/u2/_0244_ ;
wire \u0/u2/_0245_ ;
wire \u0/u2/_0246_ ;
wire \u0/u2/_0247_ ;
wire \u0/u2/_0248_ ;
wire \u0/u2/_0249_ ;
wire \u0/u2/_0250_ ;
wire \u0/u2/_0251_ ;
wire \u0/u2/_0252_ ;
wire \u0/u2/_0253_ ;
wire \u0/u2/_0254_ ;
wire \u0/u2/_0255_ ;
wire \u0/u2/_0256_ ;
wire \u0/u2/_0257_ ;
wire \u0/u2/_0258_ ;
wire \u0/u2/_0259_ ;
wire \u0/u2/_0260_ ;
wire \u0/u2/_0261_ ;
wire \u0/u2/_0263_ ;
wire \u0/u2/_0264_ ;
wire \u0/u2/_0265_ ;
wire \u0/u2/_0266_ ;
wire \u0/u2/_0267_ ;
wire \u0/u2/_0268_ ;
wire \u0/u2/_0269_ ;
wire \u0/u2/_0270_ ;
wire \u0/u2/_0271_ ;
wire \u0/u2/_0272_ ;
wire \u0/u2/_0273_ ;
wire \u0/u2/_0274_ ;
wire \u0/u2/_0275_ ;
wire \u0/u2/_0276_ ;
wire \u0/u2/_0277_ ;
wire \u0/u2/_0278_ ;
wire \u0/u2/_0279_ ;
wire \u0/u2/_0280_ ;
wire \u0/u2/_0281_ ;
wire \u0/u2/_0283_ ;
wire \u0/u2/_0284_ ;
wire \u0/u2/_0285_ ;
wire \u0/u2/_0286_ ;
wire \u0/u2/_0287_ ;
wire \u0/u2/_0288_ ;
wire \u0/u2/_0289_ ;
wire \u0/u2/_0290_ ;
wire \u0/u2/_0291_ ;
wire \u0/u2/_0293_ ;
wire \u0/u2/_0294_ ;
wire \u0/u2/_0295_ ;
wire \u0/u2/_0296_ ;
wire \u0/u2/_0297_ ;
wire \u0/u2/_0298_ ;
wire \u0/u2/_0299_ ;
wire \u0/u2/_0300_ ;
wire \u0/u2/_0301_ ;
wire \u0/u2/_0302_ ;
wire \u0/u2/_0303_ ;
wire \u0/u2/_0304_ ;
wire \u0/u2/_0305_ ;
wire \u0/u2/_0306_ ;
wire \u0/u2/_0307_ ;
wire \u0/u2/_0308_ ;
wire \u0/u2/_0309_ ;
wire \u0/u2/_0310_ ;
wire \u0/u2/_0311_ ;
wire \u0/u2/_0312_ ;
wire \u0/u2/_0313_ ;
wire \u0/u2/_0314_ ;
wire \u0/u2/_0315_ ;
wire \u0/u2/_0316_ ;
wire \u0/u2/_0317_ ;
wire \u0/u2/_0318_ ;
wire \u0/u2/_0319_ ;
wire \u0/u2/_0320_ ;
wire \u0/u2/_0321_ ;
wire \u0/u2/_0322_ ;
wire \u0/u2/_0323_ ;
wire \u0/u2/_0324_ ;
wire \u0/u2/_0325_ ;
wire \u0/u2/_0326_ ;
wire \u0/u2/_0327_ ;
wire \u0/u2/_0328_ ;
wire \u0/u2/_0329_ ;
wire \u0/u2/_0330_ ;
wire \u0/u2/_0331_ ;
wire \u0/u2/_0332_ ;
wire \u0/u2/_0333_ ;
wire \u0/u2/_0334_ ;
wire \u0/u2/_0335_ ;
wire \u0/u2/_0337_ ;
wire \u0/u2/_0338_ ;
wire \u0/u2/_0339_ ;
wire \u0/u2/_0340_ ;
wire \u0/u2/_0341_ ;
wire \u0/u2/_0342_ ;
wire \u0/u2/_0343_ ;
wire \u0/u2/_0344_ ;
wire \u0/u2/_0345_ ;
wire \u0/u2/_0347_ ;
wire \u0/u2/_0348_ ;
wire \u0/u2/_0349_ ;
wire \u0/u2/_0350_ ;
wire \u0/u2/_0351_ ;
wire \u0/u2/_0352_ ;
wire \u0/u2/_0353_ ;
wire \u0/u2/_0354_ ;
wire \u0/u2/_0355_ ;
wire \u0/u2/_0356_ ;
wire \u0/u2/_0357_ ;
wire \u0/u2/_0358_ ;
wire \u0/u2/_0359_ ;
wire \u0/u2/_0360_ ;
wire \u0/u2/_0361_ ;
wire \u0/u2/_0362_ ;
wire \u0/u2/_0363_ ;
wire \u0/u2/_0365_ ;
wire \u0/u2/_0366_ ;
wire \u0/u2/_0367_ ;
wire \u0/u2/_0368_ ;
wire \u0/u2/_0370_ ;
wire \u0/u2/_0371_ ;
wire \u0/u2/_0372_ ;
wire \u0/u2/_0373_ ;
wire \u0/u2/_0374_ ;
wire \u0/u2/_0375_ ;
wire \u0/u2/_0376_ ;
wire \u0/u2/_0377_ ;
wire \u0/u2/_0378_ ;
wire \u0/u2/_0379_ ;
wire \u0/u2/_0380_ ;
wire \u0/u2/_0381_ ;
wire \u0/u2/_0382_ ;
wire \u0/u2/_0383_ ;
wire \u0/u2/_0384_ ;
wire \u0/u2/_0385_ ;
wire \u0/u2/_0386_ ;
wire \u0/u2/_0387_ ;
wire \u0/u2/_0388_ ;
wire \u0/u2/_0389_ ;
wire \u0/u2/_0390_ ;
wire \u0/u2/_0391_ ;
wire \u0/u2/_0392_ ;
wire \u0/u2/_0393_ ;
wire \u0/u2/_0394_ ;
wire \u0/u2/_0395_ ;
wire \u0/u2/_0396_ ;
wire \u0/u2/_0397_ ;
wire \u0/u2/_0398_ ;
wire \u0/u2/_0399_ ;
wire \u0/u2/_0400_ ;
wire \u0/u2/_0401_ ;
wire \u0/u2/_0402_ ;
wire \u0/u2/_0403_ ;
wire \u0/u2/_0404_ ;
wire \u0/u2/_0405_ ;
wire \u0/u2/_0406_ ;
wire \u0/u2/_0407_ ;
wire \u0/u2/_0408_ ;
wire \u0/u2/_0409_ ;
wire \u0/u2/_0410_ ;
wire \u0/u2/_0411_ ;
wire \u0/u2/_0412_ ;
wire \u0/u2/_0413_ ;
wire \u0/u2/_0414_ ;
wire \u0/u2/_0415_ ;
wire \u0/u2/_0416_ ;
wire \u0/u2/_0417_ ;
wire \u0/u2/_0418_ ;
wire \u0/u2/_0419_ ;
wire \u0/u2/_0420_ ;
wire \u0/u2/_0421_ ;
wire \u0/u2/_0422_ ;
wire \u0/u2/_0423_ ;
wire \u0/u2/_0424_ ;
wire \u0/u2/_0425_ ;
wire \u0/u2/_0426_ ;
wire \u0/u2/_0427_ ;
wire \u0/u2/_0428_ ;
wire \u0/u2/_0429_ ;
wire \u0/u2/_0430_ ;
wire \u0/u2/_0431_ ;
wire \u0/u2/_0432_ ;
wire \u0/u2/_0433_ ;
wire \u0/u2/_0434_ ;
wire \u0/u2/_0435_ ;
wire \u0/u2/_0436_ ;
wire \u0/u2/_0437_ ;
wire \u0/u2/_0438_ ;
wire \u0/u2/_0439_ ;
wire \u0/u2/_0440_ ;
wire \u0/u2/_0441_ ;
wire \u0/u2/_0442_ ;
wire \u0/u2/_0443_ ;
wire \u0/u2/_0444_ ;
wire \u0/u2/_0446_ ;
wire \u0/u2/_0447_ ;
wire \u0/u2/_0448_ ;
wire \u0/u2/_0449_ ;
wire \u0/u2/_0450_ ;
wire \u0/u2/_0451_ ;
wire \u0/u2/_0452_ ;
wire \u0/u2/_0453_ ;
wire \u0/u2/_0454_ ;
wire \u0/u2/_0455_ ;
wire \u0/u2/_0456_ ;
wire \u0/u2/_0457_ ;
wire \u0/u2/_0458_ ;
wire \u0/u2/_0459_ ;
wire \u0/u2/_0460_ ;
wire \u0/u2/_0461_ ;
wire \u0/u2/_0462_ ;
wire \u0/u2/_0463_ ;
wire \u0/u2/_0464_ ;
wire \u0/u2/_0465_ ;
wire \u0/u2/_0466_ ;
wire \u0/u2/_0467_ ;
wire \u0/u2/_0468_ ;
wire \u0/u2/_0469_ ;
wire \u0/u2/_0470_ ;
wire \u0/u2/_0471_ ;
wire \u0/u2/_0472_ ;
wire \u0/u2/_0473_ ;
wire \u0/u2/_0474_ ;
wire \u0/u2/_0475_ ;
wire \u0/u2/_0476_ ;
wire \u0/u2/_0477_ ;
wire \u0/u2/_0478_ ;
wire \u0/u2/_0479_ ;
wire \u0/u2/_0480_ ;
wire \u0/u2/_0481_ ;
wire \u0/u2/_0482_ ;
wire \u0/u2/_0483_ ;
wire \u0/u2/_0484_ ;
wire \u0/u2/_0485_ ;
wire \u0/u2/_0486_ ;
wire \u0/u2/_0487_ ;
wire \u0/u2/_0488_ ;
wire \u0/u2/_0490_ ;
wire \u0/u2/_0491_ ;
wire \u0/u2/_0492_ ;
wire \u0/u2/_0493_ ;
wire \u0/u2/_0494_ ;
wire \u0/u2/_0495_ ;
wire \u0/u2/_0496_ ;
wire \u0/u2/_0497_ ;
wire \u0/u2/_0498_ ;
wire \u0/u2/_0499_ ;
wire \u0/u2/_0500_ ;
wire \u0/u2/_0501_ ;
wire \u0/u2/_0502_ ;
wire \u0/u2/_0503_ ;
wire \u0/u2/_0504_ ;
wire \u0/u2/_0505_ ;
wire \u0/u2/_0506_ ;
wire \u0/u2/_0507_ ;
wire \u0/u2/_0508_ ;
wire \u0/u2/_0509_ ;
wire \u0/u2/_0510_ ;
wire \u0/u2/_0511_ ;
wire \u0/u2/_0512_ ;
wire \u0/u2/_0513_ ;
wire \u0/u2/_0514_ ;
wire \u0/u2/_0515_ ;
wire \u0/u2/_0516_ ;
wire \u0/u2/_0517_ ;
wire \u0/u2/_0518_ ;
wire \u0/u2/_0519_ ;
wire \u0/u2/_0520_ ;
wire \u0/u2/_0521_ ;
wire \u0/u2/_0522_ ;
wire \u0/u2/_0523_ ;
wire \u0/u2/_0524_ ;
wire \u0/u2/_0525_ ;
wire \u0/u2/_0526_ ;
wire \u0/u2/_0527_ ;
wire \u0/u2/_0528_ ;
wire \u0/u2/_0529_ ;
wire \u0/u2/_0530_ ;
wire \u0/u2/_0531_ ;
wire \u0/u2/_0532_ ;
wire \u0/u2/_0533_ ;
wire \u0/u2/_0534_ ;
wire \u0/u2/_0535_ ;
wire \u0/u2/_0536_ ;
wire \u0/u2/_0537_ ;
wire \u0/u2/_0538_ ;
wire \u0/u2/_0539_ ;
wire \u0/u2/_0540_ ;
wire \u0/u2/_0541_ ;
wire \u0/u2/_0542_ ;
wire \u0/u2/_0543_ ;
wire \u0/u2/_0544_ ;
wire \u0/u2/_0545_ ;
wire \u0/u2/_0546_ ;
wire \u0/u2/_0547_ ;
wire \u0/u2/_0548_ ;
wire \u0/u2/_0549_ ;
wire \u0/u2/_0550_ ;
wire \u0/u2/_0551_ ;
wire \u0/u2/_0552_ ;
wire \u0/u2/_0553_ ;
wire \u0/u2/_0554_ ;
wire \u0/u2/_0555_ ;
wire \u0/u2/_0556_ ;
wire \u0/u2/_0557_ ;
wire \u0/u2/_0558_ ;
wire \u0/u2/_0559_ ;
wire \u0/u2/_0560_ ;
wire \u0/u2/_0561_ ;
wire \u0/u2/_0562_ ;
wire \u0/u2/_0563_ ;
wire \u0/u2/_0565_ ;
wire \u0/u2/_0566_ ;
wire \u0/u2/_0567_ ;
wire \u0/u2/_0568_ ;
wire \u0/u2/_0569_ ;
wire \u0/u2/_0570_ ;
wire \u0/u2/_0571_ ;
wire \u0/u2/_0572_ ;
wire \u0/u2/_0573_ ;
wire \u0/u2/_0574_ ;
wire \u0/u2/_0575_ ;
wire \u0/u2/_0576_ ;
wire \u0/u2/_0577_ ;
wire \u0/u2/_0578_ ;
wire \u0/u2/_0579_ ;
wire \u0/u2/_0580_ ;
wire \u0/u2/_0581_ ;
wire \u0/u2/_0582_ ;
wire \u0/u2/_0583_ ;
wire \u0/u2/_0584_ ;
wire \u0/u2/_0585_ ;
wire \u0/u2/_0586_ ;
wire \u0/u2/_0587_ ;
wire \u0/u2/_0588_ ;
wire \u0/u2/_0589_ ;
wire \u0/u2/_0590_ ;
wire \u0/u2/_0591_ ;
wire \u0/u2/_0592_ ;
wire \u0/u2/_0593_ ;
wire \u0/u2/_0594_ ;
wire \u0/u2/_0595_ ;
wire \u0/u2/_0596_ ;
wire \u0/u2/_0598_ ;
wire \u0/u2/_0599_ ;
wire \u0/u2/_0600_ ;
wire \u0/u2/_0601_ ;
wire \u0/u2/_0602_ ;
wire \u0/u2/_0603_ ;
wire \u0/u2/_0604_ ;
wire \u0/u2/_0605_ ;
wire \u0/u2/_0606_ ;
wire \u0/u2/_0607_ ;
wire \u0/u2/_0608_ ;
wire \u0/u2/_0609_ ;
wire \u0/u2/_0610_ ;
wire \u0/u2/_0611_ ;
wire \u0/u2/_0612_ ;
wire \u0/u2/_0613_ ;
wire \u0/u2/_0614_ ;
wire \u0/u2/_0615_ ;
wire \u0/u2/_0616_ ;
wire \u0/u2/_0617_ ;
wire \u0/u2/_0618_ ;
wire \u0/u2/_0619_ ;
wire \u0/u2/_0620_ ;
wire \u0/u2/_0621_ ;
wire \u0/u2/_0622_ ;
wire \u0/u2/_0623_ ;
wire \u0/u2/_0624_ ;
wire \u0/u2/_0625_ ;
wire \u0/u2/_0626_ ;
wire \u0/u2/_0627_ ;
wire \u0/u2/_0628_ ;
wire \u0/u2/_0629_ ;
wire \u0/u2/_0630_ ;
wire \u0/u2/_0631_ ;
wire \u0/u2/_0632_ ;
wire \u0/u2/_0633_ ;
wire \u0/u2/_0634_ ;
wire \u0/u2/_0635_ ;
wire \u0/u2/_0636_ ;
wire \u0/u2/_0637_ ;
wire \u0/u2/_0638_ ;
wire \u0/u2/_0639_ ;
wire \u0/u2/_0640_ ;
wire \u0/u2/_0641_ ;
wire \u0/u2/_0642_ ;
wire \u0/u2/_0643_ ;
wire \u0/u2/_0644_ ;
wire \u0/u2/_0645_ ;
wire \u0/u2/_0646_ ;
wire \u0/u2/_0647_ ;
wire \u0/u2/_0648_ ;
wire \u0/u2/_0649_ ;
wire \u0/u2/_0650_ ;
wire \u0/u2/_0652_ ;
wire \u0/u2/_0653_ ;
wire \u0/u2/_0654_ ;
wire \u0/u2/_0655_ ;
wire \u0/u2/_0656_ ;
wire \u0/u2/_0657_ ;
wire \u0/u2/_0658_ ;
wire \u0/u2/_0659_ ;
wire \u0/u2/_0660_ ;
wire \u0/u2/_0661_ ;
wire \u0/u2/_0662_ ;
wire \u0/u2/_0663_ ;
wire \u0/u2/_0664_ ;
wire \u0/u2/_0665_ ;
wire \u0/u2/_0666_ ;
wire \u0/u2/_0667_ ;
wire \u0/u2/_0668_ ;
wire \u0/u2/_0669_ ;
wire \u0/u2/_0670_ ;
wire \u0/u2/_0671_ ;
wire \u0/u2/_0673_ ;
wire \u0/u2/_0674_ ;
wire \u0/u2/_0675_ ;
wire \u0/u2/_0676_ ;
wire \u0/u2/_0677_ ;
wire \u0/u2/_0678_ ;
wire \u0/u2/_0679_ ;
wire \u0/u2/_0680_ ;
wire \u0/u2/_0681_ ;
wire \u0/u2/_0682_ ;
wire \u0/u2/_0683_ ;
wire \u0/u2/_0684_ ;
wire \u0/u2/_0685_ ;
wire \u0/u2/_0686_ ;
wire \u0/u2/_0687_ ;
wire \u0/u2/_0688_ ;
wire \u0/u2/_0689_ ;
wire \u0/u2/_0690_ ;
wire \u0/u2/_0691_ ;
wire \u0/u2/_0692_ ;
wire \u0/u2/_0693_ ;
wire \u0/u2/_0694_ ;
wire \u0/u2/_0695_ ;
wire \u0/u2/_0696_ ;
wire \u0/u2/_0697_ ;
wire \u0/u2/_0698_ ;
wire \u0/u2/_0699_ ;
wire \u0/u2/_0700_ ;
wire \u0/u2/_0701_ ;
wire \u0/u2/_0702_ ;
wire \u0/u2/_0703_ ;
wire \u0/u2/_0704_ ;
wire \u0/u2/_0705_ ;
wire \u0/u2/_0706_ ;
wire \u0/u2/_0707_ ;
wire \u0/u2/_0708_ ;
wire \u0/u2/_0709_ ;
wire \u0/u2/_0710_ ;
wire \u0/u2/_0711_ ;
wire \u0/u2/_0712_ ;
wire \u0/u2/_0713_ ;
wire \u0/u2/_0714_ ;
wire \u0/u2/_0715_ ;
wire \u0/u2/_0717_ ;
wire \u0/u2/_0718_ ;
wire \u0/u2/_0719_ ;
wire \u0/u2/_0720_ ;
wire \u0/u2/_0721_ ;
wire \u0/u2/_0722_ ;
wire \u0/u2/_0723_ ;
wire \u0/u2/_0724_ ;
wire \u0/u2/_0725_ ;
wire \u0/u2/_0726_ ;
wire \u0/u2/_0727_ ;
wire \u0/u2/_0728_ ;
wire \u0/u2/_0729_ ;
wire \u0/u2/_0730_ ;
wire \u0/u2/_0731_ ;
wire \u0/u2/_0733_ ;
wire \u0/u2/_0734_ ;
wire \u0/u2/_0735_ ;
wire \u0/u2/_0736_ ;
wire \u0/u2/_0738_ ;
wire \u0/u2/_0739_ ;
wire \u0/u2/_0740_ ;
wire \u0/u2/_0741_ ;
wire \u0/u2/_0742_ ;
wire \u0/u2/_0744_ ;
wire \u0/u2/_0745_ ;
wire \u0/u2/_0746_ ;
wire \u0/u2/_0748_ ;
wire \u0/u2/_0749_ ;
wire \u0/u2/_0750_ ;
wire \u0/u2/_0752_ ;
wire \u0/u3/_0007_ ;
wire \u0/u3/_0008_ ;
wire \u0/u3/_0009_ ;
wire \u0/u3/_0010_ ;
wire \u0/u3/_0011_ ;
wire \u0/u3/_0012_ ;
wire \u0/u3/_0013_ ;
wire \u0/u3/_0014_ ;
wire \u0/u3/_0015_ ;
wire \u0/u3/_0016_ ;
wire \u0/u3/_0017_ ;
wire \u0/u3/_0019_ ;
wire \u0/u3/_0020_ ;
wire \u0/u3/_0022_ ;
wire \u0/u3/_0024_ ;
wire \u0/u3/_0025_ ;
wire \u0/u3/_0026_ ;
wire \u0/u3/_0027_ ;
wire \u0/u3/_0029_ ;
wire \u0/u3/_0030_ ;
wire \u0/u3/_0032_ ;
wire \u0/u3/_0033_ ;
wire \u0/u3/_0034_ ;
wire \u0/u3/_0035_ ;
wire \u0/u3/_0037_ ;
wire \u0/u3/_0038_ ;
wire \u0/u3/_0039_ ;
wire \u0/u3/_0040_ ;
wire \u0/u3/_0041_ ;
wire \u0/u3/_0042_ ;
wire \u0/u3/_0043_ ;
wire \u0/u3/_0045_ ;
wire \u0/u3/_0046_ ;
wire \u0/u3/_0047_ ;
wire \u0/u3/_0049_ ;
wire \u0/u3/_0050_ ;
wire \u0/u3/_0051_ ;
wire \u0/u3/_0052_ ;
wire \u0/u3/_0053_ ;
wire \u0/u3/_0054_ ;
wire \u0/u3/_0057_ ;
wire \u0/u3/_0058_ ;
wire \u0/u3/_0060_ ;
wire \u0/u3/_0061_ ;
wire \u0/u3/_0062_ ;
wire \u0/u3/_0064_ ;
wire \u0/u3/_0065_ ;
wire \u0/u3/_0066_ ;
wire \u0/u3/_0067_ ;
wire \u0/u3/_0069_ ;
wire \u0/u3/_0070_ ;
wire \u0/u3/_0072_ ;
wire \u0/u3/_0073_ ;
wire \u0/u3/_0074_ ;
wire \u0/u3/_0075_ ;
wire \u0/u3/_0076_ ;
wire \u0/u3/_0077_ ;
wire \u0/u3/_0078_ ;
wire \u0/u3/_0079_ ;
wire \u0/u3/_0081_ ;
wire \u0/u3/_0082_ ;
wire \u0/u3/_0084_ ;
wire \u0/u3/_0085_ ;
wire \u0/u3/_0086_ ;
wire \u0/u3/_0087_ ;
wire \u0/u3/_0088_ ;
wire \u0/u3/_0089_ ;
wire \u0/u3/_0090_ ;
wire \u0/u3/_0091_ ;
wire \u0/u3/_0092_ ;
wire \u0/u3/_0093_ ;
wire \u0/u3/_0094_ ;
wire \u0/u3/_0095_ ;
wire \u0/u3/_0096_ ;
wire \u0/u3/_0097_ ;
wire \u0/u3/_0098_ ;
wire \u0/u3/_0100_ ;
wire \u0/u3/_0101_ ;
wire \u0/u3/_0102_ ;
wire \u0/u3/_0103_ ;
wire \u0/u3/_0104_ ;
wire \u0/u3/_0105_ ;
wire \u0/u3/_0106_ ;
wire \u0/u3/_0108_ ;
wire \u0/u3/_0109_ ;
wire \u0/u3/_0110_ ;
wire \u0/u3/_0111_ ;
wire \u0/u3/_0113_ ;
wire \u0/u3/_0114_ ;
wire \u0/u3/_0115_ ;
wire \u0/u3/_0116_ ;
wire \u0/u3/_0117_ ;
wire \u0/u3/_0118_ ;
wire \u0/u3/_0119_ ;
wire \u0/u3/_0120_ ;
wire \u0/u3/_0121_ ;
wire \u0/u3/_0122_ ;
wire \u0/u3/_0123_ ;
wire \u0/u3/_0124_ ;
wire \u0/u3/_0126_ ;
wire \u0/u3/_0127_ ;
wire \u0/u3/_0128_ ;
wire \u0/u3/_0129_ ;
wire \u0/u3/_0130_ ;
wire \u0/u3/_0132_ ;
wire \u0/u3/_0133_ ;
wire \u0/u3/_0134_ ;
wire \u0/u3/_0135_ ;
wire \u0/u3/_0136_ ;
wire \u0/u3/_0137_ ;
wire \u0/u3/_0139_ ;
wire \u0/u3/_0140_ ;
wire \u0/u3/_0141_ ;
wire \u0/u3/_0142_ ;
wire \u0/u3/_0144_ ;
wire \u0/u3/_0145_ ;
wire \u0/u3/_0146_ ;
wire \u0/u3/_0147_ ;
wire \u0/u3/_0148_ ;
wire \u0/u3/_0149_ ;
wire \u0/u3/_0150_ ;
wire \u0/u3/_0151_ ;
wire \u0/u3/_0153_ ;
wire \u0/u3/_0154_ ;
wire \u0/u3/_0155_ ;
wire \u0/u3/_0156_ ;
wire \u0/u3/_0157_ ;
wire \u0/u3/_0158_ ;
wire \u0/u3/_0159_ ;
wire \u0/u3/_0161_ ;
wire \u0/u3/_0162_ ;
wire \u0/u3/_0163_ ;
wire \u0/u3/_0164_ ;
wire \u0/u3/_0165_ ;
wire \u0/u3/_0166_ ;
wire \u0/u3/_0167_ ;
wire \u0/u3/_0168_ ;
wire \u0/u3/_0169_ ;
wire \u0/u3/_0170_ ;
wire \u0/u3/_0171_ ;
wire \u0/u3/_0172_ ;
wire \u0/u3/_0174_ ;
wire \u0/u3/_0175_ ;
wire \u0/u3/_0176_ ;
wire \u0/u3/_0177_ ;
wire \u0/u3/_0178_ ;
wire \u0/u3/_0179_ ;
wire \u0/u3/_0180_ ;
wire \u0/u3/_0181_ ;
wire \u0/u3/_0182_ ;
wire \u0/u3/_0183_ ;
wire \u0/u3/_0184_ ;
wire \u0/u3/_0185_ ;
wire \u0/u3/_0186_ ;
wire \u0/u3/_0187_ ;
wire \u0/u3/_0188_ ;
wire \u0/u3/_0189_ ;
wire \u0/u3/_0190_ ;
wire \u0/u3/_0191_ ;
wire \u0/u3/_0192_ ;
wire \u0/u3/_0193_ ;
wire \u0/u3/_0194_ ;
wire \u0/u3/_0195_ ;
wire \u0/u3/_0196_ ;
wire \u0/u3/_0197_ ;
wire \u0/u3/_0198_ ;
wire \u0/u3/_0199_ ;
wire \u0/u3/_0200_ ;
wire \u0/u3/_0201_ ;
wire \u0/u3/_0202_ ;
wire \u0/u3/_0203_ ;
wire \u0/u3/_0204_ ;
wire \u0/u3/_0205_ ;
wire \u0/u3/_0206_ ;
wire \u0/u3/_0207_ ;
wire \u0/u3/_0208_ ;
wire \u0/u3/_0209_ ;
wire \u0/u3/_0210_ ;
wire \u0/u3/_0211_ ;
wire \u0/u3/_0212_ ;
wire \u0/u3/_0213_ ;
wire \u0/u3/_0214_ ;
wire \u0/u3/_0215_ ;
wire \u0/u3/_0216_ ;
wire \u0/u3/_0217_ ;
wire \u0/u3/_0218_ ;
wire \u0/u3/_0219_ ;
wire \u0/u3/_0220_ ;
wire \u0/u3/_0221_ ;
wire \u0/u3/_0222_ ;
wire \u0/u3/_0223_ ;
wire \u0/u3/_0224_ ;
wire \u0/u3/_0225_ ;
wire \u0/u3/_0226_ ;
wire \u0/u3/_0227_ ;
wire \u0/u3/_0228_ ;
wire \u0/u3/_0229_ ;
wire \u0/u3/_0230_ ;
wire \u0/u3/_0231_ ;
wire \u0/u3/_0232_ ;
wire \u0/u3/_0233_ ;
wire \u0/u3/_0234_ ;
wire \u0/u3/_0235_ ;
wire \u0/u3/_0236_ ;
wire \u0/u3/_0237_ ;
wire \u0/u3/_0238_ ;
wire \u0/u3/_0239_ ;
wire \u0/u3/_0240_ ;
wire \u0/u3/_0241_ ;
wire \u0/u3/_0242_ ;
wire \u0/u3/_0243_ ;
wire \u0/u3/_0244_ ;
wire \u0/u3/_0245_ ;
wire \u0/u3/_0246_ ;
wire \u0/u3/_0248_ ;
wire \u0/u3/_0249_ ;
wire \u0/u3/_0250_ ;
wire \u0/u3/_0251_ ;
wire \u0/u3/_0252_ ;
wire \u0/u3/_0253_ ;
wire \u0/u3/_0254_ ;
wire \u0/u3/_0255_ ;
wire \u0/u3/_0256_ ;
wire \u0/u3/_0257_ ;
wire \u0/u3/_0258_ ;
wire \u0/u3/_0259_ ;
wire \u0/u3/_0260_ ;
wire \u0/u3/_0261_ ;
wire \u0/u3/_0263_ ;
wire \u0/u3/_0264_ ;
wire \u0/u3/_0265_ ;
wire \u0/u3/_0266_ ;
wire \u0/u3/_0267_ ;
wire \u0/u3/_0268_ ;
wire \u0/u3/_0269_ ;
wire \u0/u3/_0270_ ;
wire \u0/u3/_0271_ ;
wire \u0/u3/_0272_ ;
wire \u0/u3/_0273_ ;
wire \u0/u3/_0274_ ;
wire \u0/u3/_0275_ ;
wire \u0/u3/_0276_ ;
wire \u0/u3/_0277_ ;
wire \u0/u3/_0278_ ;
wire \u0/u3/_0279_ ;
wire \u0/u3/_0281_ ;
wire \u0/u3/_0283_ ;
wire \u0/u3/_0284_ ;
wire \u0/u3/_0285_ ;
wire \u0/u3/_0286_ ;
wire \u0/u3/_0287_ ;
wire \u0/u3/_0288_ ;
wire \u0/u3/_0289_ ;
wire \u0/u3/_0290_ ;
wire \u0/u3/_0291_ ;
wire \u0/u3/_0292_ ;
wire \u0/u3/_0293_ ;
wire \u0/u3/_0294_ ;
wire \u0/u3/_0295_ ;
wire \u0/u3/_0296_ ;
wire \u0/u3/_0297_ ;
wire \u0/u3/_0298_ ;
wire \u0/u3/_0299_ ;
wire \u0/u3/_0300_ ;
wire \u0/u3/_0301_ ;
wire \u0/u3/_0302_ ;
wire \u0/u3/_0303_ ;
wire \u0/u3/_0304_ ;
wire \u0/u3/_0305_ ;
wire \u0/u3/_0306_ ;
wire \u0/u3/_0307_ ;
wire \u0/u3/_0308_ ;
wire \u0/u3/_0309_ ;
wire \u0/u3/_0310_ ;
wire \u0/u3/_0311_ ;
wire \u0/u3/_0312_ ;
wire \u0/u3/_0313_ ;
wire \u0/u3/_0314_ ;
wire \u0/u3/_0315_ ;
wire \u0/u3/_0316_ ;
wire \u0/u3/_0317_ ;
wire \u0/u3/_0318_ ;
wire \u0/u3/_0319_ ;
wire \u0/u3/_0320_ ;
wire \u0/u3/_0321_ ;
wire \u0/u3/_0322_ ;
wire \u0/u3/_0323_ ;
wire \u0/u3/_0324_ ;
wire \u0/u3/_0325_ ;
wire \u0/u3/_0326_ ;
wire \u0/u3/_0327_ ;
wire \u0/u3/_0328_ ;
wire \u0/u3/_0329_ ;
wire \u0/u3/_0330_ ;
wire \u0/u3/_0331_ ;
wire \u0/u3/_0332_ ;
wire \u0/u3/_0333_ ;
wire \u0/u3/_0334_ ;
wire \u0/u3/_0335_ ;
wire \u0/u3/_0337_ ;
wire \u0/u3/_0338_ ;
wire \u0/u3/_0339_ ;
wire \u0/u3/_0340_ ;
wire \u0/u3/_0341_ ;
wire \u0/u3/_0342_ ;
wire \u0/u3/_0343_ ;
wire \u0/u3/_0344_ ;
wire \u0/u3/_0345_ ;
wire \u0/u3/_0347_ ;
wire \u0/u3/_0348_ ;
wire \u0/u3/_0349_ ;
wire \u0/u3/_0350_ ;
wire \u0/u3/_0351_ ;
wire \u0/u3/_0352_ ;
wire \u0/u3/_0353_ ;
wire \u0/u3/_0354_ ;
wire \u0/u3/_0355_ ;
wire \u0/u3/_0356_ ;
wire \u0/u3/_0357_ ;
wire \u0/u3/_0358_ ;
wire \u0/u3/_0359_ ;
wire \u0/u3/_0360_ ;
wire \u0/u3/_0361_ ;
wire \u0/u3/_0362_ ;
wire \u0/u3/_0363_ ;
wire \u0/u3/_0364_ ;
wire \u0/u3/_0365_ ;
wire \u0/u3/_0366_ ;
wire \u0/u3/_0367_ ;
wire \u0/u3/_0368_ ;
wire \u0/u3/_0370_ ;
wire \u0/u3/_0371_ ;
wire \u0/u3/_0372_ ;
wire \u0/u3/_0373_ ;
wire \u0/u3/_0374_ ;
wire \u0/u3/_0375_ ;
wire \u0/u3/_0376_ ;
wire \u0/u3/_0377_ ;
wire \u0/u3/_0378_ ;
wire \u0/u3/_0379_ ;
wire \u0/u3/_0380_ ;
wire \u0/u3/_0381_ ;
wire \u0/u3/_0382_ ;
wire \u0/u3/_0383_ ;
wire \u0/u3/_0384_ ;
wire \u0/u3/_0385_ ;
wire \u0/u3/_0386_ ;
wire \u0/u3/_0387_ ;
wire \u0/u3/_0388_ ;
wire \u0/u3/_0389_ ;
wire \u0/u3/_0390_ ;
wire \u0/u3/_0391_ ;
wire \u0/u3/_0392_ ;
wire \u0/u3/_0393_ ;
wire \u0/u3/_0394_ ;
wire \u0/u3/_0395_ ;
wire \u0/u3/_0396_ ;
wire \u0/u3/_0397_ ;
wire \u0/u3/_0398_ ;
wire \u0/u3/_0399_ ;
wire \u0/u3/_0400_ ;
wire \u0/u3/_0401_ ;
wire \u0/u3/_0402_ ;
wire \u0/u3/_0403_ ;
wire \u0/u3/_0404_ ;
wire \u0/u3/_0405_ ;
wire \u0/u3/_0406_ ;
wire \u0/u3/_0407_ ;
wire \u0/u3/_0408_ ;
wire \u0/u3/_0409_ ;
wire \u0/u3/_0410_ ;
wire \u0/u3/_0411_ ;
wire \u0/u3/_0412_ ;
wire \u0/u3/_0413_ ;
wire \u0/u3/_0414_ ;
wire \u0/u3/_0415_ ;
wire \u0/u3/_0416_ ;
wire \u0/u3/_0417_ ;
wire \u0/u3/_0418_ ;
wire \u0/u3/_0419_ ;
wire \u0/u3/_0420_ ;
wire \u0/u3/_0421_ ;
wire \u0/u3/_0422_ ;
wire \u0/u3/_0424_ ;
wire \u0/u3/_0425_ ;
wire \u0/u3/_0426_ ;
wire \u0/u3/_0427_ ;
wire \u0/u3/_0428_ ;
wire \u0/u3/_0429_ ;
wire \u0/u3/_0430_ ;
wire \u0/u3/_0431_ ;
wire \u0/u3/_0432_ ;
wire \u0/u3/_0433_ ;
wire \u0/u3/_0434_ ;
wire \u0/u3/_0435_ ;
wire \u0/u3/_0436_ ;
wire \u0/u3/_0437_ ;
wire \u0/u3/_0438_ ;
wire \u0/u3/_0439_ ;
wire \u0/u3/_0440_ ;
wire \u0/u3/_0441_ ;
wire \u0/u3/_0442_ ;
wire \u0/u3/_0443_ ;
wire \u0/u3/_0444_ ;
wire \u0/u3/_0446_ ;
wire \u0/u3/_0447_ ;
wire \u0/u3/_0448_ ;
wire \u0/u3/_0449_ ;
wire \u0/u3/_0450_ ;
wire \u0/u3/_0451_ ;
wire \u0/u3/_0452_ ;
wire \u0/u3/_0453_ ;
wire \u0/u3/_0454_ ;
wire \u0/u3/_0455_ ;
wire \u0/u3/_0457_ ;
wire \u0/u3/_0458_ ;
wire \u0/u3/_0459_ ;
wire \u0/u3/_0460_ ;
wire \u0/u3/_0461_ ;
wire \u0/u3/_0462_ ;
wire \u0/u3/_0463_ ;
wire \u0/u3/_0464_ ;
wire \u0/u3/_0465_ ;
wire \u0/u3/_0466_ ;
wire \u0/u3/_0467_ ;
wire \u0/u3/_0468_ ;
wire \u0/u3/_0469_ ;
wire \u0/u3/_0470_ ;
wire \u0/u3/_0471_ ;
wire \u0/u3/_0472_ ;
wire \u0/u3/_0473_ ;
wire \u0/u3/_0474_ ;
wire \u0/u3/_0475_ ;
wire \u0/u3/_0476_ ;
wire \u0/u3/_0477_ ;
wire \u0/u3/_0478_ ;
wire \u0/u3/_0479_ ;
wire \u0/u3/_0480_ ;
wire \u0/u3/_0481_ ;
wire \u0/u3/_0482_ ;
wire \u0/u3/_0483_ ;
wire \u0/u3/_0484_ ;
wire \u0/u3/_0485_ ;
wire \u0/u3/_0486_ ;
wire \u0/u3/_0487_ ;
wire \u0/u3/_0488_ ;
wire \u0/u3/_0490_ ;
wire \u0/u3/_0491_ ;
wire \u0/u3/_0492_ ;
wire \u0/u3/_0493_ ;
wire \u0/u3/_0494_ ;
wire \u0/u3/_0495_ ;
wire \u0/u3/_0496_ ;
wire \u0/u3/_0497_ ;
wire \u0/u3/_0498_ ;
wire \u0/u3/_0500_ ;
wire \u0/u3/_0501_ ;
wire \u0/u3/_0502_ ;
wire \u0/u3/_0503_ ;
wire \u0/u3/_0504_ ;
wire \u0/u3/_0505_ ;
wire \u0/u3/_0506_ ;
wire \u0/u3/_0507_ ;
wire \u0/u3/_0508_ ;
wire \u0/u3/_0509_ ;
wire \u0/u3/_0510_ ;
wire \u0/u3/_0511_ ;
wire \u0/u3/_0512_ ;
wire \u0/u3/_0513_ ;
wire \u0/u3/_0514_ ;
wire \u0/u3/_0515_ ;
wire \u0/u3/_0516_ ;
wire \u0/u3/_0517_ ;
wire \u0/u3/_0518_ ;
wire \u0/u3/_0519_ ;
wire \u0/u3/_0520_ ;
wire \u0/u3/_0521_ ;
wire \u0/u3/_0522_ ;
wire \u0/u3/_0523_ ;
wire \u0/u3/_0524_ ;
wire \u0/u3/_0525_ ;
wire \u0/u3/_0526_ ;
wire \u0/u3/_0527_ ;
wire \u0/u3/_0528_ ;
wire \u0/u3/_0529_ ;
wire \u0/u3/_0530_ ;
wire \u0/u3/_0531_ ;
wire \u0/u3/_0532_ ;
wire \u0/u3/_0533_ ;
wire \u0/u3/_0534_ ;
wire \u0/u3/_0535_ ;
wire \u0/u3/_0536_ ;
wire \u0/u3/_0537_ ;
wire \u0/u3/_0538_ ;
wire \u0/u3/_0539_ ;
wire \u0/u3/_0540_ ;
wire \u0/u3/_0541_ ;
wire \u0/u3/_0542_ ;
wire \u0/u3/_0544_ ;
wire \u0/u3/_0545_ ;
wire \u0/u3/_0546_ ;
wire \u0/u3/_0547_ ;
wire \u0/u3/_0548_ ;
wire \u0/u3/_0549_ ;
wire \u0/u3/_0550_ ;
wire \u0/u3/_0551_ ;
wire \u0/u3/_0552_ ;
wire \u0/u3/_0553_ ;
wire \u0/u3/_0554_ ;
wire \u0/u3/_0555_ ;
wire \u0/u3/_0556_ ;
wire \u0/u3/_0557_ ;
wire \u0/u3/_0558_ ;
wire \u0/u3/_0559_ ;
wire \u0/u3/_0560_ ;
wire \u0/u3/_0561_ ;
wire \u0/u3/_0562_ ;
wire \u0/u3/_0563_ ;
wire \u0/u3/_0565_ ;
wire \u0/u3/_0566_ ;
wire \u0/u3/_0567_ ;
wire \u0/u3/_0568_ ;
wire \u0/u3/_0569_ ;
wire \u0/u3/_0570_ ;
wire \u0/u3/_0571_ ;
wire \u0/u3/_0572_ ;
wire \u0/u3/_0573_ ;
wire \u0/u3/_0574_ ;
wire \u0/u3/_0575_ ;
wire \u0/u3/_0576_ ;
wire \u0/u3/_0577_ ;
wire \u0/u3/_0578_ ;
wire \u0/u3/_0579_ ;
wire \u0/u3/_0580_ ;
wire \u0/u3/_0581_ ;
wire \u0/u3/_0582_ ;
wire \u0/u3/_0583_ ;
wire \u0/u3/_0584_ ;
wire \u0/u3/_0585_ ;
wire \u0/u3/_0586_ ;
wire \u0/u3/_0587_ ;
wire \u0/u3/_0588_ ;
wire \u0/u3/_0589_ ;
wire \u0/u3/_0590_ ;
wire \u0/u3/_0591_ ;
wire \u0/u3/_0592_ ;
wire \u0/u3/_0593_ ;
wire \u0/u3/_0594_ ;
wire \u0/u3/_0595_ ;
wire \u0/u3/_0596_ ;
wire \u0/u3/_0598_ ;
wire \u0/u3/_0599_ ;
wire \u0/u3/_0600_ ;
wire \u0/u3/_0601_ ;
wire \u0/u3/_0602_ ;
wire \u0/u3/_0603_ ;
wire \u0/u3/_0604_ ;
wire \u0/u3/_0605_ ;
wire \u0/u3/_0606_ ;
wire \u0/u3/_0607_ ;
wire \u0/u3/_0608_ ;
wire \u0/u3/_0609_ ;
wire \u0/u3/_0610_ ;
wire \u0/u3/_0611_ ;
wire \u0/u3/_0612_ ;
wire \u0/u3/_0613_ ;
wire \u0/u3/_0614_ ;
wire \u0/u3/_0615_ ;
wire \u0/u3/_0616_ ;
wire \u0/u3/_0617_ ;
wire \u0/u3/_0618_ ;
wire \u0/u3/_0619_ ;
wire \u0/u3/_0620_ ;
wire \u0/u3/_0621_ ;
wire \u0/u3/_0622_ ;
wire \u0/u3/_0623_ ;
wire \u0/u3/_0624_ ;
wire \u0/u3/_0625_ ;
wire \u0/u3/_0626_ ;
wire \u0/u3/_0627_ ;
wire \u0/u3/_0628_ ;
wire \u0/u3/_0629_ ;
wire \u0/u3/_0630_ ;
wire \u0/u3/_0631_ ;
wire \u0/u3/_0632_ ;
wire \u0/u3/_0633_ ;
wire \u0/u3/_0634_ ;
wire \u0/u3/_0635_ ;
wire \u0/u3/_0636_ ;
wire \u0/u3/_0637_ ;
wire \u0/u3/_0638_ ;
wire \u0/u3/_0639_ ;
wire \u0/u3/_0640_ ;
wire \u0/u3/_0641_ ;
wire \u0/u3/_0642_ ;
wire \u0/u3/_0643_ ;
wire \u0/u3/_0644_ ;
wire \u0/u3/_0645_ ;
wire \u0/u3/_0646_ ;
wire \u0/u3/_0647_ ;
wire \u0/u3/_0648_ ;
wire \u0/u3/_0649_ ;
wire \u0/u3/_0650_ ;
wire \u0/u3/_0652_ ;
wire \u0/u3/_0653_ ;
wire \u0/u3/_0654_ ;
wire \u0/u3/_0655_ ;
wire \u0/u3/_0656_ ;
wire \u0/u3/_0657_ ;
wire \u0/u3/_0658_ ;
wire \u0/u3/_0659_ ;
wire \u0/u3/_0660_ ;
wire \u0/u3/_0661_ ;
wire \u0/u3/_0662_ ;
wire \u0/u3/_0663_ ;
wire \u0/u3/_0664_ ;
wire \u0/u3/_0665_ ;
wire \u0/u3/_0666_ ;
wire \u0/u3/_0667_ ;
wire \u0/u3/_0668_ ;
wire \u0/u3/_0669_ ;
wire \u0/u3/_0670_ ;
wire \u0/u3/_0671_ ;
wire \u0/u3/_0673_ ;
wire \u0/u3/_0674_ ;
wire \u0/u3/_0675_ ;
wire \u0/u3/_0676_ ;
wire \u0/u3/_0677_ ;
wire \u0/u3/_0678_ ;
wire \u0/u3/_0679_ ;
wire \u0/u3/_0680_ ;
wire \u0/u3/_0681_ ;
wire \u0/u3/_0682_ ;
wire \u0/u3/_0683_ ;
wire \u0/u3/_0684_ ;
wire \u0/u3/_0685_ ;
wire \u0/u3/_0686_ ;
wire \u0/u3/_0687_ ;
wire \u0/u3/_0688_ ;
wire \u0/u3/_0689_ ;
wire \u0/u3/_0690_ ;
wire \u0/u3/_0691_ ;
wire \u0/u3/_0692_ ;
wire \u0/u3/_0693_ ;
wire \u0/u3/_0694_ ;
wire \u0/u3/_0695_ ;
wire \u0/u3/_0696_ ;
wire \u0/u3/_0697_ ;
wire \u0/u3/_0698_ ;
wire \u0/u3/_0699_ ;
wire \u0/u3/_0700_ ;
wire \u0/u3/_0701_ ;
wire \u0/u3/_0702_ ;
wire \u0/u3/_0703_ ;
wire \u0/u3/_0704_ ;
wire \u0/u3/_0705_ ;
wire \u0/u3/_0706_ ;
wire \u0/u3/_0707_ ;
wire \u0/u3/_0708_ ;
wire \u0/u3/_0709_ ;
wire \u0/u3/_0710_ ;
wire \u0/u3/_0711_ ;
wire \u0/u3/_0712_ ;
wire \u0/u3/_0713_ ;
wire \u0/u3/_0714_ ;
wire \u0/u3/_0715_ ;
wire \u0/u3/_0717_ ;
wire \u0/u3/_0718_ ;
wire \u0/u3/_0719_ ;
wire \u0/u3/_0720_ ;
wire \u0/u3/_0721_ ;
wire \u0/u3/_0722_ ;
wire \u0/u3/_0723_ ;
wire \u0/u3/_0724_ ;
wire \u0/u3/_0725_ ;
wire \u0/u3/_0726_ ;
wire \u0/u3/_0727_ ;
wire \u0/u3/_0728_ ;
wire \u0/u3/_0729_ ;
wire \u0/u3/_0730_ ;
wire \u0/u3/_0731_ ;
wire \u0/u3/_0733_ ;
wire \u0/u3/_0734_ ;
wire \u0/u3/_0735_ ;
wire \u0/u3/_0736_ ;
wire \u0/u3/_0738_ ;
wire \u0/u3/_0739_ ;
wire \u0/u3/_0740_ ;
wire \u0/u3/_0741_ ;
wire \u0/u3/_0742_ ;
wire \u0/u3/_0744_ ;
wire \u0/u3/_0745_ ;
wire \u0/u3/_0746_ ;
wire \u0/u3/_0748_ ;
wire \u0/u3/_0749_ ;
wire \u0/u3/_0750_ ;
wire \u0/u3/_0752_ ;
wire \us00/_0008_ ;
wire \us00/_0009_ ;
wire \us00/_0010_ ;
wire \us00/_0011_ ;
wire \us00/_0012_ ;
wire \us00/_0013_ ;
wire \us00/_0014_ ;
wire \us00/_0015_ ;
wire \us00/_0016_ ;
wire \us00/_0017_ ;
wire \us00/_0019_ ;
wire \us00/_0020_ ;
wire \us00/_0022_ ;
wire \us00/_0024_ ;
wire \us00/_0025_ ;
wire \us00/_0026_ ;
wire \us00/_0027_ ;
wire \us00/_0030_ ;
wire \us00/_0032_ ;
wire \us00/_0033_ ;
wire \us00/_0034_ ;
wire \us00/_0035_ ;
wire \us00/_0037_ ;
wire \us00/_0038_ ;
wire \us00/_0039_ ;
wire \us00/_0040_ ;
wire \us00/_0041_ ;
wire \us00/_0042_ ;
wire \us00/_0043_ ;
wire \us00/_0045_ ;
wire \us00/_0046_ ;
wire \us00/_0047_ ;
wire \us00/_0049_ ;
wire \us00/_0050_ ;
wire \us00/_0051_ ;
wire \us00/_0052_ ;
wire \us00/_0053_ ;
wire \us00/_0054_ ;
wire \us00/_0057_ ;
wire \us00/_0058_ ;
wire \us00/_0060_ ;
wire \us00/_0061_ ;
wire \us00/_0062_ ;
wire \us00/_0064_ ;
wire \us00/_0065_ ;
wire \us00/_0066_ ;
wire \us00/_0067_ ;
wire \us00/_0069_ ;
wire \us00/_0070_ ;
wire \us00/_0072_ ;
wire \us00/_0073_ ;
wire \us00/_0074_ ;
wire \us00/_0075_ ;
wire \us00/_0076_ ;
wire \us00/_0077_ ;
wire \us00/_0078_ ;
wire \us00/_0079_ ;
wire \us00/_0081_ ;
wire \us00/_0082_ ;
wire \us00/_0084_ ;
wire \us00/_0085_ ;
wire \us00/_0086_ ;
wire \us00/_0087_ ;
wire \us00/_0088_ ;
wire \us00/_0089_ ;
wire \us00/_0090_ ;
wire \us00/_0091_ ;
wire \us00/_0092_ ;
wire \us00/_0093_ ;
wire \us00/_0094_ ;
wire \us00/_0095_ ;
wire \us00/_0096_ ;
wire \us00/_0097_ ;
wire \us00/_0098_ ;
wire \us00/_0099_ ;
wire \us00/_0100_ ;
wire \us00/_0101_ ;
wire \us00/_0102_ ;
wire \us00/_0103_ ;
wire \us00/_0104_ ;
wire \us00/_0105_ ;
wire \us00/_0106_ ;
wire \us00/_0108_ ;
wire \us00/_0109_ ;
wire \us00/_0110_ ;
wire \us00/_0111_ ;
wire \us00/_0113_ ;
wire \us00/_0114_ ;
wire \us00/_0115_ ;
wire \us00/_0116_ ;
wire \us00/_0117_ ;
wire \us00/_0118_ ;
wire \us00/_0119_ ;
wire \us00/_0120_ ;
wire \us00/_0121_ ;
wire \us00/_0122_ ;
wire \us00/_0123_ ;
wire \us00/_0124_ ;
wire \us00/_0126_ ;
wire \us00/_0127_ ;
wire \us00/_0128_ ;
wire \us00/_0129_ ;
wire \us00/_0130_ ;
wire \us00/_0132_ ;
wire \us00/_0133_ ;
wire \us00/_0134_ ;
wire \us00/_0135_ ;
wire \us00/_0136_ ;
wire \us00/_0137_ ;
wire \us00/_0139_ ;
wire \us00/_0140_ ;
wire \us00/_0141_ ;
wire \us00/_0142_ ;
wire \us00/_0144_ ;
wire \us00/_0145_ ;
wire \us00/_0146_ ;
wire \us00/_0147_ ;
wire \us00/_0148_ ;
wire \us00/_0149_ ;
wire \us00/_0150_ ;
wire \us00/_0151_ ;
wire \us00/_0153_ ;
wire \us00/_0154_ ;
wire \us00/_0155_ ;
wire \us00/_0156_ ;
wire \us00/_0157_ ;
wire \us00/_0158_ ;
wire \us00/_0159_ ;
wire \us00/_0161_ ;
wire \us00/_0162_ ;
wire \us00/_0163_ ;
wire \us00/_0164_ ;
wire \us00/_0165_ ;
wire \us00/_0166_ ;
wire \us00/_0167_ ;
wire \us00/_0168_ ;
wire \us00/_0169_ ;
wire \us00/_0170_ ;
wire \us00/_0171_ ;
wire \us00/_0172_ ;
wire \us00/_0174_ ;
wire \us00/_0175_ ;
wire \us00/_0176_ ;
wire \us00/_0177_ ;
wire \us00/_0178_ ;
wire \us00/_0179_ ;
wire \us00/_0180_ ;
wire \us00/_0181_ ;
wire \us00/_0182_ ;
wire \us00/_0183_ ;
wire \us00/_0184_ ;
wire \us00/_0185_ ;
wire \us00/_0186_ ;
wire \us00/_0187_ ;
wire \us00/_0188_ ;
wire \us00/_0189_ ;
wire \us00/_0190_ ;
wire \us00/_0191_ ;
wire \us00/_0192_ ;
wire \us00/_0193_ ;
wire \us00/_0194_ ;
wire \us00/_0195_ ;
wire \us00/_0196_ ;
wire \us00/_0197_ ;
wire \us00/_0198_ ;
wire \us00/_0199_ ;
wire \us00/_0200_ ;
wire \us00/_0201_ ;
wire \us00/_0202_ ;
wire \us00/_0203_ ;
wire \us00/_0204_ ;
wire \us00/_0205_ ;
wire \us00/_0206_ ;
wire \us00/_0207_ ;
wire \us00/_0208_ ;
wire \us00/_0209_ ;
wire \us00/_0210_ ;
wire \us00/_0211_ ;
wire \us00/_0212_ ;
wire \us00/_0213_ ;
wire \us00/_0214_ ;
wire \us00/_0215_ ;
wire \us00/_0217_ ;
wire \us00/_0218_ ;
wire \us00/_0219_ ;
wire \us00/_0220_ ;
wire \us00/_0221_ ;
wire \us00/_0222_ ;
wire \us00/_0223_ ;
wire \us00/_0224_ ;
wire \us00/_0225_ ;
wire \us00/_0226_ ;
wire \us00/_0227_ ;
wire \us00/_0228_ ;
wire \us00/_0229_ ;
wire \us00/_0230_ ;
wire \us00/_0231_ ;
wire \us00/_0232_ ;
wire \us00/_0233_ ;
wire \us00/_0234_ ;
wire \us00/_0235_ ;
wire \us00/_0236_ ;
wire \us00/_0237_ ;
wire \us00/_0238_ ;
wire \us00/_0239_ ;
wire \us00/_0240_ ;
wire \us00/_0241_ ;
wire \us00/_0242_ ;
wire \us00/_0243_ ;
wire \us00/_0244_ ;
wire \us00/_0245_ ;
wire \us00/_0246_ ;
wire \us00/_0247_ ;
wire \us00/_0248_ ;
wire \us00/_0249_ ;
wire \us00/_0250_ ;
wire \us00/_0251_ ;
wire \us00/_0252_ ;
wire \us00/_0253_ ;
wire \us00/_0254_ ;
wire \us00/_0255_ ;
wire \us00/_0256_ ;
wire \us00/_0257_ ;
wire \us00/_0258_ ;
wire \us00/_0259_ ;
wire \us00/_0260_ ;
wire \us00/_0261_ ;
wire \us00/_0263_ ;
wire \us00/_0264_ ;
wire \us00/_0265_ ;
wire \us00/_0266_ ;
wire \us00/_0267_ ;
wire \us00/_0268_ ;
wire \us00/_0269_ ;
wire \us00/_0270_ ;
wire \us00/_0271_ ;
wire \us00/_0272_ ;
wire \us00/_0273_ ;
wire \us00/_0274_ ;
wire \us00/_0275_ ;
wire \us00/_0276_ ;
wire \us00/_0277_ ;
wire \us00/_0278_ ;
wire \us00/_0279_ ;
wire \us00/_0281_ ;
wire \us00/_0283_ ;
wire \us00/_0284_ ;
wire \us00/_0285_ ;
wire \us00/_0286_ ;
wire \us00/_0287_ ;
wire \us00/_0288_ ;
wire \us00/_0289_ ;
wire \us00/_0290_ ;
wire \us00/_0291_ ;
wire \us00/_0292_ ;
wire \us00/_0293_ ;
wire \us00/_0294_ ;
wire \us00/_0295_ ;
wire \us00/_0296_ ;
wire \us00/_0297_ ;
wire \us00/_0298_ ;
wire \us00/_0299_ ;
wire \us00/_0300_ ;
wire \us00/_0301_ ;
wire \us00/_0302_ ;
wire \us00/_0303_ ;
wire \us00/_0304_ ;
wire \us00/_0305_ ;
wire \us00/_0306_ ;
wire \us00/_0307_ ;
wire \us00/_0308_ ;
wire \us00/_0309_ ;
wire \us00/_0310_ ;
wire \us00/_0311_ ;
wire \us00/_0312_ ;
wire \us00/_0313_ ;
wire \us00/_0314_ ;
wire \us00/_0315_ ;
wire \us00/_0316_ ;
wire \us00/_0317_ ;
wire \us00/_0318_ ;
wire \us00/_0319_ ;
wire \us00/_0320_ ;
wire \us00/_0321_ ;
wire \us00/_0322_ ;
wire \us00/_0323_ ;
wire \us00/_0324_ ;
wire \us00/_0325_ ;
wire \us00/_0326_ ;
wire \us00/_0327_ ;
wire \us00/_0328_ ;
wire \us00/_0329_ ;
wire \us00/_0330_ ;
wire \us00/_0331_ ;
wire \us00/_0332_ ;
wire \us00/_0333_ ;
wire \us00/_0334_ ;
wire \us00/_0335_ ;
wire \us00/_0337_ ;
wire \us00/_0338_ ;
wire \us00/_0339_ ;
wire \us00/_0340_ ;
wire \us00/_0341_ ;
wire \us00/_0342_ ;
wire \us00/_0343_ ;
wire \us00/_0344_ ;
wire \us00/_0345_ ;
wire \us00/_0347_ ;
wire \us00/_0348_ ;
wire \us00/_0349_ ;
wire \us00/_0350_ ;
wire \us00/_0351_ ;
wire \us00/_0352_ ;
wire \us00/_0353_ ;
wire \us00/_0354_ ;
wire \us00/_0355_ ;
wire \us00/_0356_ ;
wire \us00/_0357_ ;
wire \us00/_0358_ ;
wire \us00/_0359_ ;
wire \us00/_0360_ ;
wire \us00/_0361_ ;
wire \us00/_0362_ ;
wire \us00/_0363_ ;
wire \us00/_0365_ ;
wire \us00/_0366_ ;
wire \us00/_0367_ ;
wire \us00/_0368_ ;
wire \us00/_0370_ ;
wire \us00/_0371_ ;
wire \us00/_0372_ ;
wire \us00/_0373_ ;
wire \us00/_0374_ ;
wire \us00/_0375_ ;
wire \us00/_0376_ ;
wire \us00/_0377_ ;
wire \us00/_0378_ ;
wire \us00/_0379_ ;
wire \us00/_0380_ ;
wire \us00/_0381_ ;
wire \us00/_0382_ ;
wire \us00/_0383_ ;
wire \us00/_0384_ ;
wire \us00/_0385_ ;
wire \us00/_0386_ ;
wire \us00/_0387_ ;
wire \us00/_0388_ ;
wire \us00/_0389_ ;
wire \us00/_0390_ ;
wire \us00/_0391_ ;
wire \us00/_0392_ ;
wire \us00/_0393_ ;
wire \us00/_0394_ ;
wire \us00/_0395_ ;
wire \us00/_0396_ ;
wire \us00/_0397_ ;
wire \us00/_0398_ ;
wire \us00/_0399_ ;
wire \us00/_0400_ ;
wire \us00/_0401_ ;
wire \us00/_0402_ ;
wire \us00/_0403_ ;
wire \us00/_0404_ ;
wire \us00/_0405_ ;
wire \us00/_0406_ ;
wire \us00/_0407_ ;
wire \us00/_0408_ ;
wire \us00/_0409_ ;
wire \us00/_0410_ ;
wire \us00/_0411_ ;
wire \us00/_0412_ ;
wire \us00/_0413_ ;
wire \us00/_0414_ ;
wire \us00/_0415_ ;
wire \us00/_0416_ ;
wire \us00/_0417_ ;
wire \us00/_0418_ ;
wire \us00/_0419_ ;
wire \us00/_0420_ ;
wire \us00/_0421_ ;
wire \us00/_0422_ ;
wire \us00/_0424_ ;
wire \us00/_0425_ ;
wire \us00/_0426_ ;
wire \us00/_0427_ ;
wire \us00/_0428_ ;
wire \us00/_0429_ ;
wire \us00/_0430_ ;
wire \us00/_0431_ ;
wire \us00/_0432_ ;
wire \us00/_0433_ ;
wire \us00/_0434_ ;
wire \us00/_0435_ ;
wire \us00/_0436_ ;
wire \us00/_0437_ ;
wire \us00/_0438_ ;
wire \us00/_0439_ ;
wire \us00/_0440_ ;
wire \us00/_0441_ ;
wire \us00/_0442_ ;
wire \us00/_0443_ ;
wire \us00/_0444_ ;
wire \us00/_0446_ ;
wire \us00/_0447_ ;
wire \us00/_0448_ ;
wire \us00/_0449_ ;
wire \us00/_0450_ ;
wire \us00/_0451_ ;
wire \us00/_0452_ ;
wire \us00/_0453_ ;
wire \us00/_0454_ ;
wire \us00/_0455_ ;
wire \us00/_0457_ ;
wire \us00/_0458_ ;
wire \us00/_0459_ ;
wire \us00/_0460_ ;
wire \us00/_0461_ ;
wire \us00/_0462_ ;
wire \us00/_0463_ ;
wire \us00/_0464_ ;
wire \us00/_0465_ ;
wire \us00/_0466_ ;
wire \us00/_0467_ ;
wire \us00/_0468_ ;
wire \us00/_0469_ ;
wire \us00/_0470_ ;
wire \us00/_0471_ ;
wire \us00/_0472_ ;
wire \us00/_0473_ ;
wire \us00/_0474_ ;
wire \us00/_0475_ ;
wire \us00/_0476_ ;
wire \us00/_0477_ ;
wire \us00/_0478_ ;
wire \us00/_0479_ ;
wire \us00/_0480_ ;
wire \us00/_0481_ ;
wire \us00/_0482_ ;
wire \us00/_0483_ ;
wire \us00/_0484_ ;
wire \us00/_0485_ ;
wire \us00/_0486_ ;
wire \us00/_0487_ ;
wire \us00/_0488_ ;
wire \us00/_0490_ ;
wire \us00/_0491_ ;
wire \us00/_0492_ ;
wire \us00/_0493_ ;
wire \us00/_0494_ ;
wire \us00/_0495_ ;
wire \us00/_0496_ ;
wire \us00/_0497_ ;
wire \us00/_0498_ ;
wire \us00/_0500_ ;
wire \us00/_0501_ ;
wire \us00/_0502_ ;
wire \us00/_0503_ ;
wire \us00/_0504_ ;
wire \us00/_0505_ ;
wire \us00/_0506_ ;
wire \us00/_0507_ ;
wire \us00/_0508_ ;
wire \us00/_0509_ ;
wire \us00/_0510_ ;
wire \us00/_0511_ ;
wire \us00/_0512_ ;
wire \us00/_0513_ ;
wire \us00/_0514_ ;
wire \us00/_0515_ ;
wire \us00/_0516_ ;
wire \us00/_0517_ ;
wire \us00/_0518_ ;
wire \us00/_0519_ ;
wire \us00/_0520_ ;
wire \us00/_0521_ ;
wire \us00/_0522_ ;
wire \us00/_0523_ ;
wire \us00/_0524_ ;
wire \us00/_0525_ ;
wire \us00/_0526_ ;
wire \us00/_0527_ ;
wire \us00/_0528_ ;
wire \us00/_0529_ ;
wire \us00/_0530_ ;
wire \us00/_0531_ ;
wire \us00/_0532_ ;
wire \us00/_0533_ ;
wire \us00/_0534_ ;
wire \us00/_0535_ ;
wire \us00/_0536_ ;
wire \us00/_0537_ ;
wire \us00/_0538_ ;
wire \us00/_0539_ ;
wire \us00/_0540_ ;
wire \us00/_0541_ ;
wire \us00/_0542_ ;
wire \us00/_0544_ ;
wire \us00/_0545_ ;
wire \us00/_0546_ ;
wire \us00/_0547_ ;
wire \us00/_0548_ ;
wire \us00/_0549_ ;
wire \us00/_0550_ ;
wire \us00/_0551_ ;
wire \us00/_0552_ ;
wire \us00/_0553_ ;
wire \us00/_0554_ ;
wire \us00/_0555_ ;
wire \us00/_0556_ ;
wire \us00/_0557_ ;
wire \us00/_0558_ ;
wire \us00/_0559_ ;
wire \us00/_0560_ ;
wire \us00/_0561_ ;
wire \us00/_0562_ ;
wire \us00/_0563_ ;
wire \us00/_0565_ ;
wire \us00/_0566_ ;
wire \us00/_0567_ ;
wire \us00/_0568_ ;
wire \us00/_0569_ ;
wire \us00/_0570_ ;
wire \us00/_0571_ ;
wire \us00/_0572_ ;
wire \us00/_0573_ ;
wire \us00/_0574_ ;
wire \us00/_0575_ ;
wire \us00/_0576_ ;
wire \us00/_0577_ ;
wire \us00/_0578_ ;
wire \us00/_0579_ ;
wire \us00/_0580_ ;
wire \us00/_0581_ ;
wire \us00/_0582_ ;
wire \us00/_0583_ ;
wire \us00/_0584_ ;
wire \us00/_0585_ ;
wire \us00/_0586_ ;
wire \us00/_0587_ ;
wire \us00/_0588_ ;
wire \us00/_0589_ ;
wire \us00/_0590_ ;
wire \us00/_0591_ ;
wire \us00/_0592_ ;
wire \us00/_0593_ ;
wire \us00/_0594_ ;
wire \us00/_0595_ ;
wire \us00/_0596_ ;
wire \us00/_0598_ ;
wire \us00/_0599_ ;
wire \us00/_0600_ ;
wire \us00/_0601_ ;
wire \us00/_0602_ ;
wire \us00/_0603_ ;
wire \us00/_0604_ ;
wire \us00/_0605_ ;
wire \us00/_0606_ ;
wire \us00/_0607_ ;
wire \us00/_0608_ ;
wire \us00/_0609_ ;
wire \us00/_0610_ ;
wire \us00/_0611_ ;
wire \us00/_0612_ ;
wire \us00/_0613_ ;
wire \us00/_0614_ ;
wire \us00/_0615_ ;
wire \us00/_0616_ ;
wire \us00/_0617_ ;
wire \us00/_0618_ ;
wire \us00/_0619_ ;
wire \us00/_0620_ ;
wire \us00/_0621_ ;
wire \us00/_0622_ ;
wire \us00/_0623_ ;
wire \us00/_0624_ ;
wire \us00/_0625_ ;
wire \us00/_0626_ ;
wire \us00/_0627_ ;
wire \us00/_0628_ ;
wire \us00/_0629_ ;
wire \us00/_0630_ ;
wire \us00/_0631_ ;
wire \us00/_0632_ ;
wire \us00/_0633_ ;
wire \us00/_0634_ ;
wire \us00/_0635_ ;
wire \us00/_0636_ ;
wire \us00/_0637_ ;
wire \us00/_0638_ ;
wire \us00/_0639_ ;
wire \us00/_0640_ ;
wire \us00/_0641_ ;
wire \us00/_0642_ ;
wire \us00/_0643_ ;
wire \us00/_0644_ ;
wire \us00/_0645_ ;
wire \us00/_0646_ ;
wire \us00/_0647_ ;
wire \us00/_0648_ ;
wire \us00/_0649_ ;
wire \us00/_0650_ ;
wire \us00/_0652_ ;
wire \us00/_0653_ ;
wire \us00/_0654_ ;
wire \us00/_0655_ ;
wire \us00/_0656_ ;
wire \us00/_0657_ ;
wire \us00/_0658_ ;
wire \us00/_0659_ ;
wire \us00/_0660_ ;
wire \us00/_0661_ ;
wire \us00/_0662_ ;
wire \us00/_0663_ ;
wire \us00/_0664_ ;
wire \us00/_0665_ ;
wire \us00/_0666_ ;
wire \us00/_0667_ ;
wire \us00/_0668_ ;
wire \us00/_0669_ ;
wire \us00/_0670_ ;
wire \us00/_0671_ ;
wire \us00/_0673_ ;
wire \us00/_0674_ ;
wire \us00/_0675_ ;
wire \us00/_0676_ ;
wire \us00/_0677_ ;
wire \us00/_0678_ ;
wire \us00/_0679_ ;
wire \us00/_0680_ ;
wire \us00/_0681_ ;
wire \us00/_0682_ ;
wire \us00/_0683_ ;
wire \us00/_0684_ ;
wire \us00/_0685_ ;
wire \us00/_0686_ ;
wire \us00/_0687_ ;
wire \us00/_0688_ ;
wire \us00/_0689_ ;
wire \us00/_0690_ ;
wire \us00/_0691_ ;
wire \us00/_0692_ ;
wire \us00/_0693_ ;
wire \us00/_0694_ ;
wire \us00/_0695_ ;
wire \us00/_0696_ ;
wire \us00/_0697_ ;
wire \us00/_0698_ ;
wire \us00/_0699_ ;
wire \us00/_0700_ ;
wire \us00/_0701_ ;
wire \us00/_0702_ ;
wire \us00/_0703_ ;
wire \us00/_0704_ ;
wire \us00/_0705_ ;
wire \us00/_0706_ ;
wire \us00/_0707_ ;
wire \us00/_0708_ ;
wire \us00/_0709_ ;
wire \us00/_0710_ ;
wire \us00/_0711_ ;
wire \us00/_0712_ ;
wire \us00/_0713_ ;
wire \us00/_0714_ ;
wire \us00/_0715_ ;
wire \us00/_0717_ ;
wire \us00/_0718_ ;
wire \us00/_0719_ ;
wire \us00/_0720_ ;
wire \us00/_0721_ ;
wire \us00/_0722_ ;
wire \us00/_0723_ ;
wire \us00/_0724_ ;
wire \us00/_0725_ ;
wire \us00/_0726_ ;
wire \us00/_0727_ ;
wire \us00/_0728_ ;
wire \us00/_0729_ ;
wire \us00/_0730_ ;
wire \us00/_0731_ ;
wire \us00/_0732_ ;
wire \us00/_0733_ ;
wire \us00/_0734_ ;
wire \us00/_0735_ ;
wire \us00/_0736_ ;
wire \us00/_0738_ ;
wire \us00/_0739_ ;
wire \us00/_0740_ ;
wire \us00/_0741_ ;
wire \us00/_0742_ ;
wire \us00/_0744_ ;
wire \us00/_0745_ ;
wire \us00/_0746_ ;
wire \us00/_0747_ ;
wire \us00/_0748_ ;
wire \us00/_0749_ ;
wire \us00/_0750_ ;
wire \us00/_0752_ ;
wire \us01/_0008_ ;
wire \us01/_0009_ ;
wire \us01/_0010_ ;
wire \us01/_0011_ ;
wire \us01/_0012_ ;
wire \us01/_0013_ ;
wire \us01/_0014_ ;
wire \us01/_0015_ ;
wire \us01/_0016_ ;
wire \us01/_0017_ ;
wire \us01/_0019_ ;
wire \us01/_0020_ ;
wire \us01/_0022_ ;
wire \us01/_0024_ ;
wire \us01/_0025_ ;
wire \us01/_0026_ ;
wire \us01/_0027_ ;
wire \us01/_0029_ ;
wire \us01/_0030_ ;
wire \us01/_0033_ ;
wire \us01/_0034_ ;
wire \us01/_0035_ ;
wire \us01/_0037_ ;
wire \us01/_0038_ ;
wire \us01/_0039_ ;
wire \us01/_0040_ ;
wire \us01/_0041_ ;
wire \us01/_0042_ ;
wire \us01/_0043_ ;
wire \us01/_0045_ ;
wire \us01/_0046_ ;
wire \us01/_0047_ ;
wire \us01/_0049_ ;
wire \us01/_0050_ ;
wire \us01/_0051_ ;
wire \us01/_0052_ ;
wire \us01/_0053_ ;
wire \us01/_0054_ ;
wire \us01/_0057_ ;
wire \us01/_0058_ ;
wire \us01/_0060_ ;
wire \us01/_0061_ ;
wire \us01/_0062_ ;
wire \us01/_0064_ ;
wire \us01/_0065_ ;
wire \us01/_0066_ ;
wire \us01/_0067_ ;
wire \us01/_0069_ ;
wire \us01/_0070_ ;
wire \us01/_0072_ ;
wire \us01/_0073_ ;
wire \us01/_0074_ ;
wire \us01/_0075_ ;
wire \us01/_0076_ ;
wire \us01/_0077_ ;
wire \us01/_0078_ ;
wire \us01/_0079_ ;
wire \us01/_0081_ ;
wire \us01/_0082_ ;
wire \us01/_0085_ ;
wire \us01/_0086_ ;
wire \us01/_0087_ ;
wire \us01/_0088_ ;
wire \us01/_0089_ ;
wire \us01/_0090_ ;
wire \us01/_0091_ ;
wire \us01/_0092_ ;
wire \us01/_0093_ ;
wire \us01/_0094_ ;
wire \us01/_0095_ ;
wire \us01/_0096_ ;
wire \us01/_0097_ ;
wire \us01/_0098_ ;
wire \us01/_0099_ ;
wire \us01/_0100_ ;
wire \us01/_0101_ ;
wire \us01/_0102_ ;
wire \us01/_0103_ ;
wire \us01/_0104_ ;
wire \us01/_0105_ ;
wire \us01/_0106_ ;
wire \us01/_0108_ ;
wire \us01/_0109_ ;
wire \us01/_0110_ ;
wire \us01/_0111_ ;
wire \us01/_0113_ ;
wire \us01/_0114_ ;
wire \us01/_0115_ ;
wire \us01/_0116_ ;
wire \us01/_0117_ ;
wire \us01/_0118_ ;
wire \us01/_0119_ ;
wire \us01/_0120_ ;
wire \us01/_0121_ ;
wire \us01/_0122_ ;
wire \us01/_0123_ ;
wire \us01/_0124_ ;
wire \us01/_0126_ ;
wire \us01/_0127_ ;
wire \us01/_0128_ ;
wire \us01/_0129_ ;
wire \us01/_0130_ ;
wire \us01/_0132_ ;
wire \us01/_0133_ ;
wire \us01/_0134_ ;
wire \us01/_0135_ ;
wire \us01/_0136_ ;
wire \us01/_0137_ ;
wire \us01/_0139_ ;
wire \us01/_0140_ ;
wire \us01/_0141_ ;
wire \us01/_0142_ ;
wire \us01/_0144_ ;
wire \us01/_0145_ ;
wire \us01/_0146_ ;
wire \us01/_0147_ ;
wire \us01/_0148_ ;
wire \us01/_0149_ ;
wire \us01/_0150_ ;
wire \us01/_0151_ ;
wire \us01/_0153_ ;
wire \us01/_0154_ ;
wire \us01/_0155_ ;
wire \us01/_0156_ ;
wire \us01/_0157_ ;
wire \us01/_0158_ ;
wire \us01/_0159_ ;
wire \us01/_0161_ ;
wire \us01/_0162_ ;
wire \us01/_0163_ ;
wire \us01/_0164_ ;
wire \us01/_0165_ ;
wire \us01/_0166_ ;
wire \us01/_0167_ ;
wire \us01/_0168_ ;
wire \us01/_0169_ ;
wire \us01/_0170_ ;
wire \us01/_0171_ ;
wire \us01/_0172_ ;
wire \us01/_0174_ ;
wire \us01/_0175_ ;
wire \us01/_0176_ ;
wire \us01/_0177_ ;
wire \us01/_0178_ ;
wire \us01/_0179_ ;
wire \us01/_0180_ ;
wire \us01/_0181_ ;
wire \us01/_0182_ ;
wire \us01/_0183_ ;
wire \us01/_0184_ ;
wire \us01/_0185_ ;
wire \us01/_0186_ ;
wire \us01/_0187_ ;
wire \us01/_0188_ ;
wire \us01/_0189_ ;
wire \us01/_0190_ ;
wire \us01/_0191_ ;
wire \us01/_0192_ ;
wire \us01/_0193_ ;
wire \us01/_0194_ ;
wire \us01/_0195_ ;
wire \us01/_0196_ ;
wire \us01/_0197_ ;
wire \us01/_0198_ ;
wire \us01/_0199_ ;
wire \us01/_0200_ ;
wire \us01/_0201_ ;
wire \us01/_0202_ ;
wire \us01/_0203_ ;
wire \us01/_0204_ ;
wire \us01/_0205_ ;
wire \us01/_0206_ ;
wire \us01/_0207_ ;
wire \us01/_0208_ ;
wire \us01/_0209_ ;
wire \us01/_0210_ ;
wire \us01/_0211_ ;
wire \us01/_0212_ ;
wire \us01/_0213_ ;
wire \us01/_0214_ ;
wire \us01/_0215_ ;
wire \us01/_0217_ ;
wire \us01/_0218_ ;
wire \us01/_0219_ ;
wire \us01/_0220_ ;
wire \us01/_0221_ ;
wire \us01/_0222_ ;
wire \us01/_0223_ ;
wire \us01/_0224_ ;
wire \us01/_0225_ ;
wire \us01/_0226_ ;
wire \us01/_0227_ ;
wire \us01/_0228_ ;
wire \us01/_0229_ ;
wire \us01/_0230_ ;
wire \us01/_0231_ ;
wire \us01/_0232_ ;
wire \us01/_0233_ ;
wire \us01/_0234_ ;
wire \us01/_0235_ ;
wire \us01/_0236_ ;
wire \us01/_0237_ ;
wire \us01/_0238_ ;
wire \us01/_0239_ ;
wire \us01/_0240_ ;
wire \us01/_0241_ ;
wire \us01/_0242_ ;
wire \us01/_0243_ ;
wire \us01/_0244_ ;
wire \us01/_0245_ ;
wire \us01/_0246_ ;
wire \us01/_0248_ ;
wire \us01/_0249_ ;
wire \us01/_0250_ ;
wire \us01/_0251_ ;
wire \us01/_0252_ ;
wire \us01/_0253_ ;
wire \us01/_0254_ ;
wire \us01/_0255_ ;
wire \us01/_0256_ ;
wire \us01/_0257_ ;
wire \us01/_0258_ ;
wire \us01/_0259_ ;
wire \us01/_0260_ ;
wire \us01/_0261_ ;
wire \us01/_0263_ ;
wire \us01/_0264_ ;
wire \us01/_0265_ ;
wire \us01/_0266_ ;
wire \us01/_0267_ ;
wire \us01/_0268_ ;
wire \us01/_0269_ ;
wire \us01/_0270_ ;
wire \us01/_0271_ ;
wire \us01/_0272_ ;
wire \us01/_0273_ ;
wire \us01/_0274_ ;
wire \us01/_0275_ ;
wire \us01/_0276_ ;
wire \us01/_0277_ ;
wire \us01/_0278_ ;
wire \us01/_0279_ ;
wire \us01/_0280_ ;
wire \us01/_0281_ ;
wire \us01/_0283_ ;
wire \us01/_0284_ ;
wire \us01/_0285_ ;
wire \us01/_0286_ ;
wire \us01/_0287_ ;
wire \us01/_0288_ ;
wire \us01/_0289_ ;
wire \us01/_0290_ ;
wire \us01/_0291_ ;
wire \us01/_0292_ ;
wire \us01/_0293_ ;
wire \us01/_0294_ ;
wire \us01/_0295_ ;
wire \us01/_0296_ ;
wire \us01/_0297_ ;
wire \us01/_0298_ ;
wire \us01/_0299_ ;
wire \us01/_0300_ ;
wire \us01/_0301_ ;
wire \us01/_0302_ ;
wire \us01/_0303_ ;
wire \us01/_0304_ ;
wire \us01/_0305_ ;
wire \us01/_0306_ ;
wire \us01/_0307_ ;
wire \us01/_0308_ ;
wire \us01/_0309_ ;
wire \us01/_0310_ ;
wire \us01/_0311_ ;
wire \us01/_0312_ ;
wire \us01/_0313_ ;
wire \us01/_0314_ ;
wire \us01/_0315_ ;
wire \us01/_0316_ ;
wire \us01/_0317_ ;
wire \us01/_0318_ ;
wire \us01/_0319_ ;
wire \us01/_0320_ ;
wire \us01/_0321_ ;
wire \us01/_0322_ ;
wire \us01/_0323_ ;
wire \us01/_0324_ ;
wire \us01/_0325_ ;
wire \us01/_0326_ ;
wire \us01/_0327_ ;
wire \us01/_0328_ ;
wire \us01/_0329_ ;
wire \us01/_0330_ ;
wire \us01/_0331_ ;
wire \us01/_0332_ ;
wire \us01/_0333_ ;
wire \us01/_0334_ ;
wire \us01/_0335_ ;
wire \us01/_0337_ ;
wire \us01/_0338_ ;
wire \us01/_0339_ ;
wire \us01/_0340_ ;
wire \us01/_0341_ ;
wire \us01/_0342_ ;
wire \us01/_0343_ ;
wire \us01/_0344_ ;
wire \us01/_0345_ ;
wire \us01/_0347_ ;
wire \us01/_0348_ ;
wire \us01/_0349_ ;
wire \us01/_0350_ ;
wire \us01/_0351_ ;
wire \us01/_0352_ ;
wire \us01/_0353_ ;
wire \us01/_0354_ ;
wire \us01/_0355_ ;
wire \us01/_0356_ ;
wire \us01/_0357_ ;
wire \us01/_0358_ ;
wire \us01/_0359_ ;
wire \us01/_0360_ ;
wire \us01/_0361_ ;
wire \us01/_0362_ ;
wire \us01/_0363_ ;
wire \us01/_0365_ ;
wire \us01/_0366_ ;
wire \us01/_0367_ ;
wire \us01/_0368_ ;
wire \us01/_0370_ ;
wire \us01/_0371_ ;
wire \us01/_0372_ ;
wire \us01/_0373_ ;
wire \us01/_0374_ ;
wire \us01/_0375_ ;
wire \us01/_0376_ ;
wire \us01/_0377_ ;
wire \us01/_0378_ ;
wire \us01/_0379_ ;
wire \us01/_0380_ ;
wire \us01/_0381_ ;
wire \us01/_0382_ ;
wire \us01/_0383_ ;
wire \us01/_0384_ ;
wire \us01/_0385_ ;
wire \us01/_0386_ ;
wire \us01/_0387_ ;
wire \us01/_0388_ ;
wire \us01/_0389_ ;
wire \us01/_0390_ ;
wire \us01/_0391_ ;
wire \us01/_0392_ ;
wire \us01/_0393_ ;
wire \us01/_0394_ ;
wire \us01/_0395_ ;
wire \us01/_0396_ ;
wire \us01/_0397_ ;
wire \us01/_0398_ ;
wire \us01/_0399_ ;
wire \us01/_0400_ ;
wire \us01/_0401_ ;
wire \us01/_0402_ ;
wire \us01/_0403_ ;
wire \us01/_0404_ ;
wire \us01/_0405_ ;
wire \us01/_0406_ ;
wire \us01/_0407_ ;
wire \us01/_0408_ ;
wire \us01/_0409_ ;
wire \us01/_0410_ ;
wire \us01/_0411_ ;
wire \us01/_0412_ ;
wire \us01/_0413_ ;
wire \us01/_0414_ ;
wire \us01/_0415_ ;
wire \us01/_0416_ ;
wire \us01/_0417_ ;
wire \us01/_0418_ ;
wire \us01/_0419_ ;
wire \us01/_0420_ ;
wire \us01/_0421_ ;
wire \us01/_0422_ ;
wire \us01/_0424_ ;
wire \us01/_0425_ ;
wire \us01/_0426_ ;
wire \us01/_0427_ ;
wire \us01/_0428_ ;
wire \us01/_0429_ ;
wire \us01/_0430_ ;
wire \us01/_0431_ ;
wire \us01/_0432_ ;
wire \us01/_0433_ ;
wire \us01/_0434_ ;
wire \us01/_0435_ ;
wire \us01/_0436_ ;
wire \us01/_0437_ ;
wire \us01/_0438_ ;
wire \us01/_0439_ ;
wire \us01/_0440_ ;
wire \us01/_0441_ ;
wire \us01/_0442_ ;
wire \us01/_0443_ ;
wire \us01/_0444_ ;
wire \us01/_0446_ ;
wire \us01/_0447_ ;
wire \us01/_0448_ ;
wire \us01/_0449_ ;
wire \us01/_0450_ ;
wire \us01/_0451_ ;
wire \us01/_0452_ ;
wire \us01/_0453_ ;
wire \us01/_0454_ ;
wire \us01/_0455_ ;
wire \us01/_0457_ ;
wire \us01/_0458_ ;
wire \us01/_0459_ ;
wire \us01/_0460_ ;
wire \us01/_0461_ ;
wire \us01/_0462_ ;
wire \us01/_0463_ ;
wire \us01/_0464_ ;
wire \us01/_0465_ ;
wire \us01/_0466_ ;
wire \us01/_0467_ ;
wire \us01/_0468_ ;
wire \us01/_0469_ ;
wire \us01/_0470_ ;
wire \us01/_0471_ ;
wire \us01/_0472_ ;
wire \us01/_0473_ ;
wire \us01/_0474_ ;
wire \us01/_0475_ ;
wire \us01/_0476_ ;
wire \us01/_0477_ ;
wire \us01/_0478_ ;
wire \us01/_0479_ ;
wire \us01/_0480_ ;
wire \us01/_0481_ ;
wire \us01/_0482_ ;
wire \us01/_0483_ ;
wire \us01/_0484_ ;
wire \us01/_0485_ ;
wire \us01/_0486_ ;
wire \us01/_0487_ ;
wire \us01/_0488_ ;
wire \us01/_0490_ ;
wire \us01/_0491_ ;
wire \us01/_0492_ ;
wire \us01/_0493_ ;
wire \us01/_0494_ ;
wire \us01/_0495_ ;
wire \us01/_0496_ ;
wire \us01/_0497_ ;
wire \us01/_0498_ ;
wire \us01/_0500_ ;
wire \us01/_0501_ ;
wire \us01/_0502_ ;
wire \us01/_0503_ ;
wire \us01/_0504_ ;
wire \us01/_0505_ ;
wire \us01/_0506_ ;
wire \us01/_0507_ ;
wire \us01/_0508_ ;
wire \us01/_0509_ ;
wire \us01/_0510_ ;
wire \us01/_0511_ ;
wire \us01/_0512_ ;
wire \us01/_0513_ ;
wire \us01/_0514_ ;
wire \us01/_0515_ ;
wire \us01/_0516_ ;
wire \us01/_0517_ ;
wire \us01/_0518_ ;
wire \us01/_0519_ ;
wire \us01/_0520_ ;
wire \us01/_0521_ ;
wire \us01/_0522_ ;
wire \us01/_0523_ ;
wire \us01/_0524_ ;
wire \us01/_0525_ ;
wire \us01/_0526_ ;
wire \us01/_0527_ ;
wire \us01/_0528_ ;
wire \us01/_0529_ ;
wire \us01/_0530_ ;
wire \us01/_0531_ ;
wire \us01/_0532_ ;
wire \us01/_0533_ ;
wire \us01/_0534_ ;
wire \us01/_0535_ ;
wire \us01/_0536_ ;
wire \us01/_0537_ ;
wire \us01/_0538_ ;
wire \us01/_0539_ ;
wire \us01/_0540_ ;
wire \us01/_0541_ ;
wire \us01/_0542_ ;
wire \us01/_0544_ ;
wire \us01/_0545_ ;
wire \us01/_0546_ ;
wire \us01/_0547_ ;
wire \us01/_0548_ ;
wire \us01/_0549_ ;
wire \us01/_0550_ ;
wire \us01/_0551_ ;
wire \us01/_0552_ ;
wire \us01/_0553_ ;
wire \us01/_0554_ ;
wire \us01/_0555_ ;
wire \us01/_0556_ ;
wire \us01/_0557_ ;
wire \us01/_0558_ ;
wire \us01/_0559_ ;
wire \us01/_0560_ ;
wire \us01/_0561_ ;
wire \us01/_0562_ ;
wire \us01/_0563_ ;
wire \us01/_0565_ ;
wire \us01/_0566_ ;
wire \us01/_0567_ ;
wire \us01/_0568_ ;
wire \us01/_0569_ ;
wire \us01/_0570_ ;
wire \us01/_0571_ ;
wire \us01/_0572_ ;
wire \us01/_0573_ ;
wire \us01/_0574_ ;
wire \us01/_0575_ ;
wire \us01/_0576_ ;
wire \us01/_0577_ ;
wire \us01/_0578_ ;
wire \us01/_0579_ ;
wire \us01/_0580_ ;
wire \us01/_0581_ ;
wire \us01/_0582_ ;
wire \us01/_0583_ ;
wire \us01/_0584_ ;
wire \us01/_0585_ ;
wire \us01/_0586_ ;
wire \us01/_0587_ ;
wire \us01/_0588_ ;
wire \us01/_0589_ ;
wire \us01/_0590_ ;
wire \us01/_0591_ ;
wire \us01/_0592_ ;
wire \us01/_0593_ ;
wire \us01/_0594_ ;
wire \us01/_0595_ ;
wire \us01/_0596_ ;
wire \us01/_0598_ ;
wire \us01/_0599_ ;
wire \us01/_0600_ ;
wire \us01/_0601_ ;
wire \us01/_0602_ ;
wire \us01/_0603_ ;
wire \us01/_0604_ ;
wire \us01/_0605_ ;
wire \us01/_0606_ ;
wire \us01/_0607_ ;
wire \us01/_0608_ ;
wire \us01/_0609_ ;
wire \us01/_0610_ ;
wire \us01/_0611_ ;
wire \us01/_0612_ ;
wire \us01/_0613_ ;
wire \us01/_0614_ ;
wire \us01/_0615_ ;
wire \us01/_0616_ ;
wire \us01/_0617_ ;
wire \us01/_0618_ ;
wire \us01/_0619_ ;
wire \us01/_0620_ ;
wire \us01/_0621_ ;
wire \us01/_0622_ ;
wire \us01/_0623_ ;
wire \us01/_0624_ ;
wire \us01/_0625_ ;
wire \us01/_0626_ ;
wire \us01/_0627_ ;
wire \us01/_0628_ ;
wire \us01/_0629_ ;
wire \us01/_0630_ ;
wire \us01/_0631_ ;
wire \us01/_0632_ ;
wire \us01/_0633_ ;
wire \us01/_0634_ ;
wire \us01/_0635_ ;
wire \us01/_0636_ ;
wire \us01/_0637_ ;
wire \us01/_0638_ ;
wire \us01/_0639_ ;
wire \us01/_0640_ ;
wire \us01/_0641_ ;
wire \us01/_0642_ ;
wire \us01/_0643_ ;
wire \us01/_0644_ ;
wire \us01/_0645_ ;
wire \us01/_0646_ ;
wire \us01/_0647_ ;
wire \us01/_0648_ ;
wire \us01/_0649_ ;
wire \us01/_0650_ ;
wire \us01/_0652_ ;
wire \us01/_0653_ ;
wire \us01/_0654_ ;
wire \us01/_0655_ ;
wire \us01/_0656_ ;
wire \us01/_0657_ ;
wire \us01/_0658_ ;
wire \us01/_0659_ ;
wire \us01/_0660_ ;
wire \us01/_0661_ ;
wire \us01/_0662_ ;
wire \us01/_0663_ ;
wire \us01/_0664_ ;
wire \us01/_0665_ ;
wire \us01/_0666_ ;
wire \us01/_0667_ ;
wire \us01/_0668_ ;
wire \us01/_0669_ ;
wire \us01/_0670_ ;
wire \us01/_0671_ ;
wire \us01/_0673_ ;
wire \us01/_0674_ ;
wire \us01/_0675_ ;
wire \us01/_0676_ ;
wire \us01/_0677_ ;
wire \us01/_0678_ ;
wire \us01/_0679_ ;
wire \us01/_0680_ ;
wire \us01/_0681_ ;
wire \us01/_0682_ ;
wire \us01/_0683_ ;
wire \us01/_0684_ ;
wire \us01/_0685_ ;
wire \us01/_0686_ ;
wire \us01/_0687_ ;
wire \us01/_0688_ ;
wire \us01/_0689_ ;
wire \us01/_0690_ ;
wire \us01/_0691_ ;
wire \us01/_0692_ ;
wire \us01/_0693_ ;
wire \us01/_0694_ ;
wire \us01/_0695_ ;
wire \us01/_0696_ ;
wire \us01/_0697_ ;
wire \us01/_0698_ ;
wire \us01/_0699_ ;
wire \us01/_0700_ ;
wire \us01/_0701_ ;
wire \us01/_0702_ ;
wire \us01/_0703_ ;
wire \us01/_0704_ ;
wire \us01/_0705_ ;
wire \us01/_0706_ ;
wire \us01/_0707_ ;
wire \us01/_0708_ ;
wire \us01/_0709_ ;
wire \us01/_0710_ ;
wire \us01/_0711_ ;
wire \us01/_0712_ ;
wire \us01/_0713_ ;
wire \us01/_0714_ ;
wire \us01/_0715_ ;
wire \us01/_0717_ ;
wire \us01/_0718_ ;
wire \us01/_0719_ ;
wire \us01/_0720_ ;
wire \us01/_0721_ ;
wire \us01/_0722_ ;
wire \us01/_0723_ ;
wire \us01/_0724_ ;
wire \us01/_0725_ ;
wire \us01/_0726_ ;
wire \us01/_0727_ ;
wire \us01/_0728_ ;
wire \us01/_0729_ ;
wire \us01/_0730_ ;
wire \us01/_0731_ ;
wire \us01/_0733_ ;
wire \us01/_0734_ ;
wire \us01/_0735_ ;
wire \us01/_0736_ ;
wire \us01/_0738_ ;
wire \us01/_0739_ ;
wire \us01/_0740_ ;
wire \us01/_0741_ ;
wire \us01/_0742_ ;
wire \us01/_0744_ ;
wire \us01/_0745_ ;
wire \us01/_0746_ ;
wire \us01/_0748_ ;
wire \us01/_0749_ ;
wire \us01/_0750_ ;
wire \us01/_0752_ ;
wire \us02/_0008_ ;
wire \us02/_0009_ ;
wire \us02/_0010_ ;
wire \us02/_0011_ ;
wire \us02/_0012_ ;
wire \us02/_0013_ ;
wire \us02/_0014_ ;
wire \us02/_0015_ ;
wire \us02/_0016_ ;
wire \us02/_0017_ ;
wire \us02/_0019_ ;
wire \us02/_0020_ ;
wire \us02/_0022_ ;
wire \us02/_0024_ ;
wire \us02/_0025_ ;
wire \us02/_0026_ ;
wire \us02/_0027_ ;
wire \us02/_0030_ ;
wire \us02/_0032_ ;
wire \us02/_0033_ ;
wire \us02/_0034_ ;
wire \us02/_0035_ ;
wire \us02/_0037_ ;
wire \us02/_0038_ ;
wire \us02/_0039_ ;
wire \us02/_0040_ ;
wire \us02/_0041_ ;
wire \us02/_0042_ ;
wire \us02/_0043_ ;
wire \us02/_0045_ ;
wire \us02/_0046_ ;
wire \us02/_0047_ ;
wire \us02/_0049_ ;
wire \us02/_0050_ ;
wire \us02/_0051_ ;
wire \us02/_0052_ ;
wire \us02/_0053_ ;
wire \us02/_0054_ ;
wire \us02/_0056_ ;
wire \us02/_0057_ ;
wire \us02/_0058_ ;
wire \us02/_0060_ ;
wire \us02/_0061_ ;
wire \us02/_0062_ ;
wire \us02/_0064_ ;
wire \us02/_0065_ ;
wire \us02/_0066_ ;
wire \us02/_0067_ ;
wire \us02/_0069_ ;
wire \us02/_0070_ ;
wire \us02/_0072_ ;
wire \us02/_0073_ ;
wire \us02/_0074_ ;
wire \us02/_0075_ ;
wire \us02/_0076_ ;
wire \us02/_0077_ ;
wire \us02/_0078_ ;
wire \us02/_0079_ ;
wire \us02/_0081_ ;
wire \us02/_0082_ ;
wire \us02/_0084_ ;
wire \us02/_0085_ ;
wire \us02/_0086_ ;
wire \us02/_0087_ ;
wire \us02/_0088_ ;
wire \us02/_0089_ ;
wire \us02/_0090_ ;
wire \us02/_0091_ ;
wire \us02/_0092_ ;
wire \us02/_0093_ ;
wire \us02/_0094_ ;
wire \us02/_0095_ ;
wire \us02/_0096_ ;
wire \us02/_0097_ ;
wire \us02/_0098_ ;
wire \us02/_0099_ ;
wire \us02/_0100_ ;
wire \us02/_0101_ ;
wire \us02/_0102_ ;
wire \us02/_0103_ ;
wire \us02/_0104_ ;
wire \us02/_0105_ ;
wire \us02/_0106_ ;
wire \us02/_0108_ ;
wire \us02/_0109_ ;
wire \us02/_0110_ ;
wire \us02/_0111_ ;
wire \us02/_0113_ ;
wire \us02/_0114_ ;
wire \us02/_0115_ ;
wire \us02/_0116_ ;
wire \us02/_0117_ ;
wire \us02/_0118_ ;
wire \us02/_0119_ ;
wire \us02/_0120_ ;
wire \us02/_0121_ ;
wire \us02/_0122_ ;
wire \us02/_0123_ ;
wire \us02/_0124_ ;
wire \us02/_0126_ ;
wire \us02/_0127_ ;
wire \us02/_0128_ ;
wire \us02/_0129_ ;
wire \us02/_0130_ ;
wire \us02/_0132_ ;
wire \us02/_0133_ ;
wire \us02/_0134_ ;
wire \us02/_0135_ ;
wire \us02/_0136_ ;
wire \us02/_0137_ ;
wire \us02/_0139_ ;
wire \us02/_0140_ ;
wire \us02/_0141_ ;
wire \us02/_0142_ ;
wire \us02/_0144_ ;
wire \us02/_0145_ ;
wire \us02/_0146_ ;
wire \us02/_0147_ ;
wire \us02/_0148_ ;
wire \us02/_0149_ ;
wire \us02/_0150_ ;
wire \us02/_0151_ ;
wire \us02/_0153_ ;
wire \us02/_0154_ ;
wire \us02/_0155_ ;
wire \us02/_0156_ ;
wire \us02/_0157_ ;
wire \us02/_0158_ ;
wire \us02/_0159_ ;
wire \us02/_0161_ ;
wire \us02/_0162_ ;
wire \us02/_0163_ ;
wire \us02/_0164_ ;
wire \us02/_0165_ ;
wire \us02/_0166_ ;
wire \us02/_0167_ ;
wire \us02/_0168_ ;
wire \us02/_0169_ ;
wire \us02/_0170_ ;
wire \us02/_0171_ ;
wire \us02/_0172_ ;
wire \us02/_0174_ ;
wire \us02/_0175_ ;
wire \us02/_0176_ ;
wire \us02/_0177_ ;
wire \us02/_0178_ ;
wire \us02/_0179_ ;
wire \us02/_0180_ ;
wire \us02/_0181_ ;
wire \us02/_0182_ ;
wire \us02/_0183_ ;
wire \us02/_0184_ ;
wire \us02/_0185_ ;
wire \us02/_0186_ ;
wire \us02/_0187_ ;
wire \us02/_0188_ ;
wire \us02/_0189_ ;
wire \us02/_0190_ ;
wire \us02/_0191_ ;
wire \us02/_0192_ ;
wire \us02/_0193_ ;
wire \us02/_0194_ ;
wire \us02/_0195_ ;
wire \us02/_0196_ ;
wire \us02/_0197_ ;
wire \us02/_0198_ ;
wire \us02/_0199_ ;
wire \us02/_0200_ ;
wire \us02/_0201_ ;
wire \us02/_0202_ ;
wire \us02/_0203_ ;
wire \us02/_0204_ ;
wire \us02/_0205_ ;
wire \us02/_0206_ ;
wire \us02/_0207_ ;
wire \us02/_0208_ ;
wire \us02/_0209_ ;
wire \us02/_0210_ ;
wire \us02/_0211_ ;
wire \us02/_0212_ ;
wire \us02/_0213_ ;
wire \us02/_0214_ ;
wire \us02/_0215_ ;
wire \us02/_0217_ ;
wire \us02/_0218_ ;
wire \us02/_0219_ ;
wire \us02/_0220_ ;
wire \us02/_0221_ ;
wire \us02/_0222_ ;
wire \us02/_0223_ ;
wire \us02/_0224_ ;
wire \us02/_0225_ ;
wire \us02/_0226_ ;
wire \us02/_0227_ ;
wire \us02/_0228_ ;
wire \us02/_0229_ ;
wire \us02/_0230_ ;
wire \us02/_0231_ ;
wire \us02/_0232_ ;
wire \us02/_0233_ ;
wire \us02/_0234_ ;
wire \us02/_0235_ ;
wire \us02/_0236_ ;
wire \us02/_0237_ ;
wire \us02/_0238_ ;
wire \us02/_0239_ ;
wire \us02/_0240_ ;
wire \us02/_0241_ ;
wire \us02/_0242_ ;
wire \us02/_0243_ ;
wire \us02/_0244_ ;
wire \us02/_0245_ ;
wire \us02/_0246_ ;
wire \us02/_0247_ ;
wire \us02/_0248_ ;
wire \us02/_0249_ ;
wire \us02/_0250_ ;
wire \us02/_0251_ ;
wire \us02/_0252_ ;
wire \us02/_0253_ ;
wire \us02/_0254_ ;
wire \us02/_0255_ ;
wire \us02/_0256_ ;
wire \us02/_0257_ ;
wire \us02/_0258_ ;
wire \us02/_0259_ ;
wire \us02/_0260_ ;
wire \us02/_0261_ ;
wire \us02/_0263_ ;
wire \us02/_0264_ ;
wire \us02/_0265_ ;
wire \us02/_0266_ ;
wire \us02/_0267_ ;
wire \us02/_0268_ ;
wire \us02/_0269_ ;
wire \us02/_0270_ ;
wire \us02/_0271_ ;
wire \us02/_0272_ ;
wire \us02/_0273_ ;
wire \us02/_0274_ ;
wire \us02/_0275_ ;
wire \us02/_0276_ ;
wire \us02/_0277_ ;
wire \us02/_0278_ ;
wire \us02/_0279_ ;
wire \us02/_0281_ ;
wire \us02/_0283_ ;
wire \us02/_0284_ ;
wire \us02/_0285_ ;
wire \us02/_0286_ ;
wire \us02/_0287_ ;
wire \us02/_0288_ ;
wire \us02/_0289_ ;
wire \us02/_0290_ ;
wire \us02/_0291_ ;
wire \us02/_0293_ ;
wire \us02/_0294_ ;
wire \us02/_0295_ ;
wire \us02/_0296_ ;
wire \us02/_0297_ ;
wire \us02/_0298_ ;
wire \us02/_0299_ ;
wire \us02/_0300_ ;
wire \us02/_0301_ ;
wire \us02/_0302_ ;
wire \us02/_0303_ ;
wire \us02/_0304_ ;
wire \us02/_0305_ ;
wire \us02/_0306_ ;
wire \us02/_0307_ ;
wire \us02/_0308_ ;
wire \us02/_0309_ ;
wire \us02/_0310_ ;
wire \us02/_0311_ ;
wire \us02/_0312_ ;
wire \us02/_0313_ ;
wire \us02/_0314_ ;
wire \us02/_0315_ ;
wire \us02/_0316_ ;
wire \us02/_0317_ ;
wire \us02/_0318_ ;
wire \us02/_0319_ ;
wire \us02/_0320_ ;
wire \us02/_0321_ ;
wire \us02/_0322_ ;
wire \us02/_0323_ ;
wire \us02/_0324_ ;
wire \us02/_0325_ ;
wire \us02/_0326_ ;
wire \us02/_0327_ ;
wire \us02/_0328_ ;
wire \us02/_0329_ ;
wire \us02/_0330_ ;
wire \us02/_0331_ ;
wire \us02/_0332_ ;
wire \us02/_0333_ ;
wire \us02/_0334_ ;
wire \us02/_0335_ ;
wire \us02/_0337_ ;
wire \us02/_0338_ ;
wire \us02/_0339_ ;
wire \us02/_0340_ ;
wire \us02/_0341_ ;
wire \us02/_0342_ ;
wire \us02/_0343_ ;
wire \us02/_0344_ ;
wire \us02/_0345_ ;
wire \us02/_0347_ ;
wire \us02/_0348_ ;
wire \us02/_0349_ ;
wire \us02/_0350_ ;
wire \us02/_0351_ ;
wire \us02/_0352_ ;
wire \us02/_0353_ ;
wire \us02/_0354_ ;
wire \us02/_0355_ ;
wire \us02/_0356_ ;
wire \us02/_0357_ ;
wire \us02/_0358_ ;
wire \us02/_0359_ ;
wire \us02/_0360_ ;
wire \us02/_0361_ ;
wire \us02/_0362_ ;
wire \us02/_0363_ ;
wire \us02/_0365_ ;
wire \us02/_0366_ ;
wire \us02/_0367_ ;
wire \us02/_0368_ ;
wire \us02/_0370_ ;
wire \us02/_0371_ ;
wire \us02/_0372_ ;
wire \us02/_0373_ ;
wire \us02/_0374_ ;
wire \us02/_0375_ ;
wire \us02/_0376_ ;
wire \us02/_0377_ ;
wire \us02/_0378_ ;
wire \us02/_0379_ ;
wire \us02/_0380_ ;
wire \us02/_0381_ ;
wire \us02/_0382_ ;
wire \us02/_0383_ ;
wire \us02/_0384_ ;
wire \us02/_0385_ ;
wire \us02/_0386_ ;
wire \us02/_0387_ ;
wire \us02/_0388_ ;
wire \us02/_0389_ ;
wire \us02/_0390_ ;
wire \us02/_0391_ ;
wire \us02/_0392_ ;
wire \us02/_0393_ ;
wire \us02/_0394_ ;
wire \us02/_0395_ ;
wire \us02/_0396_ ;
wire \us02/_0397_ ;
wire \us02/_0398_ ;
wire \us02/_0399_ ;
wire \us02/_0400_ ;
wire \us02/_0401_ ;
wire \us02/_0402_ ;
wire \us02/_0403_ ;
wire \us02/_0404_ ;
wire \us02/_0405_ ;
wire \us02/_0406_ ;
wire \us02/_0407_ ;
wire \us02/_0408_ ;
wire \us02/_0409_ ;
wire \us02/_0410_ ;
wire \us02/_0411_ ;
wire \us02/_0412_ ;
wire \us02/_0413_ ;
wire \us02/_0414_ ;
wire \us02/_0415_ ;
wire \us02/_0416_ ;
wire \us02/_0417_ ;
wire \us02/_0418_ ;
wire \us02/_0419_ ;
wire \us02/_0420_ ;
wire \us02/_0421_ ;
wire \us02/_0422_ ;
wire \us02/_0424_ ;
wire \us02/_0425_ ;
wire \us02/_0426_ ;
wire \us02/_0427_ ;
wire \us02/_0428_ ;
wire \us02/_0429_ ;
wire \us02/_0430_ ;
wire \us02/_0431_ ;
wire \us02/_0432_ ;
wire \us02/_0433_ ;
wire \us02/_0434_ ;
wire \us02/_0435_ ;
wire \us02/_0436_ ;
wire \us02/_0437_ ;
wire \us02/_0438_ ;
wire \us02/_0439_ ;
wire \us02/_0440_ ;
wire \us02/_0441_ ;
wire \us02/_0442_ ;
wire \us02/_0443_ ;
wire \us02/_0444_ ;
wire \us02/_0446_ ;
wire \us02/_0447_ ;
wire \us02/_0448_ ;
wire \us02/_0449_ ;
wire \us02/_0450_ ;
wire \us02/_0451_ ;
wire \us02/_0452_ ;
wire \us02/_0453_ ;
wire \us02/_0454_ ;
wire \us02/_0455_ ;
wire \us02/_0457_ ;
wire \us02/_0458_ ;
wire \us02/_0459_ ;
wire \us02/_0460_ ;
wire \us02/_0461_ ;
wire \us02/_0462_ ;
wire \us02/_0463_ ;
wire \us02/_0464_ ;
wire \us02/_0465_ ;
wire \us02/_0466_ ;
wire \us02/_0467_ ;
wire \us02/_0468_ ;
wire \us02/_0469_ ;
wire \us02/_0470_ ;
wire \us02/_0471_ ;
wire \us02/_0472_ ;
wire \us02/_0473_ ;
wire \us02/_0474_ ;
wire \us02/_0475_ ;
wire \us02/_0476_ ;
wire \us02/_0477_ ;
wire \us02/_0478_ ;
wire \us02/_0479_ ;
wire \us02/_0480_ ;
wire \us02/_0481_ ;
wire \us02/_0482_ ;
wire \us02/_0483_ ;
wire \us02/_0484_ ;
wire \us02/_0485_ ;
wire \us02/_0486_ ;
wire \us02/_0487_ ;
wire \us02/_0488_ ;
wire \us02/_0490_ ;
wire \us02/_0491_ ;
wire \us02/_0492_ ;
wire \us02/_0493_ ;
wire \us02/_0494_ ;
wire \us02/_0495_ ;
wire \us02/_0496_ ;
wire \us02/_0497_ ;
wire \us02/_0498_ ;
wire \us02/_0500_ ;
wire \us02/_0501_ ;
wire \us02/_0502_ ;
wire \us02/_0503_ ;
wire \us02/_0504_ ;
wire \us02/_0505_ ;
wire \us02/_0506_ ;
wire \us02/_0507_ ;
wire \us02/_0508_ ;
wire \us02/_0509_ ;
wire \us02/_0510_ ;
wire \us02/_0511_ ;
wire \us02/_0512_ ;
wire \us02/_0513_ ;
wire \us02/_0514_ ;
wire \us02/_0515_ ;
wire \us02/_0516_ ;
wire \us02/_0517_ ;
wire \us02/_0518_ ;
wire \us02/_0519_ ;
wire \us02/_0520_ ;
wire \us02/_0521_ ;
wire \us02/_0522_ ;
wire \us02/_0523_ ;
wire \us02/_0524_ ;
wire \us02/_0525_ ;
wire \us02/_0526_ ;
wire \us02/_0527_ ;
wire \us02/_0528_ ;
wire \us02/_0529_ ;
wire \us02/_0530_ ;
wire \us02/_0531_ ;
wire \us02/_0532_ ;
wire \us02/_0533_ ;
wire \us02/_0534_ ;
wire \us02/_0535_ ;
wire \us02/_0536_ ;
wire \us02/_0537_ ;
wire \us02/_0538_ ;
wire \us02/_0539_ ;
wire \us02/_0540_ ;
wire \us02/_0541_ ;
wire \us02/_0542_ ;
wire \us02/_0544_ ;
wire \us02/_0545_ ;
wire \us02/_0546_ ;
wire \us02/_0547_ ;
wire \us02/_0548_ ;
wire \us02/_0549_ ;
wire \us02/_0550_ ;
wire \us02/_0551_ ;
wire \us02/_0552_ ;
wire \us02/_0553_ ;
wire \us02/_0554_ ;
wire \us02/_0555_ ;
wire \us02/_0556_ ;
wire \us02/_0557_ ;
wire \us02/_0558_ ;
wire \us02/_0559_ ;
wire \us02/_0560_ ;
wire \us02/_0561_ ;
wire \us02/_0562_ ;
wire \us02/_0563_ ;
wire \us02/_0565_ ;
wire \us02/_0566_ ;
wire \us02/_0567_ ;
wire \us02/_0568_ ;
wire \us02/_0569_ ;
wire \us02/_0570_ ;
wire \us02/_0571_ ;
wire \us02/_0572_ ;
wire \us02/_0573_ ;
wire \us02/_0574_ ;
wire \us02/_0575_ ;
wire \us02/_0576_ ;
wire \us02/_0577_ ;
wire \us02/_0578_ ;
wire \us02/_0579_ ;
wire \us02/_0580_ ;
wire \us02/_0581_ ;
wire \us02/_0582_ ;
wire \us02/_0583_ ;
wire \us02/_0584_ ;
wire \us02/_0585_ ;
wire \us02/_0586_ ;
wire \us02/_0587_ ;
wire \us02/_0588_ ;
wire \us02/_0589_ ;
wire \us02/_0590_ ;
wire \us02/_0591_ ;
wire \us02/_0592_ ;
wire \us02/_0593_ ;
wire \us02/_0594_ ;
wire \us02/_0595_ ;
wire \us02/_0596_ ;
wire \us02/_0598_ ;
wire \us02/_0599_ ;
wire \us02/_0600_ ;
wire \us02/_0601_ ;
wire \us02/_0602_ ;
wire \us02/_0603_ ;
wire \us02/_0604_ ;
wire \us02/_0605_ ;
wire \us02/_0606_ ;
wire \us02/_0607_ ;
wire \us02/_0608_ ;
wire \us02/_0609_ ;
wire \us02/_0610_ ;
wire \us02/_0611_ ;
wire \us02/_0612_ ;
wire \us02/_0613_ ;
wire \us02/_0614_ ;
wire \us02/_0615_ ;
wire \us02/_0616_ ;
wire \us02/_0617_ ;
wire \us02/_0618_ ;
wire \us02/_0619_ ;
wire \us02/_0620_ ;
wire \us02/_0621_ ;
wire \us02/_0622_ ;
wire \us02/_0623_ ;
wire \us02/_0624_ ;
wire \us02/_0625_ ;
wire \us02/_0626_ ;
wire \us02/_0627_ ;
wire \us02/_0628_ ;
wire \us02/_0629_ ;
wire \us02/_0630_ ;
wire \us02/_0631_ ;
wire \us02/_0632_ ;
wire \us02/_0633_ ;
wire \us02/_0634_ ;
wire \us02/_0635_ ;
wire \us02/_0636_ ;
wire \us02/_0637_ ;
wire \us02/_0638_ ;
wire \us02/_0639_ ;
wire \us02/_0640_ ;
wire \us02/_0641_ ;
wire \us02/_0642_ ;
wire \us02/_0643_ ;
wire \us02/_0644_ ;
wire \us02/_0645_ ;
wire \us02/_0646_ ;
wire \us02/_0647_ ;
wire \us02/_0648_ ;
wire \us02/_0649_ ;
wire \us02/_0650_ ;
wire \us02/_0652_ ;
wire \us02/_0653_ ;
wire \us02/_0654_ ;
wire \us02/_0655_ ;
wire \us02/_0656_ ;
wire \us02/_0657_ ;
wire \us02/_0658_ ;
wire \us02/_0659_ ;
wire \us02/_0660_ ;
wire \us02/_0661_ ;
wire \us02/_0662_ ;
wire \us02/_0663_ ;
wire \us02/_0664_ ;
wire \us02/_0665_ ;
wire \us02/_0666_ ;
wire \us02/_0667_ ;
wire \us02/_0668_ ;
wire \us02/_0669_ ;
wire \us02/_0670_ ;
wire \us02/_0671_ ;
wire \us02/_0673_ ;
wire \us02/_0674_ ;
wire \us02/_0675_ ;
wire \us02/_0676_ ;
wire \us02/_0677_ ;
wire \us02/_0678_ ;
wire \us02/_0679_ ;
wire \us02/_0680_ ;
wire \us02/_0681_ ;
wire \us02/_0682_ ;
wire \us02/_0683_ ;
wire \us02/_0684_ ;
wire \us02/_0685_ ;
wire \us02/_0686_ ;
wire \us02/_0687_ ;
wire \us02/_0688_ ;
wire \us02/_0689_ ;
wire \us02/_0690_ ;
wire \us02/_0691_ ;
wire \us02/_0692_ ;
wire \us02/_0693_ ;
wire \us02/_0694_ ;
wire \us02/_0695_ ;
wire \us02/_0696_ ;
wire \us02/_0697_ ;
wire \us02/_0698_ ;
wire \us02/_0699_ ;
wire \us02/_0700_ ;
wire \us02/_0701_ ;
wire \us02/_0702_ ;
wire \us02/_0703_ ;
wire \us02/_0704_ ;
wire \us02/_0705_ ;
wire \us02/_0706_ ;
wire \us02/_0707_ ;
wire \us02/_0708_ ;
wire \us02/_0709_ ;
wire \us02/_0710_ ;
wire \us02/_0711_ ;
wire \us02/_0712_ ;
wire \us02/_0713_ ;
wire \us02/_0714_ ;
wire \us02/_0715_ ;
wire \us02/_0717_ ;
wire \us02/_0718_ ;
wire \us02/_0719_ ;
wire \us02/_0720_ ;
wire \us02/_0721_ ;
wire \us02/_0722_ ;
wire \us02/_0723_ ;
wire \us02/_0724_ ;
wire \us02/_0725_ ;
wire \us02/_0726_ ;
wire \us02/_0727_ ;
wire \us02/_0728_ ;
wire \us02/_0729_ ;
wire \us02/_0730_ ;
wire \us02/_0731_ ;
wire \us02/_0733_ ;
wire \us02/_0734_ ;
wire \us02/_0735_ ;
wire \us02/_0736_ ;
wire \us02/_0738_ ;
wire \us02/_0739_ ;
wire \us02/_0740_ ;
wire \us02/_0741_ ;
wire \us02/_0742_ ;
wire \us02/_0744_ ;
wire \us02/_0745_ ;
wire \us02/_0746_ ;
wire \us02/_0748_ ;
wire \us02/_0749_ ;
wire \us02/_0750_ ;
wire \us02/_0752_ ;
wire \us03/_0008_ ;
wire \us03/_0009_ ;
wire \us03/_0010_ ;
wire \us03/_0011_ ;
wire \us03/_0012_ ;
wire \us03/_0013_ ;
wire \us03/_0014_ ;
wire \us03/_0015_ ;
wire \us03/_0016_ ;
wire \us03/_0017_ ;
wire \us03/_0018_ ;
wire \us03/_0019_ ;
wire \us03/_0020_ ;
wire \us03/_0022_ ;
wire \us03/_0024_ ;
wire \us03/_0025_ ;
wire \us03/_0026_ ;
wire \us03/_0027_ ;
wire \us03/_0028_ ;
wire \us03/_0030_ ;
wire \us03/_0032_ ;
wire \us03/_0033_ ;
wire \us03/_0034_ ;
wire \us03/_0035_ ;
wire \us03/_0036_ ;
wire \us03/_0037_ ;
wire \us03/_0038_ ;
wire \us03/_0039_ ;
wire \us03/_0040_ ;
wire \us03/_0041_ ;
wire \us03/_0042_ ;
wire \us03/_0043_ ;
wire \us03/_0045_ ;
wire \us03/_0046_ ;
wire \us03/_0047_ ;
wire \us03/_0048_ ;
wire \us03/_0049_ ;
wire \us03/_0050_ ;
wire \us03/_0051_ ;
wire \us03/_0052_ ;
wire \us03/_0053_ ;
wire \us03/_0054_ ;
wire \us03/_0056_ ;
wire \us03/_0057_ ;
wire \us03/_0058_ ;
wire \us03/_0060_ ;
wire \us03/_0061_ ;
wire \us03/_0062_ ;
wire \us03/_0064_ ;
wire \us03/_0065_ ;
wire \us03/_0066_ ;
wire \us03/_0067_ ;
wire \us03/_0069_ ;
wire \us03/_0070_ ;
wire \us03/_0072_ ;
wire \us03/_0073_ ;
wire \us03/_0074_ ;
wire \us03/_0075_ ;
wire \us03/_0076_ ;
wire \us03/_0077_ ;
wire \us03/_0078_ ;
wire \us03/_0079_ ;
wire \us03/_0081_ ;
wire \us03/_0082_ ;
wire \us03/_0085_ ;
wire \us03/_0086_ ;
wire \us03/_0087_ ;
wire \us03/_0088_ ;
wire \us03/_0089_ ;
wire \us03/_0090_ ;
wire \us03/_0091_ ;
wire \us03/_0092_ ;
wire \us03/_0093_ ;
wire \us03/_0094_ ;
wire \us03/_0095_ ;
wire \us03/_0096_ ;
wire \us03/_0097_ ;
wire \us03/_0098_ ;
wire \us03/_0100_ ;
wire \us03/_0101_ ;
wire \us03/_0102_ ;
wire \us03/_0103_ ;
wire \us03/_0104_ ;
wire \us03/_0105_ ;
wire \us03/_0106_ ;
wire \us03/_0108_ ;
wire \us03/_0109_ ;
wire \us03/_0110_ ;
wire \us03/_0111_ ;
wire \us03/_0113_ ;
wire \us03/_0114_ ;
wire \us03/_0115_ ;
wire \us03/_0116_ ;
wire \us03/_0117_ ;
wire \us03/_0118_ ;
wire \us03/_0119_ ;
wire \us03/_0120_ ;
wire \us03/_0121_ ;
wire \us03/_0122_ ;
wire \us03/_0123_ ;
wire \us03/_0124_ ;
wire \us03/_0126_ ;
wire \us03/_0127_ ;
wire \us03/_0128_ ;
wire \us03/_0129_ ;
wire \us03/_0130_ ;
wire \us03/_0132_ ;
wire \us03/_0133_ ;
wire \us03/_0134_ ;
wire \us03/_0135_ ;
wire \us03/_0136_ ;
wire \us03/_0137_ ;
wire \us03/_0139_ ;
wire \us03/_0140_ ;
wire \us03/_0141_ ;
wire \us03/_0142_ ;
wire \us03/_0144_ ;
wire \us03/_0145_ ;
wire \us03/_0146_ ;
wire \us03/_0147_ ;
wire \us03/_0148_ ;
wire \us03/_0149_ ;
wire \us03/_0150_ ;
wire \us03/_0151_ ;
wire \us03/_0153_ ;
wire \us03/_0154_ ;
wire \us03/_0155_ ;
wire \us03/_0156_ ;
wire \us03/_0157_ ;
wire \us03/_0158_ ;
wire \us03/_0159_ ;
wire \us03/_0161_ ;
wire \us03/_0162_ ;
wire \us03/_0163_ ;
wire \us03/_0164_ ;
wire \us03/_0165_ ;
wire \us03/_0166_ ;
wire \us03/_0167_ ;
wire \us03/_0168_ ;
wire \us03/_0169_ ;
wire \us03/_0170_ ;
wire \us03/_0171_ ;
wire \us03/_0172_ ;
wire \us03/_0174_ ;
wire \us03/_0175_ ;
wire \us03/_0176_ ;
wire \us03/_0177_ ;
wire \us03/_0178_ ;
wire \us03/_0179_ ;
wire \us03/_0180_ ;
wire \us03/_0181_ ;
wire \us03/_0182_ ;
wire \us03/_0183_ ;
wire \us03/_0184_ ;
wire \us03/_0185_ ;
wire \us03/_0186_ ;
wire \us03/_0187_ ;
wire \us03/_0188_ ;
wire \us03/_0189_ ;
wire \us03/_0190_ ;
wire \us03/_0191_ ;
wire \us03/_0192_ ;
wire \us03/_0193_ ;
wire \us03/_0194_ ;
wire \us03/_0195_ ;
wire \us03/_0196_ ;
wire \us03/_0197_ ;
wire \us03/_0198_ ;
wire \us03/_0199_ ;
wire \us03/_0200_ ;
wire \us03/_0201_ ;
wire \us03/_0202_ ;
wire \us03/_0203_ ;
wire \us03/_0204_ ;
wire \us03/_0205_ ;
wire \us03/_0206_ ;
wire \us03/_0207_ ;
wire \us03/_0208_ ;
wire \us03/_0209_ ;
wire \us03/_0210_ ;
wire \us03/_0211_ ;
wire \us03/_0212_ ;
wire \us03/_0213_ ;
wire \us03/_0214_ ;
wire \us03/_0215_ ;
wire \us03/_0216_ ;
wire \us03/_0217_ ;
wire \us03/_0219_ ;
wire \us03/_0220_ ;
wire \us03/_0221_ ;
wire \us03/_0222_ ;
wire \us03/_0223_ ;
wire \us03/_0224_ ;
wire \us03/_0225_ ;
wire \us03/_0226_ ;
wire \us03/_0227_ ;
wire \us03/_0228_ ;
wire \us03/_0229_ ;
wire \us03/_0230_ ;
wire \us03/_0231_ ;
wire \us03/_0232_ ;
wire \us03/_0233_ ;
wire \us03/_0234_ ;
wire \us03/_0235_ ;
wire \us03/_0236_ ;
wire \us03/_0237_ ;
wire \us03/_0238_ ;
wire \us03/_0239_ ;
wire \us03/_0240_ ;
wire \us03/_0241_ ;
wire \us03/_0242_ ;
wire \us03/_0243_ ;
wire \us03/_0244_ ;
wire \us03/_0245_ ;
wire \us03/_0246_ ;
wire \us03/_0247_ ;
wire \us03/_0248_ ;
wire \us03/_0249_ ;
wire \us03/_0250_ ;
wire \us03/_0251_ ;
wire \us03/_0252_ ;
wire \us03/_0253_ ;
wire \us03/_0254_ ;
wire \us03/_0255_ ;
wire \us03/_0256_ ;
wire \us03/_0257_ ;
wire \us03/_0258_ ;
wire \us03/_0259_ ;
wire \us03/_0260_ ;
wire \us03/_0261_ ;
wire \us03/_0263_ ;
wire \us03/_0264_ ;
wire \us03/_0265_ ;
wire \us03/_0266_ ;
wire \us03/_0267_ ;
wire \us03/_0268_ ;
wire \us03/_0269_ ;
wire \us03/_0270_ ;
wire \us03/_0271_ ;
wire \us03/_0272_ ;
wire \us03/_0273_ ;
wire \us03/_0274_ ;
wire \us03/_0275_ ;
wire \us03/_0276_ ;
wire \us03/_0277_ ;
wire \us03/_0278_ ;
wire \us03/_0279_ ;
wire \us03/_0280_ ;
wire \us03/_0281_ ;
wire \us03/_0283_ ;
wire \us03/_0284_ ;
wire \us03/_0285_ ;
wire \us03/_0286_ ;
wire \us03/_0287_ ;
wire \us03/_0288_ ;
wire \us03/_0289_ ;
wire \us03/_0290_ ;
wire \us03/_0291_ ;
wire \us03/_0293_ ;
wire \us03/_0294_ ;
wire \us03/_0295_ ;
wire \us03/_0296_ ;
wire \us03/_0297_ ;
wire \us03/_0298_ ;
wire \us03/_0299_ ;
wire \us03/_0300_ ;
wire \us03/_0301_ ;
wire \us03/_0302_ ;
wire \us03/_0303_ ;
wire \us03/_0304_ ;
wire \us03/_0305_ ;
wire \us03/_0306_ ;
wire \us03/_0307_ ;
wire \us03/_0308_ ;
wire \us03/_0309_ ;
wire \us03/_0310_ ;
wire \us03/_0311_ ;
wire \us03/_0312_ ;
wire \us03/_0313_ ;
wire \us03/_0314_ ;
wire \us03/_0315_ ;
wire \us03/_0316_ ;
wire \us03/_0317_ ;
wire \us03/_0318_ ;
wire \us03/_0319_ ;
wire \us03/_0320_ ;
wire \us03/_0321_ ;
wire \us03/_0322_ ;
wire \us03/_0323_ ;
wire \us03/_0324_ ;
wire \us03/_0325_ ;
wire \us03/_0326_ ;
wire \us03/_0327_ ;
wire \us03/_0328_ ;
wire \us03/_0329_ ;
wire \us03/_0330_ ;
wire \us03/_0331_ ;
wire \us03/_0332_ ;
wire \us03/_0333_ ;
wire \us03/_0334_ ;
wire \us03/_0335_ ;
wire \us03/_0337_ ;
wire \us03/_0338_ ;
wire \us03/_0339_ ;
wire \us03/_0340_ ;
wire \us03/_0341_ ;
wire \us03/_0342_ ;
wire \us03/_0343_ ;
wire \us03/_0344_ ;
wire \us03/_0345_ ;
wire \us03/_0347_ ;
wire \us03/_0348_ ;
wire \us03/_0349_ ;
wire \us03/_0350_ ;
wire \us03/_0351_ ;
wire \us03/_0352_ ;
wire \us03/_0353_ ;
wire \us03/_0354_ ;
wire \us03/_0355_ ;
wire \us03/_0356_ ;
wire \us03/_0357_ ;
wire \us03/_0358_ ;
wire \us03/_0359_ ;
wire \us03/_0360_ ;
wire \us03/_0361_ ;
wire \us03/_0362_ ;
wire \us03/_0363_ ;
wire \us03/_0364_ ;
wire \us03/_0365_ ;
wire \us03/_0366_ ;
wire \us03/_0367_ ;
wire \us03/_0368_ ;
wire \us03/_0370_ ;
wire \us03/_0371_ ;
wire \us03/_0372_ ;
wire \us03/_0373_ ;
wire \us03/_0374_ ;
wire \us03/_0375_ ;
wire \us03/_0376_ ;
wire \us03/_0377_ ;
wire \us03/_0378_ ;
wire \us03/_0379_ ;
wire \us03/_0380_ ;
wire \us03/_0381_ ;
wire \us03/_0382_ ;
wire \us03/_0383_ ;
wire \us03/_0384_ ;
wire \us03/_0385_ ;
wire \us03/_0386_ ;
wire \us03/_0387_ ;
wire \us03/_0388_ ;
wire \us03/_0389_ ;
wire \us03/_0390_ ;
wire \us03/_0391_ ;
wire \us03/_0392_ ;
wire \us03/_0393_ ;
wire \us03/_0394_ ;
wire \us03/_0395_ ;
wire \us03/_0396_ ;
wire \us03/_0397_ ;
wire \us03/_0398_ ;
wire \us03/_0399_ ;
wire \us03/_0400_ ;
wire \us03/_0401_ ;
wire \us03/_0402_ ;
wire \us03/_0403_ ;
wire \us03/_0404_ ;
wire \us03/_0405_ ;
wire \us03/_0406_ ;
wire \us03/_0407_ ;
wire \us03/_0408_ ;
wire \us03/_0409_ ;
wire \us03/_0410_ ;
wire \us03/_0411_ ;
wire \us03/_0412_ ;
wire \us03/_0413_ ;
wire \us03/_0414_ ;
wire \us03/_0415_ ;
wire \us03/_0416_ ;
wire \us03/_0417_ ;
wire \us03/_0418_ ;
wire \us03/_0419_ ;
wire \us03/_0420_ ;
wire \us03/_0421_ ;
wire \us03/_0422_ ;
wire \us03/_0424_ ;
wire \us03/_0425_ ;
wire \us03/_0426_ ;
wire \us03/_0427_ ;
wire \us03/_0428_ ;
wire \us03/_0429_ ;
wire \us03/_0430_ ;
wire \us03/_0431_ ;
wire \us03/_0432_ ;
wire \us03/_0433_ ;
wire \us03/_0434_ ;
wire \us03/_0435_ ;
wire \us03/_0436_ ;
wire \us03/_0437_ ;
wire \us03/_0438_ ;
wire \us03/_0439_ ;
wire \us03/_0440_ ;
wire \us03/_0441_ ;
wire \us03/_0442_ ;
wire \us03/_0443_ ;
wire \us03/_0444_ ;
wire \us03/_0446_ ;
wire \us03/_0447_ ;
wire \us03/_0448_ ;
wire \us03/_0449_ ;
wire \us03/_0450_ ;
wire \us03/_0451_ ;
wire \us03/_0452_ ;
wire \us03/_0453_ ;
wire \us03/_0454_ ;
wire \us03/_0455_ ;
wire \us03/_0457_ ;
wire \us03/_0458_ ;
wire \us03/_0459_ ;
wire \us03/_0460_ ;
wire \us03/_0461_ ;
wire \us03/_0462_ ;
wire \us03/_0463_ ;
wire \us03/_0464_ ;
wire \us03/_0465_ ;
wire \us03/_0466_ ;
wire \us03/_0467_ ;
wire \us03/_0468_ ;
wire \us03/_0469_ ;
wire \us03/_0470_ ;
wire \us03/_0471_ ;
wire \us03/_0472_ ;
wire \us03/_0473_ ;
wire \us03/_0474_ ;
wire \us03/_0475_ ;
wire \us03/_0476_ ;
wire \us03/_0477_ ;
wire \us03/_0478_ ;
wire \us03/_0479_ ;
wire \us03/_0480_ ;
wire \us03/_0481_ ;
wire \us03/_0482_ ;
wire \us03/_0483_ ;
wire \us03/_0484_ ;
wire \us03/_0485_ ;
wire \us03/_0486_ ;
wire \us03/_0487_ ;
wire \us03/_0488_ ;
wire \us03/_0489_ ;
wire \us03/_0490_ ;
wire \us03/_0491_ ;
wire \us03/_0492_ ;
wire \us03/_0493_ ;
wire \us03/_0494_ ;
wire \us03/_0495_ ;
wire \us03/_0496_ ;
wire \us03/_0497_ ;
wire \us03/_0498_ ;
wire \us03/_0499_ ;
wire \us03/_0500_ ;
wire \us03/_0501_ ;
wire \us03/_0502_ ;
wire \us03/_0503_ ;
wire \us03/_0504_ ;
wire \us03/_0505_ ;
wire \us03/_0506_ ;
wire \us03/_0507_ ;
wire \us03/_0508_ ;
wire \us03/_0509_ ;
wire \us03/_0510_ ;
wire \us03/_0511_ ;
wire \us03/_0512_ ;
wire \us03/_0513_ ;
wire \us03/_0514_ ;
wire \us03/_0515_ ;
wire \us03/_0516_ ;
wire \us03/_0517_ ;
wire \us03/_0518_ ;
wire \us03/_0519_ ;
wire \us03/_0520_ ;
wire \us03/_0521_ ;
wire \us03/_0522_ ;
wire \us03/_0523_ ;
wire \us03/_0524_ ;
wire \us03/_0525_ ;
wire \us03/_0526_ ;
wire \us03/_0527_ ;
wire \us03/_0528_ ;
wire \us03/_0529_ ;
wire \us03/_0530_ ;
wire \us03/_0531_ ;
wire \us03/_0532_ ;
wire \us03/_0533_ ;
wire \us03/_0534_ ;
wire \us03/_0535_ ;
wire \us03/_0536_ ;
wire \us03/_0537_ ;
wire \us03/_0538_ ;
wire \us03/_0539_ ;
wire \us03/_0540_ ;
wire \us03/_0541_ ;
wire \us03/_0542_ ;
wire \us03/_0543_ ;
wire \us03/_0544_ ;
wire \us03/_0545_ ;
wire \us03/_0546_ ;
wire \us03/_0547_ ;
wire \us03/_0548_ ;
wire \us03/_0549_ ;
wire \us03/_0550_ ;
wire \us03/_0551_ ;
wire \us03/_0552_ ;
wire \us03/_0553_ ;
wire \us03/_0554_ ;
wire \us03/_0555_ ;
wire \us03/_0556_ ;
wire \us03/_0557_ ;
wire \us03/_0558_ ;
wire \us03/_0559_ ;
wire \us03/_0560_ ;
wire \us03/_0561_ ;
wire \us03/_0562_ ;
wire \us03/_0563_ ;
wire \us03/_0565_ ;
wire \us03/_0566_ ;
wire \us03/_0567_ ;
wire \us03/_0568_ ;
wire \us03/_0569_ ;
wire \us03/_0570_ ;
wire \us03/_0571_ ;
wire \us03/_0572_ ;
wire \us03/_0573_ ;
wire \us03/_0574_ ;
wire \us03/_0575_ ;
wire \us03/_0576_ ;
wire \us03/_0577_ ;
wire \us03/_0578_ ;
wire \us03/_0579_ ;
wire \us03/_0580_ ;
wire \us03/_0581_ ;
wire \us03/_0582_ ;
wire \us03/_0583_ ;
wire \us03/_0584_ ;
wire \us03/_0585_ ;
wire \us03/_0586_ ;
wire \us03/_0587_ ;
wire \us03/_0588_ ;
wire \us03/_0589_ ;
wire \us03/_0590_ ;
wire \us03/_0591_ ;
wire \us03/_0592_ ;
wire \us03/_0593_ ;
wire \us03/_0594_ ;
wire \us03/_0595_ ;
wire \us03/_0596_ ;
wire \us03/_0598_ ;
wire \us03/_0599_ ;
wire \us03/_0600_ ;
wire \us03/_0601_ ;
wire \us03/_0602_ ;
wire \us03/_0603_ ;
wire \us03/_0604_ ;
wire \us03/_0605_ ;
wire \us03/_0606_ ;
wire \us03/_0607_ ;
wire \us03/_0608_ ;
wire \us03/_0609_ ;
wire \us03/_0610_ ;
wire \us03/_0611_ ;
wire \us03/_0612_ ;
wire \us03/_0613_ ;
wire \us03/_0614_ ;
wire \us03/_0615_ ;
wire \us03/_0616_ ;
wire \us03/_0617_ ;
wire \us03/_0618_ ;
wire \us03/_0619_ ;
wire \us03/_0620_ ;
wire \us03/_0621_ ;
wire \us03/_0622_ ;
wire \us03/_0623_ ;
wire \us03/_0624_ ;
wire \us03/_0625_ ;
wire \us03/_0626_ ;
wire \us03/_0627_ ;
wire \us03/_0628_ ;
wire \us03/_0629_ ;
wire \us03/_0630_ ;
wire \us03/_0631_ ;
wire \us03/_0632_ ;
wire \us03/_0633_ ;
wire \us03/_0634_ ;
wire \us03/_0635_ ;
wire \us03/_0636_ ;
wire \us03/_0637_ ;
wire \us03/_0638_ ;
wire \us03/_0639_ ;
wire \us03/_0640_ ;
wire \us03/_0641_ ;
wire \us03/_0642_ ;
wire \us03/_0643_ ;
wire \us03/_0644_ ;
wire \us03/_0645_ ;
wire \us03/_0646_ ;
wire \us03/_0647_ ;
wire \us03/_0648_ ;
wire \us03/_0649_ ;
wire \us03/_0650_ ;
wire \us03/_0652_ ;
wire \us03/_0653_ ;
wire \us03/_0654_ ;
wire \us03/_0655_ ;
wire \us03/_0656_ ;
wire \us03/_0657_ ;
wire \us03/_0658_ ;
wire \us03/_0659_ ;
wire \us03/_0660_ ;
wire \us03/_0661_ ;
wire \us03/_0662_ ;
wire \us03/_0663_ ;
wire \us03/_0664_ ;
wire \us03/_0665_ ;
wire \us03/_0666_ ;
wire \us03/_0667_ ;
wire \us03/_0668_ ;
wire \us03/_0669_ ;
wire \us03/_0670_ ;
wire \us03/_0671_ ;
wire \us03/_0672_ ;
wire \us03/_0673_ ;
wire \us03/_0674_ ;
wire \us03/_0675_ ;
wire \us03/_0676_ ;
wire \us03/_0677_ ;
wire \us03/_0678_ ;
wire \us03/_0679_ ;
wire \us03/_0680_ ;
wire \us03/_0681_ ;
wire \us03/_0682_ ;
wire \us03/_0683_ ;
wire \us03/_0684_ ;
wire \us03/_0685_ ;
wire \us03/_0686_ ;
wire \us03/_0687_ ;
wire \us03/_0688_ ;
wire \us03/_0689_ ;
wire \us03/_0690_ ;
wire \us03/_0691_ ;
wire \us03/_0692_ ;
wire \us03/_0693_ ;
wire \us03/_0694_ ;
wire \us03/_0695_ ;
wire \us03/_0696_ ;
wire \us03/_0697_ ;
wire \us03/_0698_ ;
wire \us03/_0699_ ;
wire \us03/_0700_ ;
wire \us03/_0701_ ;
wire \us03/_0702_ ;
wire \us03/_0703_ ;
wire \us03/_0704_ ;
wire \us03/_0705_ ;
wire \us03/_0706_ ;
wire \us03/_0707_ ;
wire \us03/_0708_ ;
wire \us03/_0709_ ;
wire \us03/_0710_ ;
wire \us03/_0711_ ;
wire \us03/_0712_ ;
wire \us03/_0713_ ;
wire \us03/_0714_ ;
wire \us03/_0715_ ;
wire \us03/_0717_ ;
wire \us03/_0718_ ;
wire \us03/_0719_ ;
wire \us03/_0720_ ;
wire \us03/_0721_ ;
wire \us03/_0722_ ;
wire \us03/_0723_ ;
wire \us03/_0724_ ;
wire \us03/_0725_ ;
wire \us03/_0726_ ;
wire \us03/_0727_ ;
wire \us03/_0728_ ;
wire \us03/_0729_ ;
wire \us03/_0730_ ;
wire \us03/_0731_ ;
wire \us03/_0732_ ;
wire \us03/_0733_ ;
wire \us03/_0734_ ;
wire \us03/_0735_ ;
wire \us03/_0736_ ;
wire \us03/_0738_ ;
wire \us03/_0739_ ;
wire \us03/_0740_ ;
wire \us03/_0741_ ;
wire \us03/_0742_ ;
wire \us03/_0744_ ;
wire \us03/_0745_ ;
wire \us03/_0746_ ;
wire \us03/_0747_ ;
wire \us03/_0748_ ;
wire \us03/_0749_ ;
wire \us03/_0750_ ;
wire \us03/_0752_ ;
wire \us10/_0008_ ;
wire \us10/_0009_ ;
wire \us10/_0010_ ;
wire \us10/_0011_ ;
wire \us10/_0012_ ;
wire \us10/_0013_ ;
wire \us10/_0014_ ;
wire \us10/_0015_ ;
wire \us10/_0016_ ;
wire \us10/_0017_ ;
wire \us10/_0018_ ;
wire \us10/_0019_ ;
wire \us10/_0020_ ;
wire \us10/_0022_ ;
wire \us10/_0023_ ;
wire \us10/_0024_ ;
wire \us10/_0025_ ;
wire \us10/_0026_ ;
wire \us10/_0027_ ;
wire \us10/_0029_ ;
wire \us10/_0030_ ;
wire \us10/_0032_ ;
wire \us10/_0033_ ;
wire \us10/_0034_ ;
wire \us10/_0035_ ;
wire \us10/_0036_ ;
wire \us10/_0037_ ;
wire \us10/_0038_ ;
wire \us10/_0039_ ;
wire \us10/_0040_ ;
wire \us10/_0041_ ;
wire \us10/_0042_ ;
wire \us10/_0043_ ;
wire \us10/_0045_ ;
wire \us10/_0046_ ;
wire \us10/_0047_ ;
wire \us10/_0048_ ;
wire \us10/_0049_ ;
wire \us10/_0050_ ;
wire \us10/_0051_ ;
wire \us10/_0052_ ;
wire \us10/_0053_ ;
wire \us10/_0054_ ;
wire \us10/_0055_ ;
wire \us10/_0056_ ;
wire \us10/_0057_ ;
wire \us10/_0058_ ;
wire \us10/_0060_ ;
wire \us10/_0061_ ;
wire \us10/_0062_ ;
wire \us10/_0064_ ;
wire \us10/_0065_ ;
wire \us10/_0066_ ;
wire \us10/_0067_ ;
wire \us10/_0069_ ;
wire \us10/_0070_ ;
wire \us10/_0072_ ;
wire \us10/_0073_ ;
wire \us10/_0074_ ;
wire \us10/_0075_ ;
wire \us10/_0076_ ;
wire \us10/_0077_ ;
wire \us10/_0078_ ;
wire \us10/_0079_ ;
wire \us10/_0081_ ;
wire \us10/_0082_ ;
wire \us10/_0083_ ;
wire \us10/_0084_ ;
wire \us10/_0085_ ;
wire \us10/_0086_ ;
wire \us10/_0087_ ;
wire \us10/_0088_ ;
wire \us10/_0089_ ;
wire \us10/_0090_ ;
wire \us10/_0091_ ;
wire \us10/_0092_ ;
wire \us10/_0093_ ;
wire \us10/_0094_ ;
wire \us10/_0095_ ;
wire \us10/_0096_ ;
wire \us10/_0097_ ;
wire \us10/_0098_ ;
wire \us10/_0099_ ;
wire \us10/_0100_ ;
wire \us10/_0101_ ;
wire \us10/_0102_ ;
wire \us10/_0103_ ;
wire \us10/_0104_ ;
wire \us10/_0105_ ;
wire \us10/_0106_ ;
wire \us10/_0108_ ;
wire \us10/_0109_ ;
wire \us10/_0110_ ;
wire \us10/_0111_ ;
wire \us10/_0113_ ;
wire \us10/_0114_ ;
wire \us10/_0115_ ;
wire \us10/_0116_ ;
wire \us10/_0117_ ;
wire \us10/_0118_ ;
wire \us10/_0119_ ;
wire \us10/_0120_ ;
wire \us10/_0121_ ;
wire \us10/_0122_ ;
wire \us10/_0123_ ;
wire \us10/_0124_ ;
wire \us10/_0126_ ;
wire \us10/_0127_ ;
wire \us10/_0128_ ;
wire \us10/_0129_ ;
wire \us10/_0130_ ;
wire \us10/_0132_ ;
wire \us10/_0133_ ;
wire \us10/_0134_ ;
wire \us10/_0135_ ;
wire \us10/_0136_ ;
wire \us10/_0137_ ;
wire \us10/_0139_ ;
wire \us10/_0140_ ;
wire \us10/_0141_ ;
wire \us10/_0142_ ;
wire \us10/_0144_ ;
wire \us10/_0145_ ;
wire \us10/_0146_ ;
wire \us10/_0147_ ;
wire \us10/_0148_ ;
wire \us10/_0149_ ;
wire \us10/_0150_ ;
wire \us10/_0151_ ;
wire \us10/_0153_ ;
wire \us10/_0154_ ;
wire \us10/_0155_ ;
wire \us10/_0156_ ;
wire \us10/_0157_ ;
wire \us10/_0158_ ;
wire \us10/_0159_ ;
wire \us10/_0161_ ;
wire \us10/_0162_ ;
wire \us10/_0163_ ;
wire \us10/_0164_ ;
wire \us10/_0165_ ;
wire \us10/_0166_ ;
wire \us10/_0167_ ;
wire \us10/_0168_ ;
wire \us10/_0169_ ;
wire \us10/_0170_ ;
wire \us10/_0171_ ;
wire \us10/_0172_ ;
wire \us10/_0174_ ;
wire \us10/_0175_ ;
wire \us10/_0176_ ;
wire \us10/_0177_ ;
wire \us10/_0178_ ;
wire \us10/_0179_ ;
wire \us10/_0180_ ;
wire \us10/_0181_ ;
wire \us10/_0182_ ;
wire \us10/_0183_ ;
wire \us10/_0184_ ;
wire \us10/_0185_ ;
wire \us10/_0186_ ;
wire \us10/_0187_ ;
wire \us10/_0188_ ;
wire \us10/_0189_ ;
wire \us10/_0190_ ;
wire \us10/_0191_ ;
wire \us10/_0192_ ;
wire \us10/_0193_ ;
wire \us10/_0194_ ;
wire \us10/_0195_ ;
wire \us10/_0196_ ;
wire \us10/_0197_ ;
wire \us10/_0198_ ;
wire \us10/_0199_ ;
wire \us10/_0200_ ;
wire \us10/_0201_ ;
wire \us10/_0202_ ;
wire \us10/_0203_ ;
wire \us10/_0204_ ;
wire \us10/_0205_ ;
wire \us10/_0206_ ;
wire \us10/_0207_ ;
wire \us10/_0208_ ;
wire \us10/_0209_ ;
wire \us10/_0210_ ;
wire \us10/_0211_ ;
wire \us10/_0212_ ;
wire \us10/_0213_ ;
wire \us10/_0214_ ;
wire \us10/_0215_ ;
wire \us10/_0216_ ;
wire \us10/_0217_ ;
wire \us10/_0218_ ;
wire \us10/_0219_ ;
wire \us10/_0220_ ;
wire \us10/_0221_ ;
wire \us10/_0222_ ;
wire \us10/_0223_ ;
wire \us10/_0224_ ;
wire \us10/_0225_ ;
wire \us10/_0226_ ;
wire \us10/_0227_ ;
wire \us10/_0228_ ;
wire \us10/_0229_ ;
wire \us10/_0230_ ;
wire \us10/_0231_ ;
wire \us10/_0232_ ;
wire \us10/_0233_ ;
wire \us10/_0234_ ;
wire \us10/_0235_ ;
wire \us10/_0236_ ;
wire \us10/_0237_ ;
wire \us10/_0238_ ;
wire \us10/_0239_ ;
wire \us10/_0240_ ;
wire \us10/_0241_ ;
wire \us10/_0242_ ;
wire \us10/_0243_ ;
wire \us10/_0244_ ;
wire \us10/_0245_ ;
wire \us10/_0246_ ;
wire \us10/_0248_ ;
wire \us10/_0249_ ;
wire \us10/_0250_ ;
wire \us10/_0251_ ;
wire \us10/_0252_ ;
wire \us10/_0253_ ;
wire \us10/_0254_ ;
wire \us10/_0255_ ;
wire \us10/_0256_ ;
wire \us10/_0257_ ;
wire \us10/_0258_ ;
wire \us10/_0259_ ;
wire \us10/_0260_ ;
wire \us10/_0261_ ;
wire \us10/_0263_ ;
wire \us10/_0264_ ;
wire \us10/_0265_ ;
wire \us10/_0266_ ;
wire \us10/_0267_ ;
wire \us10/_0268_ ;
wire \us10/_0269_ ;
wire \us10/_0270_ ;
wire \us10/_0271_ ;
wire \us10/_0272_ ;
wire \us10/_0273_ ;
wire \us10/_0274_ ;
wire \us10/_0275_ ;
wire \us10/_0276_ ;
wire \us10/_0277_ ;
wire \us10/_0278_ ;
wire \us10/_0279_ ;
wire \us10/_0281_ ;
wire \us10/_0282_ ;
wire \us10/_0283_ ;
wire \us10/_0284_ ;
wire \us10/_0285_ ;
wire \us10/_0286_ ;
wire \us10/_0287_ ;
wire \us10/_0288_ ;
wire \us10/_0289_ ;
wire \us10/_0290_ ;
wire \us10/_0291_ ;
wire \us10/_0293_ ;
wire \us10/_0294_ ;
wire \us10/_0295_ ;
wire \us10/_0296_ ;
wire \us10/_0297_ ;
wire \us10/_0298_ ;
wire \us10/_0299_ ;
wire \us10/_0300_ ;
wire \us10/_0301_ ;
wire \us10/_0302_ ;
wire \us10/_0303_ ;
wire \us10/_0304_ ;
wire \us10/_0305_ ;
wire \us10/_0306_ ;
wire \us10/_0307_ ;
wire \us10/_0308_ ;
wire \us10/_0309_ ;
wire \us10/_0310_ ;
wire \us10/_0311_ ;
wire \us10/_0312_ ;
wire \us10/_0313_ ;
wire \us10/_0314_ ;
wire \us10/_0315_ ;
wire \us10/_0316_ ;
wire \us10/_0317_ ;
wire \us10/_0318_ ;
wire \us10/_0319_ ;
wire \us10/_0320_ ;
wire \us10/_0321_ ;
wire \us10/_0322_ ;
wire \us10/_0323_ ;
wire \us10/_0324_ ;
wire \us10/_0325_ ;
wire \us10/_0326_ ;
wire \us10/_0327_ ;
wire \us10/_0328_ ;
wire \us10/_0329_ ;
wire \us10/_0330_ ;
wire \us10/_0331_ ;
wire \us10/_0332_ ;
wire \us10/_0333_ ;
wire \us10/_0334_ ;
wire \us10/_0335_ ;
wire \us10/_0337_ ;
wire \us10/_0338_ ;
wire \us10/_0339_ ;
wire \us10/_0340_ ;
wire \us10/_0341_ ;
wire \us10/_0342_ ;
wire \us10/_0343_ ;
wire \us10/_0344_ ;
wire \us10/_0345_ ;
wire \us10/_0347_ ;
wire \us10/_0348_ ;
wire \us10/_0349_ ;
wire \us10/_0350_ ;
wire \us10/_0351_ ;
wire \us10/_0352_ ;
wire \us10/_0353_ ;
wire \us10/_0354_ ;
wire \us10/_0355_ ;
wire \us10/_0356_ ;
wire \us10/_0357_ ;
wire \us10/_0358_ ;
wire \us10/_0359_ ;
wire \us10/_0360_ ;
wire \us10/_0361_ ;
wire \us10/_0362_ ;
wire \us10/_0363_ ;
wire \us10/_0365_ ;
wire \us10/_0366_ ;
wire \us10/_0367_ ;
wire \us10/_0368_ ;
wire \us10/_0370_ ;
wire \us10/_0371_ ;
wire \us10/_0372_ ;
wire \us10/_0373_ ;
wire \us10/_0374_ ;
wire \us10/_0375_ ;
wire \us10/_0376_ ;
wire \us10/_0377_ ;
wire \us10/_0378_ ;
wire \us10/_0379_ ;
wire \us10/_0380_ ;
wire \us10/_0381_ ;
wire \us10/_0382_ ;
wire \us10/_0383_ ;
wire \us10/_0384_ ;
wire \us10/_0385_ ;
wire \us10/_0386_ ;
wire \us10/_0387_ ;
wire \us10/_0388_ ;
wire \us10/_0389_ ;
wire \us10/_0390_ ;
wire \us10/_0391_ ;
wire \us10/_0392_ ;
wire \us10/_0393_ ;
wire \us10/_0394_ ;
wire \us10/_0395_ ;
wire \us10/_0396_ ;
wire \us10/_0397_ ;
wire \us10/_0398_ ;
wire \us10/_0399_ ;
wire \us10/_0400_ ;
wire \us10/_0401_ ;
wire \us10/_0402_ ;
wire \us10/_0403_ ;
wire \us10/_0404_ ;
wire \us10/_0405_ ;
wire \us10/_0406_ ;
wire \us10/_0407_ ;
wire \us10/_0408_ ;
wire \us10/_0409_ ;
wire \us10/_0410_ ;
wire \us10/_0411_ ;
wire \us10/_0412_ ;
wire \us10/_0413_ ;
wire \us10/_0414_ ;
wire \us10/_0415_ ;
wire \us10/_0416_ ;
wire \us10/_0417_ ;
wire \us10/_0418_ ;
wire \us10/_0419_ ;
wire \us10/_0420_ ;
wire \us10/_0421_ ;
wire \us10/_0422_ ;
wire \us10/_0423_ ;
wire \us10/_0424_ ;
wire \us10/_0425_ ;
wire \us10/_0426_ ;
wire \us10/_0427_ ;
wire \us10/_0428_ ;
wire \us10/_0429_ ;
wire \us10/_0430_ ;
wire \us10/_0431_ ;
wire \us10/_0432_ ;
wire \us10/_0433_ ;
wire \us10/_0434_ ;
wire \us10/_0435_ ;
wire \us10/_0436_ ;
wire \us10/_0437_ ;
wire \us10/_0438_ ;
wire \us10/_0439_ ;
wire \us10/_0440_ ;
wire \us10/_0441_ ;
wire \us10/_0442_ ;
wire \us10/_0443_ ;
wire \us10/_0444_ ;
wire \us10/_0445_ ;
wire \us10/_0446_ ;
wire \us10/_0447_ ;
wire \us10/_0448_ ;
wire \us10/_0449_ ;
wire \us10/_0450_ ;
wire \us10/_0451_ ;
wire \us10/_0452_ ;
wire \us10/_0453_ ;
wire \us10/_0454_ ;
wire \us10/_0455_ ;
wire \us10/_0457_ ;
wire \us10/_0458_ ;
wire \us10/_0459_ ;
wire \us10/_0460_ ;
wire \us10/_0461_ ;
wire \us10/_0462_ ;
wire \us10/_0463_ ;
wire \us10/_0464_ ;
wire \us10/_0465_ ;
wire \us10/_0466_ ;
wire \us10/_0467_ ;
wire \us10/_0468_ ;
wire \us10/_0469_ ;
wire \us10/_0470_ ;
wire \us10/_0471_ ;
wire \us10/_0472_ ;
wire \us10/_0473_ ;
wire \us10/_0474_ ;
wire \us10/_0475_ ;
wire \us10/_0476_ ;
wire \us10/_0477_ ;
wire \us10/_0478_ ;
wire \us10/_0479_ ;
wire \us10/_0480_ ;
wire \us10/_0481_ ;
wire \us10/_0482_ ;
wire \us10/_0483_ ;
wire \us10/_0484_ ;
wire \us10/_0485_ ;
wire \us10/_0486_ ;
wire \us10/_0487_ ;
wire \us10/_0488_ ;
wire \us10/_0489_ ;
wire \us10/_0490_ ;
wire \us10/_0491_ ;
wire \us10/_0492_ ;
wire \us10/_0493_ ;
wire \us10/_0494_ ;
wire \us10/_0495_ ;
wire \us10/_0496_ ;
wire \us10/_0497_ ;
wire \us10/_0498_ ;
wire \us10/_0500_ ;
wire \us10/_0501_ ;
wire \us10/_0502_ ;
wire \us10/_0503_ ;
wire \us10/_0504_ ;
wire \us10/_0505_ ;
wire \us10/_0506_ ;
wire \us10/_0507_ ;
wire \us10/_0508_ ;
wire \us10/_0509_ ;
wire \us10/_0510_ ;
wire \us10/_0511_ ;
wire \us10/_0512_ ;
wire \us10/_0513_ ;
wire \us10/_0514_ ;
wire \us10/_0515_ ;
wire \us10/_0516_ ;
wire \us10/_0517_ ;
wire \us10/_0518_ ;
wire \us10/_0519_ ;
wire \us10/_0520_ ;
wire \us10/_0521_ ;
wire \us10/_0522_ ;
wire \us10/_0523_ ;
wire \us10/_0524_ ;
wire \us10/_0525_ ;
wire \us10/_0526_ ;
wire \us10/_0527_ ;
wire \us10/_0528_ ;
wire \us10/_0529_ ;
wire \us10/_0530_ ;
wire \us10/_0531_ ;
wire \us10/_0532_ ;
wire \us10/_0533_ ;
wire \us10/_0534_ ;
wire \us10/_0535_ ;
wire \us10/_0536_ ;
wire \us10/_0537_ ;
wire \us10/_0538_ ;
wire \us10/_0539_ ;
wire \us10/_0540_ ;
wire \us10/_0541_ ;
wire \us10/_0542_ ;
wire \us10/_0543_ ;
wire \us10/_0544_ ;
wire \us10/_0545_ ;
wire \us10/_0546_ ;
wire \us10/_0547_ ;
wire \us10/_0548_ ;
wire \us10/_0549_ ;
wire \us10/_0550_ ;
wire \us10/_0551_ ;
wire \us10/_0552_ ;
wire \us10/_0553_ ;
wire \us10/_0554_ ;
wire \us10/_0555_ ;
wire \us10/_0556_ ;
wire \us10/_0557_ ;
wire \us10/_0558_ ;
wire \us10/_0559_ ;
wire \us10/_0560_ ;
wire \us10/_0561_ ;
wire \us10/_0562_ ;
wire \us10/_0563_ ;
wire \us10/_0565_ ;
wire \us10/_0566_ ;
wire \us10/_0567_ ;
wire \us10/_0568_ ;
wire \us10/_0569_ ;
wire \us10/_0570_ ;
wire \us10/_0571_ ;
wire \us10/_0572_ ;
wire \us10/_0573_ ;
wire \us10/_0574_ ;
wire \us10/_0575_ ;
wire \us10/_0576_ ;
wire \us10/_0577_ ;
wire \us10/_0578_ ;
wire \us10/_0579_ ;
wire \us10/_0580_ ;
wire \us10/_0581_ ;
wire \us10/_0582_ ;
wire \us10/_0583_ ;
wire \us10/_0584_ ;
wire \us10/_0585_ ;
wire \us10/_0586_ ;
wire \us10/_0587_ ;
wire \us10/_0588_ ;
wire \us10/_0589_ ;
wire \us10/_0590_ ;
wire \us10/_0591_ ;
wire \us10/_0592_ ;
wire \us10/_0593_ ;
wire \us10/_0594_ ;
wire \us10/_0595_ ;
wire \us10/_0596_ ;
wire \us10/_0598_ ;
wire \us10/_0599_ ;
wire \us10/_0600_ ;
wire \us10/_0601_ ;
wire \us10/_0602_ ;
wire \us10/_0603_ ;
wire \us10/_0604_ ;
wire \us10/_0605_ ;
wire \us10/_0606_ ;
wire \us10/_0607_ ;
wire \us10/_0608_ ;
wire \us10/_0609_ ;
wire \us10/_0610_ ;
wire \us10/_0611_ ;
wire \us10/_0612_ ;
wire \us10/_0613_ ;
wire \us10/_0614_ ;
wire \us10/_0615_ ;
wire \us10/_0616_ ;
wire \us10/_0617_ ;
wire \us10/_0618_ ;
wire \us10/_0619_ ;
wire \us10/_0620_ ;
wire \us10/_0621_ ;
wire \us10/_0622_ ;
wire \us10/_0623_ ;
wire \us10/_0624_ ;
wire \us10/_0625_ ;
wire \us10/_0626_ ;
wire \us10/_0627_ ;
wire \us10/_0628_ ;
wire \us10/_0629_ ;
wire \us10/_0630_ ;
wire \us10/_0631_ ;
wire \us10/_0632_ ;
wire \us10/_0633_ ;
wire \us10/_0634_ ;
wire \us10/_0635_ ;
wire \us10/_0636_ ;
wire \us10/_0637_ ;
wire \us10/_0638_ ;
wire \us10/_0639_ ;
wire \us10/_0640_ ;
wire \us10/_0641_ ;
wire \us10/_0642_ ;
wire \us10/_0643_ ;
wire \us10/_0644_ ;
wire \us10/_0645_ ;
wire \us10/_0646_ ;
wire \us10/_0647_ ;
wire \us10/_0648_ ;
wire \us10/_0649_ ;
wire \us10/_0650_ ;
wire \us10/_0652_ ;
wire \us10/_0653_ ;
wire \us10/_0654_ ;
wire \us10/_0655_ ;
wire \us10/_0656_ ;
wire \us10/_0657_ ;
wire \us10/_0658_ ;
wire \us10/_0659_ ;
wire \us10/_0660_ ;
wire \us10/_0661_ ;
wire \us10/_0662_ ;
wire \us10/_0663_ ;
wire \us10/_0664_ ;
wire \us10/_0665_ ;
wire \us10/_0666_ ;
wire \us10/_0667_ ;
wire \us10/_0668_ ;
wire \us10/_0669_ ;
wire \us10/_0670_ ;
wire \us10/_0671_ ;
wire \us10/_0672_ ;
wire \us10/_0673_ ;
wire \us10/_0674_ ;
wire \us10/_0675_ ;
wire \us10/_0676_ ;
wire \us10/_0677_ ;
wire \us10/_0678_ ;
wire \us10/_0679_ ;
wire \us10/_0680_ ;
wire \us10/_0681_ ;
wire \us10/_0682_ ;
wire \us10/_0683_ ;
wire \us10/_0684_ ;
wire \us10/_0685_ ;
wire \us10/_0686_ ;
wire \us10/_0687_ ;
wire \us10/_0688_ ;
wire \us10/_0689_ ;
wire \us10/_0690_ ;
wire \us10/_0691_ ;
wire \us10/_0692_ ;
wire \us10/_0693_ ;
wire \us10/_0694_ ;
wire \us10/_0695_ ;
wire \us10/_0696_ ;
wire \us10/_0697_ ;
wire \us10/_0698_ ;
wire \us10/_0699_ ;
wire \us10/_0700_ ;
wire \us10/_0701_ ;
wire \us10/_0702_ ;
wire \us10/_0703_ ;
wire \us10/_0704_ ;
wire \us10/_0705_ ;
wire \us10/_0706_ ;
wire \us10/_0707_ ;
wire \us10/_0708_ ;
wire \us10/_0709_ ;
wire \us10/_0710_ ;
wire \us10/_0711_ ;
wire \us10/_0712_ ;
wire \us10/_0713_ ;
wire \us10/_0714_ ;
wire \us10/_0715_ ;
wire \us10/_0717_ ;
wire \us10/_0718_ ;
wire \us10/_0719_ ;
wire \us10/_0720_ ;
wire \us10/_0721_ ;
wire \us10/_0722_ ;
wire \us10/_0723_ ;
wire \us10/_0724_ ;
wire \us10/_0725_ ;
wire \us10/_0726_ ;
wire \us10/_0727_ ;
wire \us10/_0728_ ;
wire \us10/_0729_ ;
wire \us10/_0730_ ;
wire \us10/_0731_ ;
wire \us10/_0732_ ;
wire \us10/_0733_ ;
wire \us10/_0734_ ;
wire \us10/_0735_ ;
wire \us10/_0736_ ;
wire \us10/_0738_ ;
wire \us10/_0739_ ;
wire \us10/_0740_ ;
wire \us10/_0741_ ;
wire \us10/_0742_ ;
wire \us10/_0744_ ;
wire \us10/_0745_ ;
wire \us10/_0746_ ;
wire \us10/_0748_ ;
wire \us10/_0749_ ;
wire \us10/_0750_ ;
wire \us10/_0752_ ;
wire \us11/_0008_ ;
wire \us11/_0009_ ;
wire \us11/_0010_ ;
wire \us11/_0011_ ;
wire \us11/_0012_ ;
wire \us11/_0013_ ;
wire \us11/_0014_ ;
wire \us11/_0015_ ;
wire \us11/_0016_ ;
wire \us11/_0017_ ;
wire \us11/_0019_ ;
wire \us11/_0020_ ;
wire \us11/_0022_ ;
wire \us11/_0024_ ;
wire \us11/_0025_ ;
wire \us11/_0026_ ;
wire \us11/_0027_ ;
wire \us11/_0030_ ;
wire \us11/_0032_ ;
wire \us11/_0033_ ;
wire \us11/_0034_ ;
wire \us11/_0035_ ;
wire \us11/_0037_ ;
wire \us11/_0038_ ;
wire \us11/_0039_ ;
wire \us11/_0040_ ;
wire \us11/_0041_ ;
wire \us11/_0042_ ;
wire \us11/_0043_ ;
wire \us11/_0045_ ;
wire \us11/_0046_ ;
wire \us11/_0047_ ;
wire \us11/_0049_ ;
wire \us11/_0050_ ;
wire \us11/_0051_ ;
wire \us11/_0052_ ;
wire \us11/_0053_ ;
wire \us11/_0054_ ;
wire \us11/_0057_ ;
wire \us11/_0058_ ;
wire \us11/_0060_ ;
wire \us11/_0061_ ;
wire \us11/_0062_ ;
wire \us11/_0064_ ;
wire \us11/_0065_ ;
wire \us11/_0066_ ;
wire \us11/_0067_ ;
wire \us11/_0069_ ;
wire \us11/_0070_ ;
wire \us11/_0072_ ;
wire \us11/_0073_ ;
wire \us11/_0074_ ;
wire \us11/_0075_ ;
wire \us11/_0076_ ;
wire \us11/_0077_ ;
wire \us11/_0078_ ;
wire \us11/_0079_ ;
wire \us11/_0081_ ;
wire \us11/_0082_ ;
wire \us11/_0084_ ;
wire \us11/_0085_ ;
wire \us11/_0086_ ;
wire \us11/_0087_ ;
wire \us11/_0088_ ;
wire \us11/_0089_ ;
wire \us11/_0090_ ;
wire \us11/_0091_ ;
wire \us11/_0092_ ;
wire \us11/_0093_ ;
wire \us11/_0094_ ;
wire \us11/_0095_ ;
wire \us11/_0096_ ;
wire \us11/_0097_ ;
wire \us11/_0098_ ;
wire \us11/_0100_ ;
wire \us11/_0101_ ;
wire \us11/_0102_ ;
wire \us11/_0103_ ;
wire \us11/_0104_ ;
wire \us11/_0105_ ;
wire \us11/_0106_ ;
wire \us11/_0108_ ;
wire \us11/_0109_ ;
wire \us11/_0110_ ;
wire \us11/_0111_ ;
wire \us11/_0113_ ;
wire \us11/_0114_ ;
wire \us11/_0115_ ;
wire \us11/_0116_ ;
wire \us11/_0117_ ;
wire \us11/_0118_ ;
wire \us11/_0119_ ;
wire \us11/_0120_ ;
wire \us11/_0121_ ;
wire \us11/_0122_ ;
wire \us11/_0123_ ;
wire \us11/_0124_ ;
wire \us11/_0126_ ;
wire \us11/_0127_ ;
wire \us11/_0128_ ;
wire \us11/_0129_ ;
wire \us11/_0130_ ;
wire \us11/_0132_ ;
wire \us11/_0133_ ;
wire \us11/_0134_ ;
wire \us11/_0135_ ;
wire \us11/_0136_ ;
wire \us11/_0137_ ;
wire \us11/_0139_ ;
wire \us11/_0140_ ;
wire \us11/_0141_ ;
wire \us11/_0142_ ;
wire \us11/_0144_ ;
wire \us11/_0145_ ;
wire \us11/_0146_ ;
wire \us11/_0147_ ;
wire \us11/_0148_ ;
wire \us11/_0149_ ;
wire \us11/_0150_ ;
wire \us11/_0151_ ;
wire \us11/_0153_ ;
wire \us11/_0154_ ;
wire \us11/_0155_ ;
wire \us11/_0156_ ;
wire \us11/_0157_ ;
wire \us11/_0158_ ;
wire \us11/_0159_ ;
wire \us11/_0161_ ;
wire \us11/_0162_ ;
wire \us11/_0163_ ;
wire \us11/_0164_ ;
wire \us11/_0165_ ;
wire \us11/_0166_ ;
wire \us11/_0167_ ;
wire \us11/_0168_ ;
wire \us11/_0169_ ;
wire \us11/_0170_ ;
wire \us11/_0171_ ;
wire \us11/_0172_ ;
wire \us11/_0174_ ;
wire \us11/_0175_ ;
wire \us11/_0176_ ;
wire \us11/_0177_ ;
wire \us11/_0178_ ;
wire \us11/_0179_ ;
wire \us11/_0180_ ;
wire \us11/_0181_ ;
wire \us11/_0182_ ;
wire \us11/_0183_ ;
wire \us11/_0184_ ;
wire \us11/_0185_ ;
wire \us11/_0186_ ;
wire \us11/_0187_ ;
wire \us11/_0188_ ;
wire \us11/_0189_ ;
wire \us11/_0190_ ;
wire \us11/_0191_ ;
wire \us11/_0192_ ;
wire \us11/_0193_ ;
wire \us11/_0194_ ;
wire \us11/_0195_ ;
wire \us11/_0196_ ;
wire \us11/_0197_ ;
wire \us11/_0198_ ;
wire \us11/_0199_ ;
wire \us11/_0200_ ;
wire \us11/_0201_ ;
wire \us11/_0202_ ;
wire \us11/_0203_ ;
wire \us11/_0204_ ;
wire \us11/_0205_ ;
wire \us11/_0206_ ;
wire \us11/_0207_ ;
wire \us11/_0208_ ;
wire \us11/_0209_ ;
wire \us11/_0210_ ;
wire \us11/_0211_ ;
wire \us11/_0212_ ;
wire \us11/_0213_ ;
wire \us11/_0214_ ;
wire \us11/_0215_ ;
wire \us11/_0216_ ;
wire \us11/_0217_ ;
wire \us11/_0219_ ;
wire \us11/_0220_ ;
wire \us11/_0221_ ;
wire \us11/_0222_ ;
wire \us11/_0223_ ;
wire \us11/_0224_ ;
wire \us11/_0225_ ;
wire \us11/_0226_ ;
wire \us11/_0227_ ;
wire \us11/_0228_ ;
wire \us11/_0229_ ;
wire \us11/_0230_ ;
wire \us11/_0231_ ;
wire \us11/_0232_ ;
wire \us11/_0233_ ;
wire \us11/_0234_ ;
wire \us11/_0235_ ;
wire \us11/_0236_ ;
wire \us11/_0237_ ;
wire \us11/_0238_ ;
wire \us11/_0239_ ;
wire \us11/_0240_ ;
wire \us11/_0241_ ;
wire \us11/_0242_ ;
wire \us11/_0243_ ;
wire \us11/_0244_ ;
wire \us11/_0245_ ;
wire \us11/_0246_ ;
wire \us11/_0247_ ;
wire \us11/_0248_ ;
wire \us11/_0249_ ;
wire \us11/_0250_ ;
wire \us11/_0251_ ;
wire \us11/_0252_ ;
wire \us11/_0253_ ;
wire \us11/_0254_ ;
wire \us11/_0255_ ;
wire \us11/_0256_ ;
wire \us11/_0257_ ;
wire \us11/_0258_ ;
wire \us11/_0259_ ;
wire \us11/_0260_ ;
wire \us11/_0261_ ;
wire \us11/_0263_ ;
wire \us11/_0264_ ;
wire \us11/_0265_ ;
wire \us11/_0266_ ;
wire \us11/_0267_ ;
wire \us11/_0268_ ;
wire \us11/_0269_ ;
wire \us11/_0270_ ;
wire \us11/_0271_ ;
wire \us11/_0272_ ;
wire \us11/_0273_ ;
wire \us11/_0274_ ;
wire \us11/_0275_ ;
wire \us11/_0276_ ;
wire \us11/_0277_ ;
wire \us11/_0278_ ;
wire \us11/_0279_ ;
wire \us11/_0281_ ;
wire \us11/_0283_ ;
wire \us11/_0284_ ;
wire \us11/_0285_ ;
wire \us11/_0286_ ;
wire \us11/_0287_ ;
wire \us11/_0288_ ;
wire \us11/_0289_ ;
wire \us11/_0290_ ;
wire \us11/_0291_ ;
wire \us11/_0292_ ;
wire \us11/_0293_ ;
wire \us11/_0294_ ;
wire \us11/_0295_ ;
wire \us11/_0296_ ;
wire \us11/_0297_ ;
wire \us11/_0298_ ;
wire \us11/_0299_ ;
wire \us11/_0300_ ;
wire \us11/_0301_ ;
wire \us11/_0302_ ;
wire \us11/_0303_ ;
wire \us11/_0304_ ;
wire \us11/_0305_ ;
wire \us11/_0306_ ;
wire \us11/_0307_ ;
wire \us11/_0308_ ;
wire \us11/_0309_ ;
wire \us11/_0310_ ;
wire \us11/_0311_ ;
wire \us11/_0312_ ;
wire \us11/_0313_ ;
wire \us11/_0314_ ;
wire \us11/_0315_ ;
wire \us11/_0316_ ;
wire \us11/_0317_ ;
wire \us11/_0318_ ;
wire \us11/_0319_ ;
wire \us11/_0320_ ;
wire \us11/_0321_ ;
wire \us11/_0322_ ;
wire \us11/_0323_ ;
wire \us11/_0324_ ;
wire \us11/_0325_ ;
wire \us11/_0326_ ;
wire \us11/_0327_ ;
wire \us11/_0328_ ;
wire \us11/_0329_ ;
wire \us11/_0330_ ;
wire \us11/_0331_ ;
wire \us11/_0332_ ;
wire \us11/_0333_ ;
wire \us11/_0334_ ;
wire \us11/_0335_ ;
wire \us11/_0337_ ;
wire \us11/_0338_ ;
wire \us11/_0339_ ;
wire \us11/_0340_ ;
wire \us11/_0341_ ;
wire \us11/_0342_ ;
wire \us11/_0343_ ;
wire \us11/_0344_ ;
wire \us11/_0345_ ;
wire \us11/_0347_ ;
wire \us11/_0348_ ;
wire \us11/_0349_ ;
wire \us11/_0350_ ;
wire \us11/_0351_ ;
wire \us11/_0352_ ;
wire \us11/_0353_ ;
wire \us11/_0354_ ;
wire \us11/_0355_ ;
wire \us11/_0356_ ;
wire \us11/_0357_ ;
wire \us11/_0358_ ;
wire \us11/_0359_ ;
wire \us11/_0360_ ;
wire \us11/_0361_ ;
wire \us11/_0362_ ;
wire \us11/_0363_ ;
wire \us11/_0364_ ;
wire \us11/_0365_ ;
wire \us11/_0366_ ;
wire \us11/_0367_ ;
wire \us11/_0368_ ;
wire \us11/_0370_ ;
wire \us11/_0371_ ;
wire \us11/_0372_ ;
wire \us11/_0373_ ;
wire \us11/_0374_ ;
wire \us11/_0375_ ;
wire \us11/_0376_ ;
wire \us11/_0377_ ;
wire \us11/_0378_ ;
wire \us11/_0379_ ;
wire \us11/_0380_ ;
wire \us11/_0381_ ;
wire \us11/_0382_ ;
wire \us11/_0383_ ;
wire \us11/_0384_ ;
wire \us11/_0385_ ;
wire \us11/_0386_ ;
wire \us11/_0387_ ;
wire \us11/_0388_ ;
wire \us11/_0389_ ;
wire \us11/_0390_ ;
wire \us11/_0391_ ;
wire \us11/_0392_ ;
wire \us11/_0393_ ;
wire \us11/_0394_ ;
wire \us11/_0395_ ;
wire \us11/_0396_ ;
wire \us11/_0397_ ;
wire \us11/_0398_ ;
wire \us11/_0399_ ;
wire \us11/_0400_ ;
wire \us11/_0401_ ;
wire \us11/_0402_ ;
wire \us11/_0403_ ;
wire \us11/_0404_ ;
wire \us11/_0405_ ;
wire \us11/_0406_ ;
wire \us11/_0407_ ;
wire \us11/_0408_ ;
wire \us11/_0409_ ;
wire \us11/_0410_ ;
wire \us11/_0411_ ;
wire \us11/_0412_ ;
wire \us11/_0413_ ;
wire \us11/_0414_ ;
wire \us11/_0415_ ;
wire \us11/_0416_ ;
wire \us11/_0417_ ;
wire \us11/_0418_ ;
wire \us11/_0419_ ;
wire \us11/_0420_ ;
wire \us11/_0421_ ;
wire \us11/_0422_ ;
wire \us11/_0423_ ;
wire \us11/_0424_ ;
wire \us11/_0425_ ;
wire \us11/_0426_ ;
wire \us11/_0427_ ;
wire \us11/_0428_ ;
wire \us11/_0429_ ;
wire \us11/_0430_ ;
wire \us11/_0431_ ;
wire \us11/_0432_ ;
wire \us11/_0433_ ;
wire \us11/_0434_ ;
wire \us11/_0435_ ;
wire \us11/_0436_ ;
wire \us11/_0437_ ;
wire \us11/_0438_ ;
wire \us11/_0439_ ;
wire \us11/_0440_ ;
wire \us11/_0441_ ;
wire \us11/_0442_ ;
wire \us11/_0443_ ;
wire \us11/_0444_ ;
wire \us11/_0446_ ;
wire \us11/_0447_ ;
wire \us11/_0448_ ;
wire \us11/_0449_ ;
wire \us11/_0450_ ;
wire \us11/_0451_ ;
wire \us11/_0452_ ;
wire \us11/_0453_ ;
wire \us11/_0454_ ;
wire \us11/_0455_ ;
wire \us11/_0457_ ;
wire \us11/_0458_ ;
wire \us11/_0459_ ;
wire \us11/_0460_ ;
wire \us11/_0461_ ;
wire \us11/_0462_ ;
wire \us11/_0463_ ;
wire \us11/_0464_ ;
wire \us11/_0465_ ;
wire \us11/_0466_ ;
wire \us11/_0467_ ;
wire \us11/_0468_ ;
wire \us11/_0469_ ;
wire \us11/_0470_ ;
wire \us11/_0471_ ;
wire \us11/_0472_ ;
wire \us11/_0473_ ;
wire \us11/_0474_ ;
wire \us11/_0475_ ;
wire \us11/_0476_ ;
wire \us11/_0477_ ;
wire \us11/_0478_ ;
wire \us11/_0479_ ;
wire \us11/_0480_ ;
wire \us11/_0481_ ;
wire \us11/_0482_ ;
wire \us11/_0483_ ;
wire \us11/_0484_ ;
wire \us11/_0485_ ;
wire \us11/_0486_ ;
wire \us11/_0487_ ;
wire \us11/_0488_ ;
wire \us11/_0490_ ;
wire \us11/_0491_ ;
wire \us11/_0492_ ;
wire \us11/_0493_ ;
wire \us11/_0494_ ;
wire \us11/_0495_ ;
wire \us11/_0496_ ;
wire \us11/_0497_ ;
wire \us11/_0498_ ;
wire \us11/_0499_ ;
wire \us11/_0500_ ;
wire \us11/_0501_ ;
wire \us11/_0502_ ;
wire \us11/_0503_ ;
wire \us11/_0504_ ;
wire \us11/_0505_ ;
wire \us11/_0506_ ;
wire \us11/_0507_ ;
wire \us11/_0508_ ;
wire \us11/_0509_ ;
wire \us11/_0510_ ;
wire \us11/_0511_ ;
wire \us11/_0512_ ;
wire \us11/_0513_ ;
wire \us11/_0514_ ;
wire \us11/_0515_ ;
wire \us11/_0516_ ;
wire \us11/_0517_ ;
wire \us11/_0518_ ;
wire \us11/_0519_ ;
wire \us11/_0520_ ;
wire \us11/_0521_ ;
wire \us11/_0522_ ;
wire \us11/_0523_ ;
wire \us11/_0524_ ;
wire \us11/_0525_ ;
wire \us11/_0526_ ;
wire \us11/_0527_ ;
wire \us11/_0528_ ;
wire \us11/_0529_ ;
wire \us11/_0530_ ;
wire \us11/_0531_ ;
wire \us11/_0532_ ;
wire \us11/_0533_ ;
wire \us11/_0534_ ;
wire \us11/_0535_ ;
wire \us11/_0536_ ;
wire \us11/_0537_ ;
wire \us11/_0538_ ;
wire \us11/_0539_ ;
wire \us11/_0540_ ;
wire \us11/_0541_ ;
wire \us11/_0542_ ;
wire \us11/_0543_ ;
wire \us11/_0544_ ;
wire \us11/_0545_ ;
wire \us11/_0546_ ;
wire \us11/_0547_ ;
wire \us11/_0548_ ;
wire \us11/_0549_ ;
wire \us11/_0550_ ;
wire \us11/_0551_ ;
wire \us11/_0552_ ;
wire \us11/_0553_ ;
wire \us11/_0554_ ;
wire \us11/_0555_ ;
wire \us11/_0556_ ;
wire \us11/_0557_ ;
wire \us11/_0558_ ;
wire \us11/_0559_ ;
wire \us11/_0560_ ;
wire \us11/_0561_ ;
wire \us11/_0562_ ;
wire \us11/_0563_ ;
wire \us11/_0565_ ;
wire \us11/_0566_ ;
wire \us11/_0567_ ;
wire \us11/_0568_ ;
wire \us11/_0569_ ;
wire \us11/_0570_ ;
wire \us11/_0571_ ;
wire \us11/_0572_ ;
wire \us11/_0573_ ;
wire \us11/_0574_ ;
wire \us11/_0575_ ;
wire \us11/_0576_ ;
wire \us11/_0577_ ;
wire \us11/_0578_ ;
wire \us11/_0579_ ;
wire \us11/_0580_ ;
wire \us11/_0581_ ;
wire \us11/_0582_ ;
wire \us11/_0583_ ;
wire \us11/_0584_ ;
wire \us11/_0585_ ;
wire \us11/_0586_ ;
wire \us11/_0587_ ;
wire \us11/_0588_ ;
wire \us11/_0589_ ;
wire \us11/_0590_ ;
wire \us11/_0591_ ;
wire \us11/_0592_ ;
wire \us11/_0593_ ;
wire \us11/_0594_ ;
wire \us11/_0595_ ;
wire \us11/_0596_ ;
wire \us11/_0598_ ;
wire \us11/_0599_ ;
wire \us11/_0600_ ;
wire \us11/_0601_ ;
wire \us11/_0602_ ;
wire \us11/_0603_ ;
wire \us11/_0604_ ;
wire \us11/_0605_ ;
wire \us11/_0606_ ;
wire \us11/_0607_ ;
wire \us11/_0608_ ;
wire \us11/_0609_ ;
wire \us11/_0610_ ;
wire \us11/_0611_ ;
wire \us11/_0612_ ;
wire \us11/_0613_ ;
wire \us11/_0614_ ;
wire \us11/_0615_ ;
wire \us11/_0616_ ;
wire \us11/_0617_ ;
wire \us11/_0618_ ;
wire \us11/_0619_ ;
wire \us11/_0620_ ;
wire \us11/_0621_ ;
wire \us11/_0622_ ;
wire \us11/_0623_ ;
wire \us11/_0624_ ;
wire \us11/_0625_ ;
wire \us11/_0626_ ;
wire \us11/_0627_ ;
wire \us11/_0628_ ;
wire \us11/_0629_ ;
wire \us11/_0630_ ;
wire \us11/_0631_ ;
wire \us11/_0632_ ;
wire \us11/_0633_ ;
wire \us11/_0634_ ;
wire \us11/_0635_ ;
wire \us11/_0636_ ;
wire \us11/_0637_ ;
wire \us11/_0638_ ;
wire \us11/_0639_ ;
wire \us11/_0640_ ;
wire \us11/_0641_ ;
wire \us11/_0642_ ;
wire \us11/_0643_ ;
wire \us11/_0644_ ;
wire \us11/_0645_ ;
wire \us11/_0646_ ;
wire \us11/_0647_ ;
wire \us11/_0648_ ;
wire \us11/_0649_ ;
wire \us11/_0650_ ;
wire \us11/_0652_ ;
wire \us11/_0653_ ;
wire \us11/_0654_ ;
wire \us11/_0655_ ;
wire \us11/_0656_ ;
wire \us11/_0657_ ;
wire \us11/_0658_ ;
wire \us11/_0659_ ;
wire \us11/_0660_ ;
wire \us11/_0661_ ;
wire \us11/_0662_ ;
wire \us11/_0663_ ;
wire \us11/_0664_ ;
wire \us11/_0665_ ;
wire \us11/_0666_ ;
wire \us11/_0667_ ;
wire \us11/_0668_ ;
wire \us11/_0669_ ;
wire \us11/_0670_ ;
wire \us11/_0671_ ;
wire \us11/_0673_ ;
wire \us11/_0674_ ;
wire \us11/_0675_ ;
wire \us11/_0676_ ;
wire \us11/_0677_ ;
wire \us11/_0678_ ;
wire \us11/_0679_ ;
wire \us11/_0680_ ;
wire \us11/_0681_ ;
wire \us11/_0682_ ;
wire \us11/_0683_ ;
wire \us11/_0684_ ;
wire \us11/_0685_ ;
wire \us11/_0686_ ;
wire \us11/_0687_ ;
wire \us11/_0688_ ;
wire \us11/_0689_ ;
wire \us11/_0690_ ;
wire \us11/_0691_ ;
wire \us11/_0692_ ;
wire \us11/_0693_ ;
wire \us11/_0694_ ;
wire \us11/_0695_ ;
wire \us11/_0696_ ;
wire \us11/_0697_ ;
wire \us11/_0698_ ;
wire \us11/_0699_ ;
wire \us11/_0700_ ;
wire \us11/_0701_ ;
wire \us11/_0702_ ;
wire \us11/_0703_ ;
wire \us11/_0704_ ;
wire \us11/_0705_ ;
wire \us11/_0706_ ;
wire \us11/_0707_ ;
wire \us11/_0708_ ;
wire \us11/_0709_ ;
wire \us11/_0710_ ;
wire \us11/_0711_ ;
wire \us11/_0712_ ;
wire \us11/_0713_ ;
wire \us11/_0714_ ;
wire \us11/_0715_ ;
wire \us11/_0717_ ;
wire \us11/_0718_ ;
wire \us11/_0719_ ;
wire \us11/_0720_ ;
wire \us11/_0721_ ;
wire \us11/_0722_ ;
wire \us11/_0723_ ;
wire \us11/_0724_ ;
wire \us11/_0725_ ;
wire \us11/_0726_ ;
wire \us11/_0727_ ;
wire \us11/_0728_ ;
wire \us11/_0729_ ;
wire \us11/_0730_ ;
wire \us11/_0731_ ;
wire \us11/_0732_ ;
wire \us11/_0733_ ;
wire \us11/_0734_ ;
wire \us11/_0735_ ;
wire \us11/_0736_ ;
wire \us11/_0738_ ;
wire \us11/_0739_ ;
wire \us11/_0740_ ;
wire \us11/_0741_ ;
wire \us11/_0742_ ;
wire \us11/_0744_ ;
wire \us11/_0745_ ;
wire \us11/_0746_ ;
wire \us11/_0748_ ;
wire \us11/_0749_ ;
wire \us11/_0750_ ;
wire \us11/_0752_ ;
wire \us12/_0008_ ;
wire \us12/_0009_ ;
wire \us12/_0010_ ;
wire \us12/_0011_ ;
wire \us12/_0012_ ;
wire \us12/_0013_ ;
wire \us12/_0014_ ;
wire \us12/_0015_ ;
wire \us12/_0016_ ;
wire \us12/_0017_ ;
wire \us12/_0018_ ;
wire \us12/_0019_ ;
wire \us12/_0020_ ;
wire \us12/_0022_ ;
wire \us12/_0024_ ;
wire \us12/_0025_ ;
wire \us12/_0026_ ;
wire \us12/_0027_ ;
wire \us12/_0029_ ;
wire \us12/_0030_ ;
wire \us12/_0032_ ;
wire \us12/_0033_ ;
wire \us12/_0034_ ;
wire \us12/_0035_ ;
wire \us12/_0037_ ;
wire \us12/_0038_ ;
wire \us12/_0039_ ;
wire \us12/_0040_ ;
wire \us12/_0041_ ;
wire \us12/_0042_ ;
wire \us12/_0043_ ;
wire \us12/_0045_ ;
wire \us12/_0046_ ;
wire \us12/_0047_ ;
wire \us12/_0049_ ;
wire \us12/_0050_ ;
wire \us12/_0051_ ;
wire \us12/_0052_ ;
wire \us12/_0053_ ;
wire \us12/_0054_ ;
wire \us12/_0056_ ;
wire \us12/_0057_ ;
wire \us12/_0058_ ;
wire \us12/_0060_ ;
wire \us12/_0061_ ;
wire \us12/_0062_ ;
wire \us12/_0064_ ;
wire \us12/_0065_ ;
wire \us12/_0066_ ;
wire \us12/_0067_ ;
wire \us12/_0069_ ;
wire \us12/_0070_ ;
wire \us12/_0072_ ;
wire \us12/_0073_ ;
wire \us12/_0074_ ;
wire \us12/_0075_ ;
wire \us12/_0076_ ;
wire \us12/_0077_ ;
wire \us12/_0078_ ;
wire \us12/_0079_ ;
wire \us12/_0081_ ;
wire \us12/_0082_ ;
wire \us12/_0084_ ;
wire \us12/_0085_ ;
wire \us12/_0086_ ;
wire \us12/_0087_ ;
wire \us12/_0088_ ;
wire \us12/_0089_ ;
wire \us12/_0090_ ;
wire \us12/_0091_ ;
wire \us12/_0092_ ;
wire \us12/_0093_ ;
wire \us12/_0094_ ;
wire \us12/_0095_ ;
wire \us12/_0096_ ;
wire \us12/_0097_ ;
wire \us12/_0098_ ;
wire \us12/_0099_ ;
wire \us12/_0100_ ;
wire \us12/_0101_ ;
wire \us12/_0102_ ;
wire \us12/_0103_ ;
wire \us12/_0104_ ;
wire \us12/_0105_ ;
wire \us12/_0106_ ;
wire \us12/_0108_ ;
wire \us12/_0109_ ;
wire \us12/_0110_ ;
wire \us12/_0111_ ;
wire \us12/_0113_ ;
wire \us12/_0114_ ;
wire \us12/_0115_ ;
wire \us12/_0116_ ;
wire \us12/_0117_ ;
wire \us12/_0118_ ;
wire \us12/_0119_ ;
wire \us12/_0120_ ;
wire \us12/_0121_ ;
wire \us12/_0122_ ;
wire \us12/_0123_ ;
wire \us12/_0124_ ;
wire \us12/_0126_ ;
wire \us12/_0127_ ;
wire \us12/_0128_ ;
wire \us12/_0129_ ;
wire \us12/_0130_ ;
wire \us12/_0132_ ;
wire \us12/_0133_ ;
wire \us12/_0134_ ;
wire \us12/_0135_ ;
wire \us12/_0136_ ;
wire \us12/_0137_ ;
wire \us12/_0139_ ;
wire \us12/_0140_ ;
wire \us12/_0141_ ;
wire \us12/_0142_ ;
wire \us12/_0144_ ;
wire \us12/_0145_ ;
wire \us12/_0146_ ;
wire \us12/_0147_ ;
wire \us12/_0148_ ;
wire \us12/_0149_ ;
wire \us12/_0150_ ;
wire \us12/_0151_ ;
wire \us12/_0153_ ;
wire \us12/_0154_ ;
wire \us12/_0155_ ;
wire \us12/_0156_ ;
wire \us12/_0157_ ;
wire \us12/_0158_ ;
wire \us12/_0159_ ;
wire \us12/_0161_ ;
wire \us12/_0162_ ;
wire \us12/_0163_ ;
wire \us12/_0164_ ;
wire \us12/_0165_ ;
wire \us12/_0166_ ;
wire \us12/_0167_ ;
wire \us12/_0168_ ;
wire \us12/_0169_ ;
wire \us12/_0170_ ;
wire \us12/_0171_ ;
wire \us12/_0172_ ;
wire \us12/_0174_ ;
wire \us12/_0175_ ;
wire \us12/_0176_ ;
wire \us12/_0177_ ;
wire \us12/_0178_ ;
wire \us12/_0179_ ;
wire \us12/_0180_ ;
wire \us12/_0181_ ;
wire \us12/_0182_ ;
wire \us12/_0183_ ;
wire \us12/_0184_ ;
wire \us12/_0185_ ;
wire \us12/_0186_ ;
wire \us12/_0187_ ;
wire \us12/_0188_ ;
wire \us12/_0189_ ;
wire \us12/_0190_ ;
wire \us12/_0191_ ;
wire \us12/_0192_ ;
wire \us12/_0193_ ;
wire \us12/_0194_ ;
wire \us12/_0195_ ;
wire \us12/_0196_ ;
wire \us12/_0197_ ;
wire \us12/_0198_ ;
wire \us12/_0199_ ;
wire \us12/_0200_ ;
wire \us12/_0201_ ;
wire \us12/_0202_ ;
wire \us12/_0203_ ;
wire \us12/_0204_ ;
wire \us12/_0205_ ;
wire \us12/_0206_ ;
wire \us12/_0207_ ;
wire \us12/_0208_ ;
wire \us12/_0209_ ;
wire \us12/_0210_ ;
wire \us12/_0211_ ;
wire \us12/_0212_ ;
wire \us12/_0213_ ;
wire \us12/_0214_ ;
wire \us12/_0215_ ;
wire \us12/_0216_ ;
wire \us12/_0217_ ;
wire \us12/_0219_ ;
wire \us12/_0220_ ;
wire \us12/_0221_ ;
wire \us12/_0222_ ;
wire \us12/_0223_ ;
wire \us12/_0224_ ;
wire \us12/_0225_ ;
wire \us12/_0226_ ;
wire \us12/_0227_ ;
wire \us12/_0228_ ;
wire \us12/_0229_ ;
wire \us12/_0230_ ;
wire \us12/_0231_ ;
wire \us12/_0232_ ;
wire \us12/_0233_ ;
wire \us12/_0234_ ;
wire \us12/_0235_ ;
wire \us12/_0236_ ;
wire \us12/_0237_ ;
wire \us12/_0238_ ;
wire \us12/_0239_ ;
wire \us12/_0240_ ;
wire \us12/_0241_ ;
wire \us12/_0242_ ;
wire \us12/_0243_ ;
wire \us12/_0244_ ;
wire \us12/_0245_ ;
wire \us12/_0246_ ;
wire \us12/_0248_ ;
wire \us12/_0249_ ;
wire \us12/_0250_ ;
wire \us12/_0251_ ;
wire \us12/_0252_ ;
wire \us12/_0253_ ;
wire \us12/_0254_ ;
wire \us12/_0255_ ;
wire \us12/_0256_ ;
wire \us12/_0257_ ;
wire \us12/_0258_ ;
wire \us12/_0259_ ;
wire \us12/_0260_ ;
wire \us12/_0261_ ;
wire \us12/_0263_ ;
wire \us12/_0264_ ;
wire \us12/_0265_ ;
wire \us12/_0266_ ;
wire \us12/_0267_ ;
wire \us12/_0268_ ;
wire \us12/_0269_ ;
wire \us12/_0270_ ;
wire \us12/_0271_ ;
wire \us12/_0272_ ;
wire \us12/_0273_ ;
wire \us12/_0274_ ;
wire \us12/_0275_ ;
wire \us12/_0276_ ;
wire \us12/_0277_ ;
wire \us12/_0278_ ;
wire \us12/_0279_ ;
wire \us12/_0281_ ;
wire \us12/_0283_ ;
wire \us12/_0284_ ;
wire \us12/_0285_ ;
wire \us12/_0286_ ;
wire \us12/_0287_ ;
wire \us12/_0288_ ;
wire \us12/_0289_ ;
wire \us12/_0290_ ;
wire \us12/_0291_ ;
wire \us12/_0293_ ;
wire \us12/_0294_ ;
wire \us12/_0295_ ;
wire \us12/_0296_ ;
wire \us12/_0297_ ;
wire \us12/_0298_ ;
wire \us12/_0299_ ;
wire \us12/_0300_ ;
wire \us12/_0301_ ;
wire \us12/_0302_ ;
wire \us12/_0303_ ;
wire \us12/_0304_ ;
wire \us12/_0305_ ;
wire \us12/_0306_ ;
wire \us12/_0307_ ;
wire \us12/_0308_ ;
wire \us12/_0309_ ;
wire \us12/_0310_ ;
wire \us12/_0311_ ;
wire \us12/_0312_ ;
wire \us12/_0313_ ;
wire \us12/_0314_ ;
wire \us12/_0315_ ;
wire \us12/_0316_ ;
wire \us12/_0317_ ;
wire \us12/_0318_ ;
wire \us12/_0319_ ;
wire \us12/_0320_ ;
wire \us12/_0321_ ;
wire \us12/_0322_ ;
wire \us12/_0323_ ;
wire \us12/_0324_ ;
wire \us12/_0325_ ;
wire \us12/_0326_ ;
wire \us12/_0327_ ;
wire \us12/_0328_ ;
wire \us12/_0329_ ;
wire \us12/_0330_ ;
wire \us12/_0331_ ;
wire \us12/_0332_ ;
wire \us12/_0333_ ;
wire \us12/_0334_ ;
wire \us12/_0335_ ;
wire \us12/_0337_ ;
wire \us12/_0338_ ;
wire \us12/_0339_ ;
wire \us12/_0340_ ;
wire \us12/_0341_ ;
wire \us12/_0342_ ;
wire \us12/_0343_ ;
wire \us12/_0344_ ;
wire \us12/_0345_ ;
wire \us12/_0347_ ;
wire \us12/_0348_ ;
wire \us12/_0349_ ;
wire \us12/_0350_ ;
wire \us12/_0351_ ;
wire \us12/_0352_ ;
wire \us12/_0353_ ;
wire \us12/_0354_ ;
wire \us12/_0355_ ;
wire \us12/_0356_ ;
wire \us12/_0357_ ;
wire \us12/_0358_ ;
wire \us12/_0359_ ;
wire \us12/_0360_ ;
wire \us12/_0361_ ;
wire \us12/_0362_ ;
wire \us12/_0363_ ;
wire \us12/_0365_ ;
wire \us12/_0366_ ;
wire \us12/_0367_ ;
wire \us12/_0368_ ;
wire \us12/_0370_ ;
wire \us12/_0371_ ;
wire \us12/_0372_ ;
wire \us12/_0373_ ;
wire \us12/_0374_ ;
wire \us12/_0375_ ;
wire \us12/_0376_ ;
wire \us12/_0377_ ;
wire \us12/_0378_ ;
wire \us12/_0379_ ;
wire \us12/_0380_ ;
wire \us12/_0381_ ;
wire \us12/_0382_ ;
wire \us12/_0383_ ;
wire \us12/_0384_ ;
wire \us12/_0385_ ;
wire \us12/_0386_ ;
wire \us12/_0387_ ;
wire \us12/_0388_ ;
wire \us12/_0389_ ;
wire \us12/_0390_ ;
wire \us12/_0391_ ;
wire \us12/_0392_ ;
wire \us12/_0393_ ;
wire \us12/_0394_ ;
wire \us12/_0395_ ;
wire \us12/_0396_ ;
wire \us12/_0397_ ;
wire \us12/_0398_ ;
wire \us12/_0399_ ;
wire \us12/_0400_ ;
wire \us12/_0401_ ;
wire \us12/_0402_ ;
wire \us12/_0403_ ;
wire \us12/_0404_ ;
wire \us12/_0405_ ;
wire \us12/_0406_ ;
wire \us12/_0407_ ;
wire \us12/_0408_ ;
wire \us12/_0409_ ;
wire \us12/_0410_ ;
wire \us12/_0411_ ;
wire \us12/_0412_ ;
wire \us12/_0413_ ;
wire \us12/_0414_ ;
wire \us12/_0415_ ;
wire \us12/_0416_ ;
wire \us12/_0417_ ;
wire \us12/_0418_ ;
wire \us12/_0419_ ;
wire \us12/_0420_ ;
wire \us12/_0421_ ;
wire \us12/_0422_ ;
wire \us12/_0423_ ;
wire \us12/_0424_ ;
wire \us12/_0425_ ;
wire \us12/_0426_ ;
wire \us12/_0427_ ;
wire \us12/_0428_ ;
wire \us12/_0429_ ;
wire \us12/_0430_ ;
wire \us12/_0431_ ;
wire \us12/_0432_ ;
wire \us12/_0433_ ;
wire \us12/_0434_ ;
wire \us12/_0435_ ;
wire \us12/_0436_ ;
wire \us12/_0437_ ;
wire \us12/_0438_ ;
wire \us12/_0439_ ;
wire \us12/_0440_ ;
wire \us12/_0441_ ;
wire \us12/_0442_ ;
wire \us12/_0443_ ;
wire \us12/_0444_ ;
wire \us12/_0446_ ;
wire \us12/_0447_ ;
wire \us12/_0448_ ;
wire \us12/_0449_ ;
wire \us12/_0450_ ;
wire \us12/_0451_ ;
wire \us12/_0452_ ;
wire \us12/_0453_ ;
wire \us12/_0454_ ;
wire \us12/_0455_ ;
wire \us12/_0457_ ;
wire \us12/_0458_ ;
wire \us12/_0459_ ;
wire \us12/_0460_ ;
wire \us12/_0461_ ;
wire \us12/_0462_ ;
wire \us12/_0463_ ;
wire \us12/_0464_ ;
wire \us12/_0465_ ;
wire \us12/_0466_ ;
wire \us12/_0467_ ;
wire \us12/_0468_ ;
wire \us12/_0469_ ;
wire \us12/_0470_ ;
wire \us12/_0471_ ;
wire \us12/_0472_ ;
wire \us12/_0473_ ;
wire \us12/_0474_ ;
wire \us12/_0475_ ;
wire \us12/_0476_ ;
wire \us12/_0477_ ;
wire \us12/_0478_ ;
wire \us12/_0479_ ;
wire \us12/_0480_ ;
wire \us12/_0481_ ;
wire \us12/_0482_ ;
wire \us12/_0483_ ;
wire \us12/_0484_ ;
wire \us12/_0485_ ;
wire \us12/_0486_ ;
wire \us12/_0487_ ;
wire \us12/_0488_ ;
wire \us12/_0489_ ;
wire \us12/_0490_ ;
wire \us12/_0491_ ;
wire \us12/_0492_ ;
wire \us12/_0493_ ;
wire \us12/_0494_ ;
wire \us12/_0495_ ;
wire \us12/_0496_ ;
wire \us12/_0497_ ;
wire \us12/_0498_ ;
wire \us12/_0499_ ;
wire \us12/_0500_ ;
wire \us12/_0501_ ;
wire \us12/_0502_ ;
wire \us12/_0503_ ;
wire \us12/_0504_ ;
wire \us12/_0505_ ;
wire \us12/_0506_ ;
wire \us12/_0507_ ;
wire \us12/_0508_ ;
wire \us12/_0509_ ;
wire \us12/_0510_ ;
wire \us12/_0511_ ;
wire \us12/_0512_ ;
wire \us12/_0513_ ;
wire \us12/_0514_ ;
wire \us12/_0515_ ;
wire \us12/_0516_ ;
wire \us12/_0517_ ;
wire \us12/_0518_ ;
wire \us12/_0519_ ;
wire \us12/_0520_ ;
wire \us12/_0521_ ;
wire \us12/_0522_ ;
wire \us12/_0523_ ;
wire \us12/_0524_ ;
wire \us12/_0525_ ;
wire \us12/_0526_ ;
wire \us12/_0527_ ;
wire \us12/_0528_ ;
wire \us12/_0529_ ;
wire \us12/_0530_ ;
wire \us12/_0531_ ;
wire \us12/_0532_ ;
wire \us12/_0533_ ;
wire \us12/_0534_ ;
wire \us12/_0535_ ;
wire \us12/_0536_ ;
wire \us12/_0537_ ;
wire \us12/_0538_ ;
wire \us12/_0539_ ;
wire \us12/_0540_ ;
wire \us12/_0541_ ;
wire \us12/_0542_ ;
wire \us12/_0543_ ;
wire \us12/_0544_ ;
wire \us12/_0545_ ;
wire \us12/_0546_ ;
wire \us12/_0547_ ;
wire \us12/_0548_ ;
wire \us12/_0549_ ;
wire \us12/_0550_ ;
wire \us12/_0551_ ;
wire \us12/_0552_ ;
wire \us12/_0553_ ;
wire \us12/_0554_ ;
wire \us12/_0555_ ;
wire \us12/_0556_ ;
wire \us12/_0557_ ;
wire \us12/_0558_ ;
wire \us12/_0559_ ;
wire \us12/_0560_ ;
wire \us12/_0561_ ;
wire \us12/_0562_ ;
wire \us12/_0563_ ;
wire \us12/_0565_ ;
wire \us12/_0566_ ;
wire \us12/_0567_ ;
wire \us12/_0568_ ;
wire \us12/_0569_ ;
wire \us12/_0570_ ;
wire \us12/_0571_ ;
wire \us12/_0572_ ;
wire \us12/_0573_ ;
wire \us12/_0574_ ;
wire \us12/_0575_ ;
wire \us12/_0576_ ;
wire \us12/_0577_ ;
wire \us12/_0578_ ;
wire \us12/_0579_ ;
wire \us12/_0580_ ;
wire \us12/_0581_ ;
wire \us12/_0582_ ;
wire \us12/_0583_ ;
wire \us12/_0584_ ;
wire \us12/_0585_ ;
wire \us12/_0586_ ;
wire \us12/_0587_ ;
wire \us12/_0588_ ;
wire \us12/_0589_ ;
wire \us12/_0590_ ;
wire \us12/_0591_ ;
wire \us12/_0592_ ;
wire \us12/_0593_ ;
wire \us12/_0594_ ;
wire \us12/_0595_ ;
wire \us12/_0596_ ;
wire \us12/_0598_ ;
wire \us12/_0599_ ;
wire \us12/_0600_ ;
wire \us12/_0601_ ;
wire \us12/_0602_ ;
wire \us12/_0603_ ;
wire \us12/_0604_ ;
wire \us12/_0605_ ;
wire \us12/_0606_ ;
wire \us12/_0607_ ;
wire \us12/_0608_ ;
wire \us12/_0609_ ;
wire \us12/_0610_ ;
wire \us12/_0611_ ;
wire \us12/_0612_ ;
wire \us12/_0613_ ;
wire \us12/_0614_ ;
wire \us12/_0615_ ;
wire \us12/_0616_ ;
wire \us12/_0617_ ;
wire \us12/_0618_ ;
wire \us12/_0619_ ;
wire \us12/_0620_ ;
wire \us12/_0621_ ;
wire \us12/_0622_ ;
wire \us12/_0623_ ;
wire \us12/_0624_ ;
wire \us12/_0625_ ;
wire \us12/_0626_ ;
wire \us12/_0627_ ;
wire \us12/_0628_ ;
wire \us12/_0629_ ;
wire \us12/_0630_ ;
wire \us12/_0631_ ;
wire \us12/_0632_ ;
wire \us12/_0633_ ;
wire \us12/_0634_ ;
wire \us12/_0635_ ;
wire \us12/_0636_ ;
wire \us12/_0637_ ;
wire \us12/_0638_ ;
wire \us12/_0639_ ;
wire \us12/_0640_ ;
wire \us12/_0641_ ;
wire \us12/_0642_ ;
wire \us12/_0643_ ;
wire \us12/_0644_ ;
wire \us12/_0645_ ;
wire \us12/_0646_ ;
wire \us12/_0647_ ;
wire \us12/_0648_ ;
wire \us12/_0649_ ;
wire \us12/_0650_ ;
wire \us12/_0652_ ;
wire \us12/_0653_ ;
wire \us12/_0654_ ;
wire \us12/_0655_ ;
wire \us12/_0656_ ;
wire \us12/_0657_ ;
wire \us12/_0658_ ;
wire \us12/_0659_ ;
wire \us12/_0660_ ;
wire \us12/_0661_ ;
wire \us12/_0662_ ;
wire \us12/_0663_ ;
wire \us12/_0664_ ;
wire \us12/_0665_ ;
wire \us12/_0666_ ;
wire \us12/_0667_ ;
wire \us12/_0668_ ;
wire \us12/_0669_ ;
wire \us12/_0670_ ;
wire \us12/_0671_ ;
wire \us12/_0673_ ;
wire \us12/_0674_ ;
wire \us12/_0675_ ;
wire \us12/_0676_ ;
wire \us12/_0677_ ;
wire \us12/_0678_ ;
wire \us12/_0679_ ;
wire \us12/_0680_ ;
wire \us12/_0681_ ;
wire \us12/_0682_ ;
wire \us12/_0683_ ;
wire \us12/_0684_ ;
wire \us12/_0685_ ;
wire \us12/_0686_ ;
wire \us12/_0687_ ;
wire \us12/_0688_ ;
wire \us12/_0689_ ;
wire \us12/_0690_ ;
wire \us12/_0691_ ;
wire \us12/_0692_ ;
wire \us12/_0693_ ;
wire \us12/_0694_ ;
wire \us12/_0695_ ;
wire \us12/_0696_ ;
wire \us12/_0697_ ;
wire \us12/_0698_ ;
wire \us12/_0699_ ;
wire \us12/_0700_ ;
wire \us12/_0701_ ;
wire \us12/_0702_ ;
wire \us12/_0703_ ;
wire \us12/_0704_ ;
wire \us12/_0705_ ;
wire \us12/_0706_ ;
wire \us12/_0707_ ;
wire \us12/_0708_ ;
wire \us12/_0709_ ;
wire \us12/_0710_ ;
wire \us12/_0711_ ;
wire \us12/_0712_ ;
wire \us12/_0713_ ;
wire \us12/_0714_ ;
wire \us12/_0715_ ;
wire \us12/_0717_ ;
wire \us12/_0718_ ;
wire \us12/_0719_ ;
wire \us12/_0720_ ;
wire \us12/_0721_ ;
wire \us12/_0722_ ;
wire \us12/_0723_ ;
wire \us12/_0724_ ;
wire \us12/_0725_ ;
wire \us12/_0726_ ;
wire \us12/_0727_ ;
wire \us12/_0728_ ;
wire \us12/_0729_ ;
wire \us12/_0730_ ;
wire \us12/_0731_ ;
wire \us12/_0732_ ;
wire \us12/_0733_ ;
wire \us12/_0734_ ;
wire \us12/_0735_ ;
wire \us12/_0736_ ;
wire \us12/_0738_ ;
wire \us12/_0739_ ;
wire \us12/_0740_ ;
wire \us12/_0741_ ;
wire \us12/_0742_ ;
wire \us12/_0744_ ;
wire \us12/_0745_ ;
wire \us12/_0746_ ;
wire \us12/_0747_ ;
wire \us12/_0748_ ;
wire \us12/_0749_ ;
wire \us12/_0750_ ;
wire \us12/_0752_ ;
wire \us13/_0008_ ;
wire \us13/_0009_ ;
wire \us13/_0010_ ;
wire \us13/_0011_ ;
wire \us13/_0012_ ;
wire \us13/_0013_ ;
wire \us13/_0014_ ;
wire \us13/_0015_ ;
wire \us13/_0016_ ;
wire \us13/_0017_ ;
wire \us13/_0018_ ;
wire \us13/_0019_ ;
wire \us13/_0020_ ;
wire \us13/_0022_ ;
wire \us13/_0024_ ;
wire \us13/_0025_ ;
wire \us13/_0026_ ;
wire \us13/_0027_ ;
wire \us13/_0029_ ;
wire \us13/_0030_ ;
wire \us13/_0032_ ;
wire \us13/_0033_ ;
wire \us13/_0034_ ;
wire \us13/_0035_ ;
wire \us13/_0036_ ;
wire \us13/_0037_ ;
wire \us13/_0038_ ;
wire \us13/_0039_ ;
wire \us13/_0040_ ;
wire \us13/_0041_ ;
wire \us13/_0042_ ;
wire \us13/_0043_ ;
wire \us13/_0045_ ;
wire \us13/_0046_ ;
wire \us13/_0047_ ;
wire \us13/_0048_ ;
wire \us13/_0049_ ;
wire \us13/_0050_ ;
wire \us13/_0051_ ;
wire \us13/_0052_ ;
wire \us13/_0053_ ;
wire \us13/_0054_ ;
wire \us13/_0056_ ;
wire \us13/_0057_ ;
wire \us13/_0058_ ;
wire \us13/_0060_ ;
wire \us13/_0061_ ;
wire \us13/_0062_ ;
wire \us13/_0064_ ;
wire \us13/_0065_ ;
wire \us13/_0066_ ;
wire \us13/_0067_ ;
wire \us13/_0069_ ;
wire \us13/_0070_ ;
wire \us13/_0072_ ;
wire \us13/_0073_ ;
wire \us13/_0074_ ;
wire \us13/_0075_ ;
wire \us13/_0076_ ;
wire \us13/_0077_ ;
wire \us13/_0078_ ;
wire \us13/_0079_ ;
wire \us13/_0081_ ;
wire \us13/_0082_ ;
wire \us13/_0083_ ;
wire \us13/_0084_ ;
wire \us13/_0085_ ;
wire \us13/_0086_ ;
wire \us13/_0087_ ;
wire \us13/_0088_ ;
wire \us13/_0089_ ;
wire \us13/_0090_ ;
wire \us13/_0091_ ;
wire \us13/_0092_ ;
wire \us13/_0093_ ;
wire \us13/_0094_ ;
wire \us13/_0095_ ;
wire \us13/_0096_ ;
wire \us13/_0097_ ;
wire \us13/_0098_ ;
wire \us13/_0099_ ;
wire \us13/_0100_ ;
wire \us13/_0101_ ;
wire \us13/_0102_ ;
wire \us13/_0103_ ;
wire \us13/_0104_ ;
wire \us13/_0105_ ;
wire \us13/_0106_ ;
wire \us13/_0108_ ;
wire \us13/_0109_ ;
wire \us13/_0110_ ;
wire \us13/_0111_ ;
wire \us13/_0113_ ;
wire \us13/_0114_ ;
wire \us13/_0115_ ;
wire \us13/_0116_ ;
wire \us13/_0117_ ;
wire \us13/_0118_ ;
wire \us13/_0119_ ;
wire \us13/_0120_ ;
wire \us13/_0121_ ;
wire \us13/_0122_ ;
wire \us13/_0123_ ;
wire \us13/_0124_ ;
wire \us13/_0126_ ;
wire \us13/_0127_ ;
wire \us13/_0128_ ;
wire \us13/_0129_ ;
wire \us13/_0130_ ;
wire \us13/_0132_ ;
wire \us13/_0133_ ;
wire \us13/_0134_ ;
wire \us13/_0135_ ;
wire \us13/_0136_ ;
wire \us13/_0137_ ;
wire \us13/_0139_ ;
wire \us13/_0140_ ;
wire \us13/_0141_ ;
wire \us13/_0142_ ;
wire \us13/_0144_ ;
wire \us13/_0145_ ;
wire \us13/_0146_ ;
wire \us13/_0147_ ;
wire \us13/_0148_ ;
wire \us13/_0149_ ;
wire \us13/_0150_ ;
wire \us13/_0151_ ;
wire \us13/_0153_ ;
wire \us13/_0154_ ;
wire \us13/_0155_ ;
wire \us13/_0156_ ;
wire \us13/_0157_ ;
wire \us13/_0158_ ;
wire \us13/_0159_ ;
wire \us13/_0161_ ;
wire \us13/_0162_ ;
wire \us13/_0163_ ;
wire \us13/_0164_ ;
wire \us13/_0165_ ;
wire \us13/_0166_ ;
wire \us13/_0167_ ;
wire \us13/_0168_ ;
wire \us13/_0169_ ;
wire \us13/_0170_ ;
wire \us13/_0171_ ;
wire \us13/_0172_ ;
wire \us13/_0174_ ;
wire \us13/_0175_ ;
wire \us13/_0176_ ;
wire \us13/_0177_ ;
wire \us13/_0178_ ;
wire \us13/_0179_ ;
wire \us13/_0180_ ;
wire \us13/_0181_ ;
wire \us13/_0182_ ;
wire \us13/_0183_ ;
wire \us13/_0184_ ;
wire \us13/_0185_ ;
wire \us13/_0186_ ;
wire \us13/_0187_ ;
wire \us13/_0188_ ;
wire \us13/_0189_ ;
wire \us13/_0190_ ;
wire \us13/_0191_ ;
wire \us13/_0192_ ;
wire \us13/_0193_ ;
wire \us13/_0194_ ;
wire \us13/_0195_ ;
wire \us13/_0196_ ;
wire \us13/_0197_ ;
wire \us13/_0198_ ;
wire \us13/_0199_ ;
wire \us13/_0200_ ;
wire \us13/_0201_ ;
wire \us13/_0202_ ;
wire \us13/_0203_ ;
wire \us13/_0204_ ;
wire \us13/_0205_ ;
wire \us13/_0206_ ;
wire \us13/_0207_ ;
wire \us13/_0208_ ;
wire \us13/_0209_ ;
wire \us13/_0210_ ;
wire \us13/_0211_ ;
wire \us13/_0212_ ;
wire \us13/_0213_ ;
wire \us13/_0214_ ;
wire \us13/_0215_ ;
wire \us13/_0216_ ;
wire \us13/_0217_ ;
wire \us13/_0219_ ;
wire \us13/_0220_ ;
wire \us13/_0221_ ;
wire \us13/_0222_ ;
wire \us13/_0223_ ;
wire \us13/_0224_ ;
wire \us13/_0225_ ;
wire \us13/_0226_ ;
wire \us13/_0227_ ;
wire \us13/_0228_ ;
wire \us13/_0229_ ;
wire \us13/_0230_ ;
wire \us13/_0231_ ;
wire \us13/_0232_ ;
wire \us13/_0233_ ;
wire \us13/_0234_ ;
wire \us13/_0235_ ;
wire \us13/_0236_ ;
wire \us13/_0237_ ;
wire \us13/_0238_ ;
wire \us13/_0239_ ;
wire \us13/_0240_ ;
wire \us13/_0241_ ;
wire \us13/_0242_ ;
wire \us13/_0243_ ;
wire \us13/_0244_ ;
wire \us13/_0245_ ;
wire \us13/_0246_ ;
wire \us13/_0248_ ;
wire \us13/_0249_ ;
wire \us13/_0250_ ;
wire \us13/_0251_ ;
wire \us13/_0252_ ;
wire \us13/_0253_ ;
wire \us13/_0254_ ;
wire \us13/_0255_ ;
wire \us13/_0256_ ;
wire \us13/_0257_ ;
wire \us13/_0258_ ;
wire \us13/_0259_ ;
wire \us13/_0260_ ;
wire \us13/_0261_ ;
wire \us13/_0263_ ;
wire \us13/_0264_ ;
wire \us13/_0265_ ;
wire \us13/_0266_ ;
wire \us13/_0267_ ;
wire \us13/_0268_ ;
wire \us13/_0269_ ;
wire \us13/_0270_ ;
wire \us13/_0271_ ;
wire \us13/_0272_ ;
wire \us13/_0273_ ;
wire \us13/_0274_ ;
wire \us13/_0275_ ;
wire \us13/_0276_ ;
wire \us13/_0277_ ;
wire \us13/_0278_ ;
wire \us13/_0279_ ;
wire \us13/_0281_ ;
wire \us13/_0283_ ;
wire \us13/_0284_ ;
wire \us13/_0285_ ;
wire \us13/_0286_ ;
wire \us13/_0287_ ;
wire \us13/_0288_ ;
wire \us13/_0289_ ;
wire \us13/_0290_ ;
wire \us13/_0291_ ;
wire \us13/_0293_ ;
wire \us13/_0294_ ;
wire \us13/_0295_ ;
wire \us13/_0296_ ;
wire \us13/_0297_ ;
wire \us13/_0298_ ;
wire \us13/_0299_ ;
wire \us13/_0300_ ;
wire \us13/_0301_ ;
wire \us13/_0302_ ;
wire \us13/_0303_ ;
wire \us13/_0304_ ;
wire \us13/_0305_ ;
wire \us13/_0306_ ;
wire \us13/_0307_ ;
wire \us13/_0308_ ;
wire \us13/_0309_ ;
wire \us13/_0310_ ;
wire \us13/_0311_ ;
wire \us13/_0312_ ;
wire \us13/_0313_ ;
wire \us13/_0314_ ;
wire \us13/_0315_ ;
wire \us13/_0316_ ;
wire \us13/_0317_ ;
wire \us13/_0318_ ;
wire \us13/_0319_ ;
wire \us13/_0320_ ;
wire \us13/_0321_ ;
wire \us13/_0322_ ;
wire \us13/_0323_ ;
wire \us13/_0324_ ;
wire \us13/_0325_ ;
wire \us13/_0326_ ;
wire \us13/_0327_ ;
wire \us13/_0328_ ;
wire \us13/_0329_ ;
wire \us13/_0330_ ;
wire \us13/_0331_ ;
wire \us13/_0332_ ;
wire \us13/_0333_ ;
wire \us13/_0334_ ;
wire \us13/_0335_ ;
wire \us13/_0337_ ;
wire \us13/_0338_ ;
wire \us13/_0339_ ;
wire \us13/_0340_ ;
wire \us13/_0341_ ;
wire \us13/_0342_ ;
wire \us13/_0343_ ;
wire \us13/_0344_ ;
wire \us13/_0345_ ;
wire \us13/_0347_ ;
wire \us13/_0348_ ;
wire \us13/_0349_ ;
wire \us13/_0350_ ;
wire \us13/_0351_ ;
wire \us13/_0352_ ;
wire \us13/_0353_ ;
wire \us13/_0354_ ;
wire \us13/_0355_ ;
wire \us13/_0356_ ;
wire \us13/_0357_ ;
wire \us13/_0358_ ;
wire \us13/_0359_ ;
wire \us13/_0360_ ;
wire \us13/_0361_ ;
wire \us13/_0362_ ;
wire \us13/_0363_ ;
wire \us13/_0365_ ;
wire \us13/_0366_ ;
wire \us13/_0367_ ;
wire \us13/_0368_ ;
wire \us13/_0370_ ;
wire \us13/_0371_ ;
wire \us13/_0372_ ;
wire \us13/_0373_ ;
wire \us13/_0374_ ;
wire \us13/_0375_ ;
wire \us13/_0376_ ;
wire \us13/_0377_ ;
wire \us13/_0378_ ;
wire \us13/_0379_ ;
wire \us13/_0380_ ;
wire \us13/_0381_ ;
wire \us13/_0382_ ;
wire \us13/_0383_ ;
wire \us13/_0384_ ;
wire \us13/_0385_ ;
wire \us13/_0386_ ;
wire \us13/_0387_ ;
wire \us13/_0388_ ;
wire \us13/_0389_ ;
wire \us13/_0390_ ;
wire \us13/_0391_ ;
wire \us13/_0392_ ;
wire \us13/_0393_ ;
wire \us13/_0394_ ;
wire \us13/_0395_ ;
wire \us13/_0396_ ;
wire \us13/_0397_ ;
wire \us13/_0398_ ;
wire \us13/_0399_ ;
wire \us13/_0400_ ;
wire \us13/_0401_ ;
wire \us13/_0402_ ;
wire \us13/_0403_ ;
wire \us13/_0404_ ;
wire \us13/_0405_ ;
wire \us13/_0406_ ;
wire \us13/_0407_ ;
wire \us13/_0408_ ;
wire \us13/_0409_ ;
wire \us13/_0410_ ;
wire \us13/_0411_ ;
wire \us13/_0412_ ;
wire \us13/_0413_ ;
wire \us13/_0414_ ;
wire \us13/_0415_ ;
wire \us13/_0416_ ;
wire \us13/_0417_ ;
wire \us13/_0418_ ;
wire \us13/_0419_ ;
wire \us13/_0420_ ;
wire \us13/_0421_ ;
wire \us13/_0422_ ;
wire \us13/_0423_ ;
wire \us13/_0424_ ;
wire \us13/_0425_ ;
wire \us13/_0426_ ;
wire \us13/_0427_ ;
wire \us13/_0428_ ;
wire \us13/_0429_ ;
wire \us13/_0430_ ;
wire \us13/_0431_ ;
wire \us13/_0432_ ;
wire \us13/_0433_ ;
wire \us13/_0434_ ;
wire \us13/_0435_ ;
wire \us13/_0436_ ;
wire \us13/_0437_ ;
wire \us13/_0438_ ;
wire \us13/_0439_ ;
wire \us13/_0440_ ;
wire \us13/_0441_ ;
wire \us13/_0442_ ;
wire \us13/_0443_ ;
wire \us13/_0444_ ;
wire \us13/_0446_ ;
wire \us13/_0447_ ;
wire \us13/_0448_ ;
wire \us13/_0449_ ;
wire \us13/_0450_ ;
wire \us13/_0451_ ;
wire \us13/_0452_ ;
wire \us13/_0453_ ;
wire \us13/_0454_ ;
wire \us13/_0455_ ;
wire \us13/_0457_ ;
wire \us13/_0458_ ;
wire \us13/_0459_ ;
wire \us13/_0460_ ;
wire \us13/_0461_ ;
wire \us13/_0462_ ;
wire \us13/_0463_ ;
wire \us13/_0464_ ;
wire \us13/_0465_ ;
wire \us13/_0466_ ;
wire \us13/_0467_ ;
wire \us13/_0468_ ;
wire \us13/_0469_ ;
wire \us13/_0470_ ;
wire \us13/_0471_ ;
wire \us13/_0472_ ;
wire \us13/_0473_ ;
wire \us13/_0474_ ;
wire \us13/_0475_ ;
wire \us13/_0476_ ;
wire \us13/_0477_ ;
wire \us13/_0478_ ;
wire \us13/_0479_ ;
wire \us13/_0480_ ;
wire \us13/_0481_ ;
wire \us13/_0482_ ;
wire \us13/_0483_ ;
wire \us13/_0484_ ;
wire \us13/_0485_ ;
wire \us13/_0486_ ;
wire \us13/_0487_ ;
wire \us13/_0488_ ;
wire \us13/_0490_ ;
wire \us13/_0491_ ;
wire \us13/_0492_ ;
wire \us13/_0493_ ;
wire \us13/_0494_ ;
wire \us13/_0495_ ;
wire \us13/_0496_ ;
wire \us13/_0497_ ;
wire \us13/_0498_ ;
wire \us13/_0499_ ;
wire \us13/_0500_ ;
wire \us13/_0501_ ;
wire \us13/_0502_ ;
wire \us13/_0503_ ;
wire \us13/_0504_ ;
wire \us13/_0505_ ;
wire \us13/_0506_ ;
wire \us13/_0507_ ;
wire \us13/_0508_ ;
wire \us13/_0509_ ;
wire \us13/_0510_ ;
wire \us13/_0511_ ;
wire \us13/_0512_ ;
wire \us13/_0513_ ;
wire \us13/_0514_ ;
wire \us13/_0515_ ;
wire \us13/_0516_ ;
wire \us13/_0517_ ;
wire \us13/_0518_ ;
wire \us13/_0519_ ;
wire \us13/_0520_ ;
wire \us13/_0521_ ;
wire \us13/_0522_ ;
wire \us13/_0523_ ;
wire \us13/_0524_ ;
wire \us13/_0525_ ;
wire \us13/_0526_ ;
wire \us13/_0527_ ;
wire \us13/_0528_ ;
wire \us13/_0529_ ;
wire \us13/_0530_ ;
wire \us13/_0531_ ;
wire \us13/_0532_ ;
wire \us13/_0533_ ;
wire \us13/_0534_ ;
wire \us13/_0535_ ;
wire \us13/_0536_ ;
wire \us13/_0537_ ;
wire \us13/_0538_ ;
wire \us13/_0539_ ;
wire \us13/_0540_ ;
wire \us13/_0541_ ;
wire \us13/_0542_ ;
wire \us13/_0543_ ;
wire \us13/_0544_ ;
wire \us13/_0545_ ;
wire \us13/_0546_ ;
wire \us13/_0547_ ;
wire \us13/_0548_ ;
wire \us13/_0549_ ;
wire \us13/_0550_ ;
wire \us13/_0551_ ;
wire \us13/_0552_ ;
wire \us13/_0553_ ;
wire \us13/_0554_ ;
wire \us13/_0555_ ;
wire \us13/_0556_ ;
wire \us13/_0557_ ;
wire \us13/_0558_ ;
wire \us13/_0559_ ;
wire \us13/_0560_ ;
wire \us13/_0561_ ;
wire \us13/_0562_ ;
wire \us13/_0563_ ;
wire \us13/_0565_ ;
wire \us13/_0566_ ;
wire \us13/_0567_ ;
wire \us13/_0568_ ;
wire \us13/_0569_ ;
wire \us13/_0570_ ;
wire \us13/_0571_ ;
wire \us13/_0572_ ;
wire \us13/_0573_ ;
wire \us13/_0574_ ;
wire \us13/_0575_ ;
wire \us13/_0576_ ;
wire \us13/_0577_ ;
wire \us13/_0578_ ;
wire \us13/_0579_ ;
wire \us13/_0580_ ;
wire \us13/_0581_ ;
wire \us13/_0582_ ;
wire \us13/_0583_ ;
wire \us13/_0584_ ;
wire \us13/_0585_ ;
wire \us13/_0586_ ;
wire \us13/_0587_ ;
wire \us13/_0588_ ;
wire \us13/_0589_ ;
wire \us13/_0590_ ;
wire \us13/_0591_ ;
wire \us13/_0592_ ;
wire \us13/_0593_ ;
wire \us13/_0594_ ;
wire \us13/_0595_ ;
wire \us13/_0596_ ;
wire \us13/_0598_ ;
wire \us13/_0599_ ;
wire \us13/_0600_ ;
wire \us13/_0601_ ;
wire \us13/_0602_ ;
wire \us13/_0603_ ;
wire \us13/_0604_ ;
wire \us13/_0605_ ;
wire \us13/_0606_ ;
wire \us13/_0607_ ;
wire \us13/_0608_ ;
wire \us13/_0609_ ;
wire \us13/_0610_ ;
wire \us13/_0611_ ;
wire \us13/_0612_ ;
wire \us13/_0613_ ;
wire \us13/_0614_ ;
wire \us13/_0615_ ;
wire \us13/_0616_ ;
wire \us13/_0617_ ;
wire \us13/_0618_ ;
wire \us13/_0619_ ;
wire \us13/_0620_ ;
wire \us13/_0621_ ;
wire \us13/_0622_ ;
wire \us13/_0623_ ;
wire \us13/_0624_ ;
wire \us13/_0625_ ;
wire \us13/_0626_ ;
wire \us13/_0627_ ;
wire \us13/_0628_ ;
wire \us13/_0629_ ;
wire \us13/_0630_ ;
wire \us13/_0631_ ;
wire \us13/_0632_ ;
wire \us13/_0633_ ;
wire \us13/_0634_ ;
wire \us13/_0635_ ;
wire \us13/_0636_ ;
wire \us13/_0637_ ;
wire \us13/_0638_ ;
wire \us13/_0639_ ;
wire \us13/_0640_ ;
wire \us13/_0641_ ;
wire \us13/_0642_ ;
wire \us13/_0643_ ;
wire \us13/_0644_ ;
wire \us13/_0645_ ;
wire \us13/_0646_ ;
wire \us13/_0647_ ;
wire \us13/_0648_ ;
wire \us13/_0649_ ;
wire \us13/_0650_ ;
wire \us13/_0652_ ;
wire \us13/_0653_ ;
wire \us13/_0654_ ;
wire \us13/_0655_ ;
wire \us13/_0656_ ;
wire \us13/_0657_ ;
wire \us13/_0658_ ;
wire \us13/_0659_ ;
wire \us13/_0660_ ;
wire \us13/_0661_ ;
wire \us13/_0662_ ;
wire \us13/_0663_ ;
wire \us13/_0664_ ;
wire \us13/_0665_ ;
wire \us13/_0666_ ;
wire \us13/_0667_ ;
wire \us13/_0668_ ;
wire \us13/_0669_ ;
wire \us13/_0670_ ;
wire \us13/_0671_ ;
wire \us13/_0673_ ;
wire \us13/_0674_ ;
wire \us13/_0675_ ;
wire \us13/_0676_ ;
wire \us13/_0677_ ;
wire \us13/_0678_ ;
wire \us13/_0679_ ;
wire \us13/_0680_ ;
wire \us13/_0681_ ;
wire \us13/_0682_ ;
wire \us13/_0683_ ;
wire \us13/_0684_ ;
wire \us13/_0685_ ;
wire \us13/_0686_ ;
wire \us13/_0687_ ;
wire \us13/_0688_ ;
wire \us13/_0689_ ;
wire \us13/_0690_ ;
wire \us13/_0691_ ;
wire \us13/_0692_ ;
wire \us13/_0693_ ;
wire \us13/_0694_ ;
wire \us13/_0695_ ;
wire \us13/_0696_ ;
wire \us13/_0697_ ;
wire \us13/_0698_ ;
wire \us13/_0699_ ;
wire \us13/_0700_ ;
wire \us13/_0701_ ;
wire \us13/_0702_ ;
wire \us13/_0703_ ;
wire \us13/_0704_ ;
wire \us13/_0705_ ;
wire \us13/_0706_ ;
wire \us13/_0707_ ;
wire \us13/_0708_ ;
wire \us13/_0709_ ;
wire \us13/_0710_ ;
wire \us13/_0711_ ;
wire \us13/_0712_ ;
wire \us13/_0713_ ;
wire \us13/_0714_ ;
wire \us13/_0715_ ;
wire \us13/_0716_ ;
wire \us13/_0717_ ;
wire \us13/_0718_ ;
wire \us13/_0719_ ;
wire \us13/_0720_ ;
wire \us13/_0721_ ;
wire \us13/_0722_ ;
wire \us13/_0723_ ;
wire \us13/_0724_ ;
wire \us13/_0725_ ;
wire \us13/_0726_ ;
wire \us13/_0727_ ;
wire \us13/_0728_ ;
wire \us13/_0729_ ;
wire \us13/_0730_ ;
wire \us13/_0731_ ;
wire \us13/_0732_ ;
wire \us13/_0733_ ;
wire \us13/_0734_ ;
wire \us13/_0735_ ;
wire \us13/_0736_ ;
wire \us13/_0738_ ;
wire \us13/_0739_ ;
wire \us13/_0740_ ;
wire \us13/_0741_ ;
wire \us13/_0742_ ;
wire \us13/_0744_ ;
wire \us13/_0745_ ;
wire \us13/_0746_ ;
wire \us13/_0747_ ;
wire \us13/_0748_ ;
wire \us13/_0749_ ;
wire \us13/_0750_ ;
wire \us13/_0752_ ;
wire \us20/_0008_ ;
wire \us20/_0009_ ;
wire \us20/_0010_ ;
wire \us20/_0011_ ;
wire \us20/_0012_ ;
wire \us20/_0013_ ;
wire \us20/_0014_ ;
wire \us20/_0015_ ;
wire \us20/_0016_ ;
wire \us20/_0017_ ;
wire \us20/_0019_ ;
wire \us20/_0020_ ;
wire \us20/_0022_ ;
wire \us20/_0024_ ;
wire \us20/_0025_ ;
wire \us20/_0026_ ;
wire \us20/_0027_ ;
wire \us20/_0030_ ;
wire \us20/_0032_ ;
wire \us20/_0033_ ;
wire \us20/_0034_ ;
wire \us20/_0035_ ;
wire \us20/_0037_ ;
wire \us20/_0038_ ;
wire \us20/_0039_ ;
wire \us20/_0040_ ;
wire \us20/_0041_ ;
wire \us20/_0042_ ;
wire \us20/_0043_ ;
wire \us20/_0045_ ;
wire \us20/_0046_ ;
wire \us20/_0047_ ;
wire \us20/_0049_ ;
wire \us20/_0050_ ;
wire \us20/_0051_ ;
wire \us20/_0052_ ;
wire \us20/_0053_ ;
wire \us20/_0054_ ;
wire \us20/_0057_ ;
wire \us20/_0058_ ;
wire \us20/_0060_ ;
wire \us20/_0061_ ;
wire \us20/_0062_ ;
wire \us20/_0064_ ;
wire \us20/_0065_ ;
wire \us20/_0066_ ;
wire \us20/_0067_ ;
wire \us20/_0069_ ;
wire \us20/_0070_ ;
wire \us20/_0072_ ;
wire \us20/_0073_ ;
wire \us20/_0074_ ;
wire \us20/_0075_ ;
wire \us20/_0076_ ;
wire \us20/_0077_ ;
wire \us20/_0078_ ;
wire \us20/_0079_ ;
wire \us20/_0081_ ;
wire \us20/_0082_ ;
wire \us20/_0084_ ;
wire \us20/_0085_ ;
wire \us20/_0086_ ;
wire \us20/_0087_ ;
wire \us20/_0088_ ;
wire \us20/_0089_ ;
wire \us20/_0090_ ;
wire \us20/_0091_ ;
wire \us20/_0092_ ;
wire \us20/_0093_ ;
wire \us20/_0094_ ;
wire \us20/_0095_ ;
wire \us20/_0096_ ;
wire \us20/_0097_ ;
wire \us20/_0098_ ;
wire \us20/_0099_ ;
wire \us20/_0100_ ;
wire \us20/_0101_ ;
wire \us20/_0102_ ;
wire \us20/_0103_ ;
wire \us20/_0104_ ;
wire \us20/_0105_ ;
wire \us20/_0106_ ;
wire \us20/_0107_ ;
wire \us20/_0108_ ;
wire \us20/_0109_ ;
wire \us20/_0110_ ;
wire \us20/_0111_ ;
wire \us20/_0113_ ;
wire \us20/_0114_ ;
wire \us20/_0115_ ;
wire \us20/_0116_ ;
wire \us20/_0117_ ;
wire \us20/_0118_ ;
wire \us20/_0119_ ;
wire \us20/_0120_ ;
wire \us20/_0121_ ;
wire \us20/_0122_ ;
wire \us20/_0123_ ;
wire \us20/_0124_ ;
wire \us20/_0126_ ;
wire \us20/_0127_ ;
wire \us20/_0128_ ;
wire \us20/_0129_ ;
wire \us20/_0130_ ;
wire \us20/_0132_ ;
wire \us20/_0133_ ;
wire \us20/_0134_ ;
wire \us20/_0135_ ;
wire \us20/_0136_ ;
wire \us20/_0137_ ;
wire \us20/_0139_ ;
wire \us20/_0140_ ;
wire \us20/_0141_ ;
wire \us20/_0142_ ;
wire \us20/_0144_ ;
wire \us20/_0145_ ;
wire \us20/_0146_ ;
wire \us20/_0147_ ;
wire \us20/_0148_ ;
wire \us20/_0149_ ;
wire \us20/_0150_ ;
wire \us20/_0151_ ;
wire \us20/_0153_ ;
wire \us20/_0154_ ;
wire \us20/_0155_ ;
wire \us20/_0156_ ;
wire \us20/_0157_ ;
wire \us20/_0158_ ;
wire \us20/_0159_ ;
wire \us20/_0161_ ;
wire \us20/_0162_ ;
wire \us20/_0163_ ;
wire \us20/_0164_ ;
wire \us20/_0165_ ;
wire \us20/_0166_ ;
wire \us20/_0167_ ;
wire \us20/_0168_ ;
wire \us20/_0169_ ;
wire \us20/_0170_ ;
wire \us20/_0171_ ;
wire \us20/_0172_ ;
wire \us20/_0174_ ;
wire \us20/_0175_ ;
wire \us20/_0176_ ;
wire \us20/_0177_ ;
wire \us20/_0178_ ;
wire \us20/_0179_ ;
wire \us20/_0180_ ;
wire \us20/_0181_ ;
wire \us20/_0182_ ;
wire \us20/_0183_ ;
wire \us20/_0184_ ;
wire \us20/_0185_ ;
wire \us20/_0186_ ;
wire \us20/_0187_ ;
wire \us20/_0188_ ;
wire \us20/_0189_ ;
wire \us20/_0190_ ;
wire \us20/_0191_ ;
wire \us20/_0192_ ;
wire \us20/_0193_ ;
wire \us20/_0194_ ;
wire \us20/_0195_ ;
wire \us20/_0196_ ;
wire \us20/_0197_ ;
wire \us20/_0198_ ;
wire \us20/_0199_ ;
wire \us20/_0200_ ;
wire \us20/_0201_ ;
wire \us20/_0202_ ;
wire \us20/_0203_ ;
wire \us20/_0204_ ;
wire \us20/_0205_ ;
wire \us20/_0206_ ;
wire \us20/_0207_ ;
wire \us20/_0208_ ;
wire \us20/_0209_ ;
wire \us20/_0210_ ;
wire \us20/_0211_ ;
wire \us20/_0212_ ;
wire \us20/_0213_ ;
wire \us20/_0214_ ;
wire \us20/_0215_ ;
wire \us20/_0216_ ;
wire \us20/_0217_ ;
wire \us20/_0218_ ;
wire \us20/_0219_ ;
wire \us20/_0220_ ;
wire \us20/_0221_ ;
wire \us20/_0222_ ;
wire \us20/_0223_ ;
wire \us20/_0224_ ;
wire \us20/_0225_ ;
wire \us20/_0226_ ;
wire \us20/_0227_ ;
wire \us20/_0228_ ;
wire \us20/_0229_ ;
wire \us20/_0230_ ;
wire \us20/_0231_ ;
wire \us20/_0232_ ;
wire \us20/_0233_ ;
wire \us20/_0234_ ;
wire \us20/_0235_ ;
wire \us20/_0236_ ;
wire \us20/_0237_ ;
wire \us20/_0238_ ;
wire \us20/_0239_ ;
wire \us20/_0240_ ;
wire \us20/_0241_ ;
wire \us20/_0242_ ;
wire \us20/_0243_ ;
wire \us20/_0244_ ;
wire \us20/_0245_ ;
wire \us20/_0246_ ;
wire \us20/_0247_ ;
wire \us20/_0248_ ;
wire \us20/_0249_ ;
wire \us20/_0250_ ;
wire \us20/_0251_ ;
wire \us20/_0252_ ;
wire \us20/_0253_ ;
wire \us20/_0254_ ;
wire \us20/_0255_ ;
wire \us20/_0256_ ;
wire \us20/_0257_ ;
wire \us20/_0258_ ;
wire \us20/_0259_ ;
wire \us20/_0260_ ;
wire \us20/_0261_ ;
wire \us20/_0263_ ;
wire \us20/_0264_ ;
wire \us20/_0265_ ;
wire \us20/_0266_ ;
wire \us20/_0267_ ;
wire \us20/_0268_ ;
wire \us20/_0269_ ;
wire \us20/_0270_ ;
wire \us20/_0271_ ;
wire \us20/_0272_ ;
wire \us20/_0273_ ;
wire \us20/_0274_ ;
wire \us20/_0275_ ;
wire \us20/_0276_ ;
wire \us20/_0277_ ;
wire \us20/_0278_ ;
wire \us20/_0279_ ;
wire \us20/_0281_ ;
wire \us20/_0283_ ;
wire \us20/_0284_ ;
wire \us20/_0285_ ;
wire \us20/_0286_ ;
wire \us20/_0287_ ;
wire \us20/_0288_ ;
wire \us20/_0289_ ;
wire \us20/_0290_ ;
wire \us20/_0291_ ;
wire \us20/_0292_ ;
wire \us20/_0293_ ;
wire \us20/_0294_ ;
wire \us20/_0295_ ;
wire \us20/_0296_ ;
wire \us20/_0297_ ;
wire \us20/_0298_ ;
wire \us20/_0299_ ;
wire \us20/_0300_ ;
wire \us20/_0301_ ;
wire \us20/_0302_ ;
wire \us20/_0303_ ;
wire \us20/_0304_ ;
wire \us20/_0305_ ;
wire \us20/_0306_ ;
wire \us20/_0307_ ;
wire \us20/_0308_ ;
wire \us20/_0309_ ;
wire \us20/_0310_ ;
wire \us20/_0311_ ;
wire \us20/_0312_ ;
wire \us20/_0313_ ;
wire \us20/_0314_ ;
wire \us20/_0315_ ;
wire \us20/_0316_ ;
wire \us20/_0317_ ;
wire \us20/_0318_ ;
wire \us20/_0319_ ;
wire \us20/_0320_ ;
wire \us20/_0321_ ;
wire \us20/_0322_ ;
wire \us20/_0323_ ;
wire \us20/_0324_ ;
wire \us20/_0325_ ;
wire \us20/_0326_ ;
wire \us20/_0327_ ;
wire \us20/_0328_ ;
wire \us20/_0329_ ;
wire \us20/_0330_ ;
wire \us20/_0331_ ;
wire \us20/_0332_ ;
wire \us20/_0333_ ;
wire \us20/_0334_ ;
wire \us20/_0335_ ;
wire \us20/_0337_ ;
wire \us20/_0338_ ;
wire \us20/_0339_ ;
wire \us20/_0340_ ;
wire \us20/_0341_ ;
wire \us20/_0342_ ;
wire \us20/_0343_ ;
wire \us20/_0344_ ;
wire \us20/_0345_ ;
wire \us20/_0347_ ;
wire \us20/_0348_ ;
wire \us20/_0349_ ;
wire \us20/_0350_ ;
wire \us20/_0351_ ;
wire \us20/_0352_ ;
wire \us20/_0353_ ;
wire \us20/_0354_ ;
wire \us20/_0355_ ;
wire \us20/_0356_ ;
wire \us20/_0357_ ;
wire \us20/_0358_ ;
wire \us20/_0359_ ;
wire \us20/_0360_ ;
wire \us20/_0361_ ;
wire \us20/_0362_ ;
wire \us20/_0363_ ;
wire \us20/_0365_ ;
wire \us20/_0366_ ;
wire \us20/_0367_ ;
wire \us20/_0368_ ;
wire \us20/_0370_ ;
wire \us20/_0371_ ;
wire \us20/_0372_ ;
wire \us20/_0373_ ;
wire \us20/_0374_ ;
wire \us20/_0375_ ;
wire \us20/_0376_ ;
wire \us20/_0377_ ;
wire \us20/_0378_ ;
wire \us20/_0379_ ;
wire \us20/_0380_ ;
wire \us20/_0381_ ;
wire \us20/_0382_ ;
wire \us20/_0383_ ;
wire \us20/_0384_ ;
wire \us20/_0385_ ;
wire \us20/_0386_ ;
wire \us20/_0387_ ;
wire \us20/_0388_ ;
wire \us20/_0389_ ;
wire \us20/_0390_ ;
wire \us20/_0391_ ;
wire \us20/_0392_ ;
wire \us20/_0393_ ;
wire \us20/_0394_ ;
wire \us20/_0395_ ;
wire \us20/_0396_ ;
wire \us20/_0397_ ;
wire \us20/_0398_ ;
wire \us20/_0399_ ;
wire \us20/_0400_ ;
wire \us20/_0401_ ;
wire \us20/_0402_ ;
wire \us20/_0403_ ;
wire \us20/_0404_ ;
wire \us20/_0405_ ;
wire \us20/_0406_ ;
wire \us20/_0407_ ;
wire \us20/_0408_ ;
wire \us20/_0409_ ;
wire \us20/_0410_ ;
wire \us20/_0411_ ;
wire \us20/_0412_ ;
wire \us20/_0413_ ;
wire \us20/_0414_ ;
wire \us20/_0415_ ;
wire \us20/_0416_ ;
wire \us20/_0417_ ;
wire \us20/_0418_ ;
wire \us20/_0419_ ;
wire \us20/_0420_ ;
wire \us20/_0421_ ;
wire \us20/_0422_ ;
wire \us20/_0423_ ;
wire \us20/_0424_ ;
wire \us20/_0425_ ;
wire \us20/_0426_ ;
wire \us20/_0427_ ;
wire \us20/_0428_ ;
wire \us20/_0429_ ;
wire \us20/_0430_ ;
wire \us20/_0431_ ;
wire \us20/_0432_ ;
wire \us20/_0433_ ;
wire \us20/_0434_ ;
wire \us20/_0435_ ;
wire \us20/_0436_ ;
wire \us20/_0437_ ;
wire \us20/_0438_ ;
wire \us20/_0439_ ;
wire \us20/_0440_ ;
wire \us20/_0441_ ;
wire \us20/_0442_ ;
wire \us20/_0443_ ;
wire \us20/_0444_ ;
wire \us20/_0446_ ;
wire \us20/_0447_ ;
wire \us20/_0448_ ;
wire \us20/_0449_ ;
wire \us20/_0450_ ;
wire \us20/_0451_ ;
wire \us20/_0452_ ;
wire \us20/_0453_ ;
wire \us20/_0454_ ;
wire \us20/_0455_ ;
wire \us20/_0457_ ;
wire \us20/_0458_ ;
wire \us20/_0459_ ;
wire \us20/_0460_ ;
wire \us20/_0461_ ;
wire \us20/_0462_ ;
wire \us20/_0463_ ;
wire \us20/_0464_ ;
wire \us20/_0465_ ;
wire \us20/_0466_ ;
wire \us20/_0467_ ;
wire \us20/_0468_ ;
wire \us20/_0469_ ;
wire \us20/_0470_ ;
wire \us20/_0471_ ;
wire \us20/_0472_ ;
wire \us20/_0473_ ;
wire \us20/_0474_ ;
wire \us20/_0475_ ;
wire \us20/_0476_ ;
wire \us20/_0477_ ;
wire \us20/_0478_ ;
wire \us20/_0479_ ;
wire \us20/_0480_ ;
wire \us20/_0481_ ;
wire \us20/_0482_ ;
wire \us20/_0483_ ;
wire \us20/_0484_ ;
wire \us20/_0485_ ;
wire \us20/_0486_ ;
wire \us20/_0487_ ;
wire \us20/_0488_ ;
wire \us20/_0490_ ;
wire \us20/_0491_ ;
wire \us20/_0492_ ;
wire \us20/_0493_ ;
wire \us20/_0494_ ;
wire \us20/_0495_ ;
wire \us20/_0496_ ;
wire \us20/_0497_ ;
wire \us20/_0498_ ;
wire \us20/_0500_ ;
wire \us20/_0501_ ;
wire \us20/_0502_ ;
wire \us20/_0503_ ;
wire \us20/_0504_ ;
wire \us20/_0505_ ;
wire \us20/_0506_ ;
wire \us20/_0507_ ;
wire \us20/_0508_ ;
wire \us20/_0509_ ;
wire \us20/_0510_ ;
wire \us20/_0511_ ;
wire \us20/_0512_ ;
wire \us20/_0513_ ;
wire \us20/_0514_ ;
wire \us20/_0515_ ;
wire \us20/_0516_ ;
wire \us20/_0517_ ;
wire \us20/_0518_ ;
wire \us20/_0519_ ;
wire \us20/_0520_ ;
wire \us20/_0521_ ;
wire \us20/_0522_ ;
wire \us20/_0523_ ;
wire \us20/_0524_ ;
wire \us20/_0525_ ;
wire \us20/_0526_ ;
wire \us20/_0527_ ;
wire \us20/_0528_ ;
wire \us20/_0529_ ;
wire \us20/_0530_ ;
wire \us20/_0531_ ;
wire \us20/_0532_ ;
wire \us20/_0533_ ;
wire \us20/_0534_ ;
wire \us20/_0535_ ;
wire \us20/_0536_ ;
wire \us20/_0537_ ;
wire \us20/_0538_ ;
wire \us20/_0539_ ;
wire \us20/_0540_ ;
wire \us20/_0541_ ;
wire \us20/_0542_ ;
wire \us20/_0543_ ;
wire \us20/_0544_ ;
wire \us20/_0545_ ;
wire \us20/_0546_ ;
wire \us20/_0547_ ;
wire \us20/_0548_ ;
wire \us20/_0549_ ;
wire \us20/_0550_ ;
wire \us20/_0551_ ;
wire \us20/_0552_ ;
wire \us20/_0553_ ;
wire \us20/_0554_ ;
wire \us20/_0555_ ;
wire \us20/_0556_ ;
wire \us20/_0557_ ;
wire \us20/_0558_ ;
wire \us20/_0559_ ;
wire \us20/_0560_ ;
wire \us20/_0561_ ;
wire \us20/_0562_ ;
wire \us20/_0563_ ;
wire \us20/_0565_ ;
wire \us20/_0566_ ;
wire \us20/_0567_ ;
wire \us20/_0568_ ;
wire \us20/_0569_ ;
wire \us20/_0570_ ;
wire \us20/_0571_ ;
wire \us20/_0572_ ;
wire \us20/_0573_ ;
wire \us20/_0574_ ;
wire \us20/_0575_ ;
wire \us20/_0576_ ;
wire \us20/_0577_ ;
wire \us20/_0578_ ;
wire \us20/_0579_ ;
wire \us20/_0580_ ;
wire \us20/_0581_ ;
wire \us20/_0582_ ;
wire \us20/_0583_ ;
wire \us20/_0584_ ;
wire \us20/_0585_ ;
wire \us20/_0586_ ;
wire \us20/_0587_ ;
wire \us20/_0588_ ;
wire \us20/_0589_ ;
wire \us20/_0590_ ;
wire \us20/_0591_ ;
wire \us20/_0592_ ;
wire \us20/_0593_ ;
wire \us20/_0594_ ;
wire \us20/_0595_ ;
wire \us20/_0596_ ;
wire \us20/_0598_ ;
wire \us20/_0599_ ;
wire \us20/_0600_ ;
wire \us20/_0601_ ;
wire \us20/_0602_ ;
wire \us20/_0603_ ;
wire \us20/_0604_ ;
wire \us20/_0605_ ;
wire \us20/_0606_ ;
wire \us20/_0607_ ;
wire \us20/_0608_ ;
wire \us20/_0609_ ;
wire \us20/_0610_ ;
wire \us20/_0611_ ;
wire \us20/_0612_ ;
wire \us20/_0613_ ;
wire \us20/_0614_ ;
wire \us20/_0615_ ;
wire \us20/_0616_ ;
wire \us20/_0617_ ;
wire \us20/_0618_ ;
wire \us20/_0619_ ;
wire \us20/_0620_ ;
wire \us20/_0621_ ;
wire \us20/_0622_ ;
wire \us20/_0623_ ;
wire \us20/_0624_ ;
wire \us20/_0625_ ;
wire \us20/_0626_ ;
wire \us20/_0627_ ;
wire \us20/_0628_ ;
wire \us20/_0629_ ;
wire \us20/_0630_ ;
wire \us20/_0631_ ;
wire \us20/_0632_ ;
wire \us20/_0633_ ;
wire \us20/_0634_ ;
wire \us20/_0635_ ;
wire \us20/_0636_ ;
wire \us20/_0637_ ;
wire \us20/_0638_ ;
wire \us20/_0639_ ;
wire \us20/_0640_ ;
wire \us20/_0641_ ;
wire \us20/_0642_ ;
wire \us20/_0643_ ;
wire \us20/_0644_ ;
wire \us20/_0645_ ;
wire \us20/_0646_ ;
wire \us20/_0647_ ;
wire \us20/_0648_ ;
wire \us20/_0649_ ;
wire \us20/_0650_ ;
wire \us20/_0652_ ;
wire \us20/_0653_ ;
wire \us20/_0654_ ;
wire \us20/_0655_ ;
wire \us20/_0656_ ;
wire \us20/_0657_ ;
wire \us20/_0658_ ;
wire \us20/_0659_ ;
wire \us20/_0660_ ;
wire \us20/_0661_ ;
wire \us20/_0662_ ;
wire \us20/_0663_ ;
wire \us20/_0664_ ;
wire \us20/_0665_ ;
wire \us20/_0666_ ;
wire \us20/_0667_ ;
wire \us20/_0668_ ;
wire \us20/_0669_ ;
wire \us20/_0670_ ;
wire \us20/_0671_ ;
wire \us20/_0672_ ;
wire \us20/_0673_ ;
wire \us20/_0674_ ;
wire \us20/_0675_ ;
wire \us20/_0676_ ;
wire \us20/_0677_ ;
wire \us20/_0678_ ;
wire \us20/_0679_ ;
wire \us20/_0680_ ;
wire \us20/_0681_ ;
wire \us20/_0682_ ;
wire \us20/_0683_ ;
wire \us20/_0684_ ;
wire \us20/_0685_ ;
wire \us20/_0686_ ;
wire \us20/_0687_ ;
wire \us20/_0688_ ;
wire \us20/_0689_ ;
wire \us20/_0690_ ;
wire \us20/_0691_ ;
wire \us20/_0692_ ;
wire \us20/_0693_ ;
wire \us20/_0694_ ;
wire \us20/_0695_ ;
wire \us20/_0696_ ;
wire \us20/_0697_ ;
wire \us20/_0698_ ;
wire \us20/_0699_ ;
wire \us20/_0700_ ;
wire \us20/_0701_ ;
wire \us20/_0702_ ;
wire \us20/_0703_ ;
wire \us20/_0704_ ;
wire \us20/_0705_ ;
wire \us20/_0706_ ;
wire \us20/_0707_ ;
wire \us20/_0708_ ;
wire \us20/_0709_ ;
wire \us20/_0710_ ;
wire \us20/_0711_ ;
wire \us20/_0712_ ;
wire \us20/_0713_ ;
wire \us20/_0714_ ;
wire \us20/_0715_ ;
wire \us20/_0717_ ;
wire \us20/_0718_ ;
wire \us20/_0719_ ;
wire \us20/_0720_ ;
wire \us20/_0721_ ;
wire \us20/_0722_ ;
wire \us20/_0723_ ;
wire \us20/_0724_ ;
wire \us20/_0725_ ;
wire \us20/_0726_ ;
wire \us20/_0727_ ;
wire \us20/_0728_ ;
wire \us20/_0729_ ;
wire \us20/_0730_ ;
wire \us20/_0731_ ;
wire \us20/_0732_ ;
wire \us20/_0733_ ;
wire \us20/_0734_ ;
wire \us20/_0735_ ;
wire \us20/_0736_ ;
wire \us20/_0738_ ;
wire \us20/_0739_ ;
wire \us20/_0740_ ;
wire \us20/_0741_ ;
wire \us20/_0742_ ;
wire \us20/_0744_ ;
wire \us20/_0745_ ;
wire \us20/_0746_ ;
wire \us20/_0748_ ;
wire \us20/_0749_ ;
wire \us20/_0750_ ;
wire \us20/_0752_ ;
wire \us21/_0008_ ;
wire \us21/_0009_ ;
wire \us21/_0010_ ;
wire \us21/_0011_ ;
wire \us21/_0012_ ;
wire \us21/_0013_ ;
wire \us21/_0014_ ;
wire \us21/_0015_ ;
wire \us21/_0016_ ;
wire \us21/_0017_ ;
wire \us21/_0019_ ;
wire \us21/_0020_ ;
wire \us21/_0022_ ;
wire \us21/_0024_ ;
wire \us21/_0025_ ;
wire \us21/_0026_ ;
wire \us21/_0027_ ;
wire \us21/_0030_ ;
wire \us21/_0032_ ;
wire \us21/_0033_ ;
wire \us21/_0034_ ;
wire \us21/_0035_ ;
wire \us21/_0037_ ;
wire \us21/_0038_ ;
wire \us21/_0039_ ;
wire \us21/_0040_ ;
wire \us21/_0041_ ;
wire \us21/_0042_ ;
wire \us21/_0043_ ;
wire \us21/_0045_ ;
wire \us21/_0046_ ;
wire \us21/_0047_ ;
wire \us21/_0049_ ;
wire \us21/_0050_ ;
wire \us21/_0051_ ;
wire \us21/_0052_ ;
wire \us21/_0053_ ;
wire \us21/_0054_ ;
wire \us21/_0056_ ;
wire \us21/_0057_ ;
wire \us21/_0058_ ;
wire \us21/_0060_ ;
wire \us21/_0061_ ;
wire \us21/_0062_ ;
wire \us21/_0064_ ;
wire \us21/_0065_ ;
wire \us21/_0066_ ;
wire \us21/_0067_ ;
wire \us21/_0069_ ;
wire \us21/_0070_ ;
wire \us21/_0072_ ;
wire \us21/_0073_ ;
wire \us21/_0074_ ;
wire \us21/_0075_ ;
wire \us21/_0076_ ;
wire \us21/_0077_ ;
wire \us21/_0078_ ;
wire \us21/_0079_ ;
wire \us21/_0081_ ;
wire \us21/_0082_ ;
wire \us21/_0084_ ;
wire \us21/_0085_ ;
wire \us21/_0086_ ;
wire \us21/_0087_ ;
wire \us21/_0088_ ;
wire \us21/_0089_ ;
wire \us21/_0090_ ;
wire \us21/_0091_ ;
wire \us21/_0092_ ;
wire \us21/_0093_ ;
wire \us21/_0094_ ;
wire \us21/_0095_ ;
wire \us21/_0096_ ;
wire \us21/_0097_ ;
wire \us21/_0098_ ;
wire \us21/_0099_ ;
wire \us21/_0100_ ;
wire \us21/_0101_ ;
wire \us21/_0102_ ;
wire \us21/_0103_ ;
wire \us21/_0104_ ;
wire \us21/_0105_ ;
wire \us21/_0106_ ;
wire \us21/_0108_ ;
wire \us21/_0109_ ;
wire \us21/_0110_ ;
wire \us21/_0111_ ;
wire \us21/_0113_ ;
wire \us21/_0114_ ;
wire \us21/_0115_ ;
wire \us21/_0116_ ;
wire \us21/_0117_ ;
wire \us21/_0118_ ;
wire \us21/_0119_ ;
wire \us21/_0120_ ;
wire \us21/_0121_ ;
wire \us21/_0122_ ;
wire \us21/_0123_ ;
wire \us21/_0124_ ;
wire \us21/_0126_ ;
wire \us21/_0127_ ;
wire \us21/_0128_ ;
wire \us21/_0129_ ;
wire \us21/_0130_ ;
wire \us21/_0132_ ;
wire \us21/_0133_ ;
wire \us21/_0134_ ;
wire \us21/_0135_ ;
wire \us21/_0136_ ;
wire \us21/_0137_ ;
wire \us21/_0139_ ;
wire \us21/_0140_ ;
wire \us21/_0141_ ;
wire \us21/_0142_ ;
wire \us21/_0144_ ;
wire \us21/_0145_ ;
wire \us21/_0146_ ;
wire \us21/_0147_ ;
wire \us21/_0148_ ;
wire \us21/_0149_ ;
wire \us21/_0150_ ;
wire \us21/_0151_ ;
wire \us21/_0153_ ;
wire \us21/_0154_ ;
wire \us21/_0155_ ;
wire \us21/_0156_ ;
wire \us21/_0157_ ;
wire \us21/_0158_ ;
wire \us21/_0159_ ;
wire \us21/_0161_ ;
wire \us21/_0162_ ;
wire \us21/_0163_ ;
wire \us21/_0164_ ;
wire \us21/_0165_ ;
wire \us21/_0166_ ;
wire \us21/_0167_ ;
wire \us21/_0168_ ;
wire \us21/_0169_ ;
wire \us21/_0170_ ;
wire \us21/_0171_ ;
wire \us21/_0172_ ;
wire \us21/_0174_ ;
wire \us21/_0175_ ;
wire \us21/_0176_ ;
wire \us21/_0177_ ;
wire \us21/_0178_ ;
wire \us21/_0179_ ;
wire \us21/_0180_ ;
wire \us21/_0181_ ;
wire \us21/_0182_ ;
wire \us21/_0183_ ;
wire \us21/_0184_ ;
wire \us21/_0185_ ;
wire \us21/_0186_ ;
wire \us21/_0187_ ;
wire \us21/_0188_ ;
wire \us21/_0189_ ;
wire \us21/_0190_ ;
wire \us21/_0191_ ;
wire \us21/_0192_ ;
wire \us21/_0193_ ;
wire \us21/_0194_ ;
wire \us21/_0195_ ;
wire \us21/_0196_ ;
wire \us21/_0197_ ;
wire \us21/_0198_ ;
wire \us21/_0199_ ;
wire \us21/_0200_ ;
wire \us21/_0201_ ;
wire \us21/_0202_ ;
wire \us21/_0203_ ;
wire \us21/_0204_ ;
wire \us21/_0205_ ;
wire \us21/_0206_ ;
wire \us21/_0207_ ;
wire \us21/_0208_ ;
wire \us21/_0209_ ;
wire \us21/_0210_ ;
wire \us21/_0211_ ;
wire \us21/_0212_ ;
wire \us21/_0213_ ;
wire \us21/_0214_ ;
wire \us21/_0215_ ;
wire \us21/_0217_ ;
wire \us21/_0218_ ;
wire \us21/_0219_ ;
wire \us21/_0220_ ;
wire \us21/_0221_ ;
wire \us21/_0222_ ;
wire \us21/_0223_ ;
wire \us21/_0224_ ;
wire \us21/_0225_ ;
wire \us21/_0226_ ;
wire \us21/_0227_ ;
wire \us21/_0228_ ;
wire \us21/_0229_ ;
wire \us21/_0230_ ;
wire \us21/_0231_ ;
wire \us21/_0232_ ;
wire \us21/_0233_ ;
wire \us21/_0234_ ;
wire \us21/_0235_ ;
wire \us21/_0236_ ;
wire \us21/_0237_ ;
wire \us21/_0238_ ;
wire \us21/_0239_ ;
wire \us21/_0240_ ;
wire \us21/_0241_ ;
wire \us21/_0242_ ;
wire \us21/_0243_ ;
wire \us21/_0244_ ;
wire \us21/_0245_ ;
wire \us21/_0246_ ;
wire \us21/_0247_ ;
wire \us21/_0248_ ;
wire \us21/_0249_ ;
wire \us21/_0250_ ;
wire \us21/_0251_ ;
wire \us21/_0252_ ;
wire \us21/_0253_ ;
wire \us21/_0254_ ;
wire \us21/_0255_ ;
wire \us21/_0256_ ;
wire \us21/_0257_ ;
wire \us21/_0258_ ;
wire \us21/_0259_ ;
wire \us21/_0260_ ;
wire \us21/_0261_ ;
wire \us21/_0263_ ;
wire \us21/_0264_ ;
wire \us21/_0265_ ;
wire \us21/_0266_ ;
wire \us21/_0267_ ;
wire \us21/_0268_ ;
wire \us21/_0269_ ;
wire \us21/_0270_ ;
wire \us21/_0271_ ;
wire \us21/_0272_ ;
wire \us21/_0273_ ;
wire \us21/_0274_ ;
wire \us21/_0275_ ;
wire \us21/_0276_ ;
wire \us21/_0277_ ;
wire \us21/_0278_ ;
wire \us21/_0279_ ;
wire \us21/_0281_ ;
wire \us21/_0283_ ;
wire \us21/_0284_ ;
wire \us21/_0285_ ;
wire \us21/_0286_ ;
wire \us21/_0287_ ;
wire \us21/_0288_ ;
wire \us21/_0289_ ;
wire \us21/_0290_ ;
wire \us21/_0291_ ;
wire \us21/_0293_ ;
wire \us21/_0294_ ;
wire \us21/_0295_ ;
wire \us21/_0296_ ;
wire \us21/_0297_ ;
wire \us21/_0298_ ;
wire \us21/_0299_ ;
wire \us21/_0300_ ;
wire \us21/_0301_ ;
wire \us21/_0302_ ;
wire \us21/_0303_ ;
wire \us21/_0304_ ;
wire \us21/_0305_ ;
wire \us21/_0306_ ;
wire \us21/_0307_ ;
wire \us21/_0308_ ;
wire \us21/_0309_ ;
wire \us21/_0310_ ;
wire \us21/_0311_ ;
wire \us21/_0312_ ;
wire \us21/_0313_ ;
wire \us21/_0314_ ;
wire \us21/_0315_ ;
wire \us21/_0316_ ;
wire \us21/_0317_ ;
wire \us21/_0318_ ;
wire \us21/_0319_ ;
wire \us21/_0320_ ;
wire \us21/_0321_ ;
wire \us21/_0322_ ;
wire \us21/_0323_ ;
wire \us21/_0324_ ;
wire \us21/_0325_ ;
wire \us21/_0326_ ;
wire \us21/_0327_ ;
wire \us21/_0328_ ;
wire \us21/_0329_ ;
wire \us21/_0330_ ;
wire \us21/_0331_ ;
wire \us21/_0332_ ;
wire \us21/_0333_ ;
wire \us21/_0334_ ;
wire \us21/_0335_ ;
wire \us21/_0337_ ;
wire \us21/_0338_ ;
wire \us21/_0339_ ;
wire \us21/_0340_ ;
wire \us21/_0341_ ;
wire \us21/_0342_ ;
wire \us21/_0343_ ;
wire \us21/_0344_ ;
wire \us21/_0345_ ;
wire \us21/_0347_ ;
wire \us21/_0348_ ;
wire \us21/_0349_ ;
wire \us21/_0350_ ;
wire \us21/_0351_ ;
wire \us21/_0352_ ;
wire \us21/_0353_ ;
wire \us21/_0354_ ;
wire \us21/_0355_ ;
wire \us21/_0356_ ;
wire \us21/_0357_ ;
wire \us21/_0358_ ;
wire \us21/_0359_ ;
wire \us21/_0360_ ;
wire \us21/_0361_ ;
wire \us21/_0362_ ;
wire \us21/_0363_ ;
wire \us21/_0365_ ;
wire \us21/_0366_ ;
wire \us21/_0367_ ;
wire \us21/_0368_ ;
wire \us21/_0370_ ;
wire \us21/_0371_ ;
wire \us21/_0372_ ;
wire \us21/_0373_ ;
wire \us21/_0374_ ;
wire \us21/_0375_ ;
wire \us21/_0376_ ;
wire \us21/_0377_ ;
wire \us21/_0378_ ;
wire \us21/_0379_ ;
wire \us21/_0380_ ;
wire \us21/_0381_ ;
wire \us21/_0382_ ;
wire \us21/_0383_ ;
wire \us21/_0384_ ;
wire \us21/_0385_ ;
wire \us21/_0386_ ;
wire \us21/_0387_ ;
wire \us21/_0388_ ;
wire \us21/_0389_ ;
wire \us21/_0390_ ;
wire \us21/_0391_ ;
wire \us21/_0392_ ;
wire \us21/_0393_ ;
wire \us21/_0394_ ;
wire \us21/_0395_ ;
wire \us21/_0396_ ;
wire \us21/_0397_ ;
wire \us21/_0398_ ;
wire \us21/_0399_ ;
wire \us21/_0400_ ;
wire \us21/_0401_ ;
wire \us21/_0402_ ;
wire \us21/_0403_ ;
wire \us21/_0404_ ;
wire \us21/_0405_ ;
wire \us21/_0406_ ;
wire \us21/_0407_ ;
wire \us21/_0408_ ;
wire \us21/_0409_ ;
wire \us21/_0410_ ;
wire \us21/_0411_ ;
wire \us21/_0412_ ;
wire \us21/_0413_ ;
wire \us21/_0414_ ;
wire \us21/_0415_ ;
wire \us21/_0416_ ;
wire \us21/_0417_ ;
wire \us21/_0418_ ;
wire \us21/_0419_ ;
wire \us21/_0420_ ;
wire \us21/_0421_ ;
wire \us21/_0422_ ;
wire \us21/_0424_ ;
wire \us21/_0425_ ;
wire \us21/_0426_ ;
wire \us21/_0427_ ;
wire \us21/_0428_ ;
wire \us21/_0429_ ;
wire \us21/_0430_ ;
wire \us21/_0431_ ;
wire \us21/_0432_ ;
wire \us21/_0433_ ;
wire \us21/_0434_ ;
wire \us21/_0435_ ;
wire \us21/_0436_ ;
wire \us21/_0437_ ;
wire \us21/_0438_ ;
wire \us21/_0439_ ;
wire \us21/_0440_ ;
wire \us21/_0441_ ;
wire \us21/_0442_ ;
wire \us21/_0443_ ;
wire \us21/_0444_ ;
wire \us21/_0446_ ;
wire \us21/_0447_ ;
wire \us21/_0448_ ;
wire \us21/_0449_ ;
wire \us21/_0450_ ;
wire \us21/_0451_ ;
wire \us21/_0452_ ;
wire \us21/_0453_ ;
wire \us21/_0454_ ;
wire \us21/_0455_ ;
wire \us21/_0457_ ;
wire \us21/_0458_ ;
wire \us21/_0459_ ;
wire \us21/_0460_ ;
wire \us21/_0461_ ;
wire \us21/_0462_ ;
wire \us21/_0463_ ;
wire \us21/_0464_ ;
wire \us21/_0465_ ;
wire \us21/_0466_ ;
wire \us21/_0467_ ;
wire \us21/_0468_ ;
wire \us21/_0469_ ;
wire \us21/_0470_ ;
wire \us21/_0471_ ;
wire \us21/_0472_ ;
wire \us21/_0473_ ;
wire \us21/_0474_ ;
wire \us21/_0475_ ;
wire \us21/_0476_ ;
wire \us21/_0477_ ;
wire \us21/_0478_ ;
wire \us21/_0479_ ;
wire \us21/_0480_ ;
wire \us21/_0481_ ;
wire \us21/_0482_ ;
wire \us21/_0483_ ;
wire \us21/_0484_ ;
wire \us21/_0485_ ;
wire \us21/_0486_ ;
wire \us21/_0487_ ;
wire \us21/_0488_ ;
wire \us21/_0490_ ;
wire \us21/_0491_ ;
wire \us21/_0492_ ;
wire \us21/_0493_ ;
wire \us21/_0494_ ;
wire \us21/_0495_ ;
wire \us21/_0496_ ;
wire \us21/_0497_ ;
wire \us21/_0498_ ;
wire \us21/_0500_ ;
wire \us21/_0501_ ;
wire \us21/_0502_ ;
wire \us21/_0503_ ;
wire \us21/_0504_ ;
wire \us21/_0505_ ;
wire \us21/_0506_ ;
wire \us21/_0507_ ;
wire \us21/_0508_ ;
wire \us21/_0509_ ;
wire \us21/_0510_ ;
wire \us21/_0511_ ;
wire \us21/_0512_ ;
wire \us21/_0513_ ;
wire \us21/_0514_ ;
wire \us21/_0515_ ;
wire \us21/_0516_ ;
wire \us21/_0517_ ;
wire \us21/_0518_ ;
wire \us21/_0519_ ;
wire \us21/_0520_ ;
wire \us21/_0521_ ;
wire \us21/_0522_ ;
wire \us21/_0523_ ;
wire \us21/_0524_ ;
wire \us21/_0525_ ;
wire \us21/_0526_ ;
wire \us21/_0527_ ;
wire \us21/_0528_ ;
wire \us21/_0529_ ;
wire \us21/_0530_ ;
wire \us21/_0531_ ;
wire \us21/_0532_ ;
wire \us21/_0533_ ;
wire \us21/_0534_ ;
wire \us21/_0535_ ;
wire \us21/_0536_ ;
wire \us21/_0537_ ;
wire \us21/_0538_ ;
wire \us21/_0539_ ;
wire \us21/_0540_ ;
wire \us21/_0541_ ;
wire \us21/_0542_ ;
wire \us21/_0544_ ;
wire \us21/_0545_ ;
wire \us21/_0546_ ;
wire \us21/_0547_ ;
wire \us21/_0548_ ;
wire \us21/_0549_ ;
wire \us21/_0550_ ;
wire \us21/_0551_ ;
wire \us21/_0552_ ;
wire \us21/_0553_ ;
wire \us21/_0554_ ;
wire \us21/_0555_ ;
wire \us21/_0556_ ;
wire \us21/_0557_ ;
wire \us21/_0558_ ;
wire \us21/_0559_ ;
wire \us21/_0560_ ;
wire \us21/_0561_ ;
wire \us21/_0562_ ;
wire \us21/_0563_ ;
wire \us21/_0565_ ;
wire \us21/_0566_ ;
wire \us21/_0567_ ;
wire \us21/_0568_ ;
wire \us21/_0569_ ;
wire \us21/_0570_ ;
wire \us21/_0571_ ;
wire \us21/_0572_ ;
wire \us21/_0573_ ;
wire \us21/_0574_ ;
wire \us21/_0575_ ;
wire \us21/_0576_ ;
wire \us21/_0577_ ;
wire \us21/_0578_ ;
wire \us21/_0579_ ;
wire \us21/_0580_ ;
wire \us21/_0581_ ;
wire \us21/_0582_ ;
wire \us21/_0583_ ;
wire \us21/_0584_ ;
wire \us21/_0585_ ;
wire \us21/_0586_ ;
wire \us21/_0587_ ;
wire \us21/_0588_ ;
wire \us21/_0589_ ;
wire \us21/_0590_ ;
wire \us21/_0591_ ;
wire \us21/_0592_ ;
wire \us21/_0593_ ;
wire \us21/_0594_ ;
wire \us21/_0595_ ;
wire \us21/_0596_ ;
wire \us21/_0598_ ;
wire \us21/_0599_ ;
wire \us21/_0600_ ;
wire \us21/_0601_ ;
wire \us21/_0602_ ;
wire \us21/_0603_ ;
wire \us21/_0604_ ;
wire \us21/_0605_ ;
wire \us21/_0606_ ;
wire \us21/_0607_ ;
wire \us21/_0608_ ;
wire \us21/_0609_ ;
wire \us21/_0610_ ;
wire \us21/_0611_ ;
wire \us21/_0612_ ;
wire \us21/_0613_ ;
wire \us21/_0614_ ;
wire \us21/_0615_ ;
wire \us21/_0616_ ;
wire \us21/_0617_ ;
wire \us21/_0618_ ;
wire \us21/_0619_ ;
wire \us21/_0620_ ;
wire \us21/_0621_ ;
wire \us21/_0622_ ;
wire \us21/_0623_ ;
wire \us21/_0624_ ;
wire \us21/_0625_ ;
wire \us21/_0626_ ;
wire \us21/_0627_ ;
wire \us21/_0628_ ;
wire \us21/_0629_ ;
wire \us21/_0630_ ;
wire \us21/_0631_ ;
wire \us21/_0632_ ;
wire \us21/_0633_ ;
wire \us21/_0634_ ;
wire \us21/_0635_ ;
wire \us21/_0636_ ;
wire \us21/_0637_ ;
wire \us21/_0638_ ;
wire \us21/_0639_ ;
wire \us21/_0640_ ;
wire \us21/_0641_ ;
wire \us21/_0642_ ;
wire \us21/_0643_ ;
wire \us21/_0644_ ;
wire \us21/_0645_ ;
wire \us21/_0646_ ;
wire \us21/_0647_ ;
wire \us21/_0648_ ;
wire \us21/_0649_ ;
wire \us21/_0650_ ;
wire \us21/_0652_ ;
wire \us21/_0653_ ;
wire \us21/_0654_ ;
wire \us21/_0655_ ;
wire \us21/_0656_ ;
wire \us21/_0657_ ;
wire \us21/_0658_ ;
wire \us21/_0659_ ;
wire \us21/_0660_ ;
wire \us21/_0661_ ;
wire \us21/_0662_ ;
wire \us21/_0663_ ;
wire \us21/_0664_ ;
wire \us21/_0665_ ;
wire \us21/_0666_ ;
wire \us21/_0667_ ;
wire \us21/_0668_ ;
wire \us21/_0669_ ;
wire \us21/_0670_ ;
wire \us21/_0671_ ;
wire \us21/_0673_ ;
wire \us21/_0674_ ;
wire \us21/_0675_ ;
wire \us21/_0676_ ;
wire \us21/_0677_ ;
wire \us21/_0678_ ;
wire \us21/_0679_ ;
wire \us21/_0680_ ;
wire \us21/_0681_ ;
wire \us21/_0682_ ;
wire \us21/_0683_ ;
wire \us21/_0684_ ;
wire \us21/_0685_ ;
wire \us21/_0686_ ;
wire \us21/_0687_ ;
wire \us21/_0688_ ;
wire \us21/_0689_ ;
wire \us21/_0690_ ;
wire \us21/_0691_ ;
wire \us21/_0692_ ;
wire \us21/_0693_ ;
wire \us21/_0694_ ;
wire \us21/_0695_ ;
wire \us21/_0696_ ;
wire \us21/_0697_ ;
wire \us21/_0698_ ;
wire \us21/_0699_ ;
wire \us21/_0700_ ;
wire \us21/_0701_ ;
wire \us21/_0702_ ;
wire \us21/_0703_ ;
wire \us21/_0704_ ;
wire \us21/_0705_ ;
wire \us21/_0706_ ;
wire \us21/_0707_ ;
wire \us21/_0708_ ;
wire \us21/_0709_ ;
wire \us21/_0710_ ;
wire \us21/_0711_ ;
wire \us21/_0712_ ;
wire \us21/_0713_ ;
wire \us21/_0714_ ;
wire \us21/_0715_ ;
wire \us21/_0717_ ;
wire \us21/_0718_ ;
wire \us21/_0719_ ;
wire \us21/_0720_ ;
wire \us21/_0721_ ;
wire \us21/_0722_ ;
wire \us21/_0723_ ;
wire \us21/_0724_ ;
wire \us21/_0725_ ;
wire \us21/_0726_ ;
wire \us21/_0727_ ;
wire \us21/_0728_ ;
wire \us21/_0729_ ;
wire \us21/_0730_ ;
wire \us21/_0731_ ;
wire \us21/_0733_ ;
wire \us21/_0734_ ;
wire \us21/_0735_ ;
wire \us21/_0736_ ;
wire \us21/_0738_ ;
wire \us21/_0739_ ;
wire \us21/_0740_ ;
wire \us21/_0741_ ;
wire \us21/_0742_ ;
wire \us21/_0744_ ;
wire \us21/_0745_ ;
wire \us21/_0746_ ;
wire \us21/_0747_ ;
wire \us21/_0748_ ;
wire \us21/_0749_ ;
wire \us21/_0750_ ;
wire \us21/_0752_ ;
wire \us22/_0008_ ;
wire \us22/_0009_ ;
wire \us22/_0010_ ;
wire \us22/_0011_ ;
wire \us22/_0012_ ;
wire \us22/_0013_ ;
wire \us22/_0014_ ;
wire \us22/_0015_ ;
wire \us22/_0016_ ;
wire \us22/_0017_ ;
wire \us22/_0018_ ;
wire \us22/_0019_ ;
wire \us22/_0020_ ;
wire \us22/_0021_ ;
wire \us22/_0022_ ;
wire \us22/_0023_ ;
wire \us22/_0024_ ;
wire \us22/_0025_ ;
wire \us22/_0026_ ;
wire \us22/_0027_ ;
wire \us22/_0030_ ;
wire \us22/_0032_ ;
wire \us22/_0033_ ;
wire \us22/_0034_ ;
wire \us22/_0035_ ;
wire \us22/_0036_ ;
wire \us22/_0037_ ;
wire \us22/_0038_ ;
wire \us22/_0039_ ;
wire \us22/_0040_ ;
wire \us22/_0041_ ;
wire \us22/_0042_ ;
wire \us22/_0043_ ;
wire \us22/_0045_ ;
wire \us22/_0046_ ;
wire \us22/_0047_ ;
wire \us22/_0049_ ;
wire \us22/_0050_ ;
wire \us22/_0051_ ;
wire \us22/_0052_ ;
wire \us22/_0053_ ;
wire \us22/_0054_ ;
wire \us22/_0056_ ;
wire \us22/_0057_ ;
wire \us22/_0058_ ;
wire \us22/_0060_ ;
wire \us22/_0061_ ;
wire \us22/_0062_ ;
wire \us22/_0064_ ;
wire \us22/_0065_ ;
wire \us22/_0066_ ;
wire \us22/_0067_ ;
wire \us22/_0069_ ;
wire \us22/_0070_ ;
wire \us22/_0072_ ;
wire \us22/_0073_ ;
wire \us22/_0074_ ;
wire \us22/_0075_ ;
wire \us22/_0076_ ;
wire \us22/_0077_ ;
wire \us22/_0078_ ;
wire \us22/_0079_ ;
wire \us22/_0080_ ;
wire \us22/_0081_ ;
wire \us22/_0082_ ;
wire \us22/_0084_ ;
wire \us22/_0085_ ;
wire \us22/_0086_ ;
wire \us22/_0087_ ;
wire \us22/_0088_ ;
wire \us22/_0089_ ;
wire \us22/_0090_ ;
wire \us22/_0091_ ;
wire \us22/_0092_ ;
wire \us22/_0093_ ;
wire \us22/_0094_ ;
wire \us22/_0095_ ;
wire \us22/_0096_ ;
wire \us22/_0097_ ;
wire \us22/_0098_ ;
wire \us22/_0099_ ;
wire \us22/_0100_ ;
wire \us22/_0101_ ;
wire \us22/_0102_ ;
wire \us22/_0103_ ;
wire \us22/_0104_ ;
wire \us22/_0105_ ;
wire \us22/_0106_ ;
wire \us22/_0108_ ;
wire \us22/_0109_ ;
wire \us22/_0110_ ;
wire \us22/_0111_ ;
wire \us22/_0113_ ;
wire \us22/_0114_ ;
wire \us22/_0115_ ;
wire \us22/_0116_ ;
wire \us22/_0117_ ;
wire \us22/_0118_ ;
wire \us22/_0119_ ;
wire \us22/_0120_ ;
wire \us22/_0121_ ;
wire \us22/_0122_ ;
wire \us22/_0123_ ;
wire \us22/_0124_ ;
wire \us22/_0126_ ;
wire \us22/_0127_ ;
wire \us22/_0128_ ;
wire \us22/_0129_ ;
wire \us22/_0130_ ;
wire \us22/_0132_ ;
wire \us22/_0133_ ;
wire \us22/_0134_ ;
wire \us22/_0135_ ;
wire \us22/_0136_ ;
wire \us22/_0137_ ;
wire \us22/_0139_ ;
wire \us22/_0140_ ;
wire \us22/_0141_ ;
wire \us22/_0142_ ;
wire \us22/_0144_ ;
wire \us22/_0145_ ;
wire \us22/_0146_ ;
wire \us22/_0147_ ;
wire \us22/_0148_ ;
wire \us22/_0149_ ;
wire \us22/_0150_ ;
wire \us22/_0151_ ;
wire \us22/_0153_ ;
wire \us22/_0154_ ;
wire \us22/_0155_ ;
wire \us22/_0156_ ;
wire \us22/_0157_ ;
wire \us22/_0158_ ;
wire \us22/_0159_ ;
wire \us22/_0161_ ;
wire \us22/_0162_ ;
wire \us22/_0163_ ;
wire \us22/_0164_ ;
wire \us22/_0165_ ;
wire \us22/_0166_ ;
wire \us22/_0167_ ;
wire \us22/_0168_ ;
wire \us22/_0169_ ;
wire \us22/_0170_ ;
wire \us22/_0171_ ;
wire \us22/_0172_ ;
wire \us22/_0174_ ;
wire \us22/_0175_ ;
wire \us22/_0176_ ;
wire \us22/_0177_ ;
wire \us22/_0178_ ;
wire \us22/_0179_ ;
wire \us22/_0180_ ;
wire \us22/_0181_ ;
wire \us22/_0182_ ;
wire \us22/_0183_ ;
wire \us22/_0184_ ;
wire \us22/_0185_ ;
wire \us22/_0186_ ;
wire \us22/_0187_ ;
wire \us22/_0188_ ;
wire \us22/_0189_ ;
wire \us22/_0190_ ;
wire \us22/_0191_ ;
wire \us22/_0192_ ;
wire \us22/_0193_ ;
wire \us22/_0194_ ;
wire \us22/_0195_ ;
wire \us22/_0196_ ;
wire \us22/_0197_ ;
wire \us22/_0198_ ;
wire \us22/_0199_ ;
wire \us22/_0200_ ;
wire \us22/_0201_ ;
wire \us22/_0202_ ;
wire \us22/_0203_ ;
wire \us22/_0204_ ;
wire \us22/_0205_ ;
wire \us22/_0206_ ;
wire \us22/_0207_ ;
wire \us22/_0208_ ;
wire \us22/_0209_ ;
wire \us22/_0210_ ;
wire \us22/_0211_ ;
wire \us22/_0212_ ;
wire \us22/_0213_ ;
wire \us22/_0214_ ;
wire \us22/_0215_ ;
wire \us22/_0216_ ;
wire \us22/_0217_ ;
wire \us22/_0218_ ;
wire \us22/_0219_ ;
wire \us22/_0220_ ;
wire \us22/_0221_ ;
wire \us22/_0222_ ;
wire \us22/_0223_ ;
wire \us22/_0224_ ;
wire \us22/_0225_ ;
wire \us22/_0226_ ;
wire \us22/_0227_ ;
wire \us22/_0228_ ;
wire \us22/_0229_ ;
wire \us22/_0230_ ;
wire \us22/_0231_ ;
wire \us22/_0232_ ;
wire \us22/_0233_ ;
wire \us22/_0234_ ;
wire \us22/_0235_ ;
wire \us22/_0236_ ;
wire \us22/_0237_ ;
wire \us22/_0238_ ;
wire \us22/_0239_ ;
wire \us22/_0240_ ;
wire \us22/_0241_ ;
wire \us22/_0242_ ;
wire \us22/_0243_ ;
wire \us22/_0244_ ;
wire \us22/_0245_ ;
wire \us22/_0246_ ;
wire \us22/_0247_ ;
wire \us22/_0248_ ;
wire \us22/_0249_ ;
wire \us22/_0250_ ;
wire \us22/_0251_ ;
wire \us22/_0252_ ;
wire \us22/_0253_ ;
wire \us22/_0254_ ;
wire \us22/_0255_ ;
wire \us22/_0256_ ;
wire \us22/_0257_ ;
wire \us22/_0258_ ;
wire \us22/_0259_ ;
wire \us22/_0260_ ;
wire \us22/_0261_ ;
wire \us22/_0263_ ;
wire \us22/_0264_ ;
wire \us22/_0265_ ;
wire \us22/_0266_ ;
wire \us22/_0267_ ;
wire \us22/_0268_ ;
wire \us22/_0269_ ;
wire \us22/_0270_ ;
wire \us22/_0271_ ;
wire \us22/_0272_ ;
wire \us22/_0273_ ;
wire \us22/_0274_ ;
wire \us22/_0275_ ;
wire \us22/_0276_ ;
wire \us22/_0277_ ;
wire \us22/_0278_ ;
wire \us22/_0279_ ;
wire \us22/_0281_ ;
wire \us22/_0283_ ;
wire \us22/_0284_ ;
wire \us22/_0285_ ;
wire \us22/_0286_ ;
wire \us22/_0287_ ;
wire \us22/_0288_ ;
wire \us22/_0289_ ;
wire \us22/_0290_ ;
wire \us22/_0291_ ;
wire \us22/_0293_ ;
wire \us22/_0294_ ;
wire \us22/_0295_ ;
wire \us22/_0296_ ;
wire \us22/_0297_ ;
wire \us22/_0298_ ;
wire \us22/_0299_ ;
wire \us22/_0300_ ;
wire \us22/_0301_ ;
wire \us22/_0302_ ;
wire \us22/_0303_ ;
wire \us22/_0304_ ;
wire \us22/_0305_ ;
wire \us22/_0306_ ;
wire \us22/_0307_ ;
wire \us22/_0308_ ;
wire \us22/_0309_ ;
wire \us22/_0310_ ;
wire \us22/_0311_ ;
wire \us22/_0312_ ;
wire \us22/_0313_ ;
wire \us22/_0314_ ;
wire \us22/_0315_ ;
wire \us22/_0316_ ;
wire \us22/_0317_ ;
wire \us22/_0318_ ;
wire \us22/_0319_ ;
wire \us22/_0320_ ;
wire \us22/_0321_ ;
wire \us22/_0322_ ;
wire \us22/_0323_ ;
wire \us22/_0324_ ;
wire \us22/_0325_ ;
wire \us22/_0326_ ;
wire \us22/_0327_ ;
wire \us22/_0328_ ;
wire \us22/_0329_ ;
wire \us22/_0330_ ;
wire \us22/_0331_ ;
wire \us22/_0332_ ;
wire \us22/_0333_ ;
wire \us22/_0334_ ;
wire \us22/_0335_ ;
wire \us22/_0337_ ;
wire \us22/_0338_ ;
wire \us22/_0339_ ;
wire \us22/_0340_ ;
wire \us22/_0341_ ;
wire \us22/_0342_ ;
wire \us22/_0343_ ;
wire \us22/_0344_ ;
wire \us22/_0345_ ;
wire \us22/_0347_ ;
wire \us22/_0348_ ;
wire \us22/_0349_ ;
wire \us22/_0350_ ;
wire \us22/_0351_ ;
wire \us22/_0352_ ;
wire \us22/_0353_ ;
wire \us22/_0354_ ;
wire \us22/_0355_ ;
wire \us22/_0356_ ;
wire \us22/_0357_ ;
wire \us22/_0358_ ;
wire \us22/_0359_ ;
wire \us22/_0360_ ;
wire \us22/_0361_ ;
wire \us22/_0362_ ;
wire \us22/_0363_ ;
wire \us22/_0365_ ;
wire \us22/_0366_ ;
wire \us22/_0367_ ;
wire \us22/_0368_ ;
wire \us22/_0370_ ;
wire \us22/_0371_ ;
wire \us22/_0372_ ;
wire \us22/_0373_ ;
wire \us22/_0374_ ;
wire \us22/_0375_ ;
wire \us22/_0376_ ;
wire \us22/_0377_ ;
wire \us22/_0378_ ;
wire \us22/_0379_ ;
wire \us22/_0380_ ;
wire \us22/_0381_ ;
wire \us22/_0382_ ;
wire \us22/_0383_ ;
wire \us22/_0384_ ;
wire \us22/_0385_ ;
wire \us22/_0386_ ;
wire \us22/_0387_ ;
wire \us22/_0388_ ;
wire \us22/_0389_ ;
wire \us22/_0390_ ;
wire \us22/_0391_ ;
wire \us22/_0392_ ;
wire \us22/_0393_ ;
wire \us22/_0394_ ;
wire \us22/_0395_ ;
wire \us22/_0396_ ;
wire \us22/_0397_ ;
wire \us22/_0398_ ;
wire \us22/_0399_ ;
wire \us22/_0400_ ;
wire \us22/_0401_ ;
wire \us22/_0402_ ;
wire \us22/_0403_ ;
wire \us22/_0404_ ;
wire \us22/_0405_ ;
wire \us22/_0406_ ;
wire \us22/_0407_ ;
wire \us22/_0408_ ;
wire \us22/_0409_ ;
wire \us22/_0410_ ;
wire \us22/_0411_ ;
wire \us22/_0412_ ;
wire \us22/_0413_ ;
wire \us22/_0414_ ;
wire \us22/_0415_ ;
wire \us22/_0416_ ;
wire \us22/_0417_ ;
wire \us22/_0418_ ;
wire \us22/_0419_ ;
wire \us22/_0420_ ;
wire \us22/_0421_ ;
wire \us22/_0422_ ;
wire \us22/_0423_ ;
wire \us22/_0424_ ;
wire \us22/_0425_ ;
wire \us22/_0426_ ;
wire \us22/_0427_ ;
wire \us22/_0428_ ;
wire \us22/_0429_ ;
wire \us22/_0430_ ;
wire \us22/_0431_ ;
wire \us22/_0432_ ;
wire \us22/_0433_ ;
wire \us22/_0434_ ;
wire \us22/_0435_ ;
wire \us22/_0436_ ;
wire \us22/_0437_ ;
wire \us22/_0438_ ;
wire \us22/_0439_ ;
wire \us22/_0440_ ;
wire \us22/_0441_ ;
wire \us22/_0442_ ;
wire \us22/_0443_ ;
wire \us22/_0444_ ;
wire \us22/_0446_ ;
wire \us22/_0447_ ;
wire \us22/_0448_ ;
wire \us22/_0449_ ;
wire \us22/_0450_ ;
wire \us22/_0451_ ;
wire \us22/_0452_ ;
wire \us22/_0453_ ;
wire \us22/_0454_ ;
wire \us22/_0455_ ;
wire \us22/_0457_ ;
wire \us22/_0458_ ;
wire \us22/_0459_ ;
wire \us22/_0460_ ;
wire \us22/_0461_ ;
wire \us22/_0462_ ;
wire \us22/_0463_ ;
wire \us22/_0464_ ;
wire \us22/_0465_ ;
wire \us22/_0466_ ;
wire \us22/_0467_ ;
wire \us22/_0468_ ;
wire \us22/_0469_ ;
wire \us22/_0470_ ;
wire \us22/_0471_ ;
wire \us22/_0472_ ;
wire \us22/_0473_ ;
wire \us22/_0474_ ;
wire \us22/_0475_ ;
wire \us22/_0476_ ;
wire \us22/_0477_ ;
wire \us22/_0478_ ;
wire \us22/_0479_ ;
wire \us22/_0480_ ;
wire \us22/_0481_ ;
wire \us22/_0482_ ;
wire \us22/_0483_ ;
wire \us22/_0484_ ;
wire \us22/_0485_ ;
wire \us22/_0486_ ;
wire \us22/_0487_ ;
wire \us22/_0488_ ;
wire \us22/_0490_ ;
wire \us22/_0491_ ;
wire \us22/_0492_ ;
wire \us22/_0493_ ;
wire \us22/_0494_ ;
wire \us22/_0495_ ;
wire \us22/_0496_ ;
wire \us22/_0497_ ;
wire \us22/_0498_ ;
wire \us22/_0500_ ;
wire \us22/_0501_ ;
wire \us22/_0502_ ;
wire \us22/_0503_ ;
wire \us22/_0504_ ;
wire \us22/_0505_ ;
wire \us22/_0506_ ;
wire \us22/_0507_ ;
wire \us22/_0508_ ;
wire \us22/_0509_ ;
wire \us22/_0510_ ;
wire \us22/_0511_ ;
wire \us22/_0512_ ;
wire \us22/_0513_ ;
wire \us22/_0514_ ;
wire \us22/_0515_ ;
wire \us22/_0516_ ;
wire \us22/_0517_ ;
wire \us22/_0518_ ;
wire \us22/_0519_ ;
wire \us22/_0520_ ;
wire \us22/_0521_ ;
wire \us22/_0522_ ;
wire \us22/_0523_ ;
wire \us22/_0524_ ;
wire \us22/_0525_ ;
wire \us22/_0526_ ;
wire \us22/_0527_ ;
wire \us22/_0528_ ;
wire \us22/_0529_ ;
wire \us22/_0530_ ;
wire \us22/_0531_ ;
wire \us22/_0532_ ;
wire \us22/_0533_ ;
wire \us22/_0534_ ;
wire \us22/_0535_ ;
wire \us22/_0536_ ;
wire \us22/_0537_ ;
wire \us22/_0538_ ;
wire \us22/_0539_ ;
wire \us22/_0540_ ;
wire \us22/_0541_ ;
wire \us22/_0542_ ;
wire \us22/_0543_ ;
wire \us22/_0544_ ;
wire \us22/_0545_ ;
wire \us22/_0546_ ;
wire \us22/_0547_ ;
wire \us22/_0548_ ;
wire \us22/_0549_ ;
wire \us22/_0550_ ;
wire \us22/_0551_ ;
wire \us22/_0552_ ;
wire \us22/_0553_ ;
wire \us22/_0554_ ;
wire \us22/_0555_ ;
wire \us22/_0556_ ;
wire \us22/_0557_ ;
wire \us22/_0558_ ;
wire \us22/_0559_ ;
wire \us22/_0560_ ;
wire \us22/_0561_ ;
wire \us22/_0562_ ;
wire \us22/_0563_ ;
wire \us22/_0565_ ;
wire \us22/_0566_ ;
wire \us22/_0567_ ;
wire \us22/_0568_ ;
wire \us22/_0569_ ;
wire \us22/_0570_ ;
wire \us22/_0571_ ;
wire \us22/_0572_ ;
wire \us22/_0573_ ;
wire \us22/_0574_ ;
wire \us22/_0575_ ;
wire \us22/_0576_ ;
wire \us22/_0577_ ;
wire \us22/_0578_ ;
wire \us22/_0579_ ;
wire \us22/_0580_ ;
wire \us22/_0581_ ;
wire \us22/_0582_ ;
wire \us22/_0583_ ;
wire \us22/_0584_ ;
wire \us22/_0585_ ;
wire \us22/_0586_ ;
wire \us22/_0587_ ;
wire \us22/_0588_ ;
wire \us22/_0589_ ;
wire \us22/_0590_ ;
wire \us22/_0591_ ;
wire \us22/_0592_ ;
wire \us22/_0593_ ;
wire \us22/_0594_ ;
wire \us22/_0595_ ;
wire \us22/_0596_ ;
wire \us22/_0598_ ;
wire \us22/_0599_ ;
wire \us22/_0600_ ;
wire \us22/_0601_ ;
wire \us22/_0602_ ;
wire \us22/_0603_ ;
wire \us22/_0604_ ;
wire \us22/_0605_ ;
wire \us22/_0606_ ;
wire \us22/_0607_ ;
wire \us22/_0608_ ;
wire \us22/_0609_ ;
wire \us22/_0610_ ;
wire \us22/_0611_ ;
wire \us22/_0612_ ;
wire \us22/_0613_ ;
wire \us22/_0614_ ;
wire \us22/_0615_ ;
wire \us22/_0616_ ;
wire \us22/_0617_ ;
wire \us22/_0618_ ;
wire \us22/_0619_ ;
wire \us22/_0620_ ;
wire \us22/_0621_ ;
wire \us22/_0622_ ;
wire \us22/_0623_ ;
wire \us22/_0624_ ;
wire \us22/_0625_ ;
wire \us22/_0626_ ;
wire \us22/_0627_ ;
wire \us22/_0628_ ;
wire \us22/_0629_ ;
wire \us22/_0630_ ;
wire \us22/_0631_ ;
wire \us22/_0632_ ;
wire \us22/_0633_ ;
wire \us22/_0634_ ;
wire \us22/_0635_ ;
wire \us22/_0636_ ;
wire \us22/_0637_ ;
wire \us22/_0638_ ;
wire \us22/_0639_ ;
wire \us22/_0640_ ;
wire \us22/_0641_ ;
wire \us22/_0642_ ;
wire \us22/_0643_ ;
wire \us22/_0644_ ;
wire \us22/_0645_ ;
wire \us22/_0646_ ;
wire \us22/_0647_ ;
wire \us22/_0648_ ;
wire \us22/_0649_ ;
wire \us22/_0650_ ;
wire \us22/_0651_ ;
wire \us22/_0652_ ;
wire \us22/_0653_ ;
wire \us22/_0654_ ;
wire \us22/_0655_ ;
wire \us22/_0656_ ;
wire \us22/_0657_ ;
wire \us22/_0658_ ;
wire \us22/_0659_ ;
wire \us22/_0660_ ;
wire \us22/_0661_ ;
wire \us22/_0662_ ;
wire \us22/_0663_ ;
wire \us22/_0664_ ;
wire \us22/_0665_ ;
wire \us22/_0666_ ;
wire \us22/_0667_ ;
wire \us22/_0668_ ;
wire \us22/_0669_ ;
wire \us22/_0670_ ;
wire \us22/_0671_ ;
wire \us22/_0672_ ;
wire \us22/_0673_ ;
wire \us22/_0674_ ;
wire \us22/_0675_ ;
wire \us22/_0676_ ;
wire \us22/_0677_ ;
wire \us22/_0678_ ;
wire \us22/_0679_ ;
wire \us22/_0680_ ;
wire \us22/_0681_ ;
wire \us22/_0682_ ;
wire \us22/_0683_ ;
wire \us22/_0684_ ;
wire \us22/_0685_ ;
wire \us22/_0686_ ;
wire \us22/_0687_ ;
wire \us22/_0688_ ;
wire \us22/_0689_ ;
wire \us22/_0690_ ;
wire \us22/_0691_ ;
wire \us22/_0692_ ;
wire \us22/_0693_ ;
wire \us22/_0694_ ;
wire \us22/_0695_ ;
wire \us22/_0696_ ;
wire \us22/_0697_ ;
wire \us22/_0698_ ;
wire \us22/_0699_ ;
wire \us22/_0700_ ;
wire \us22/_0701_ ;
wire \us22/_0702_ ;
wire \us22/_0703_ ;
wire \us22/_0704_ ;
wire \us22/_0705_ ;
wire \us22/_0706_ ;
wire \us22/_0707_ ;
wire \us22/_0708_ ;
wire \us22/_0709_ ;
wire \us22/_0710_ ;
wire \us22/_0711_ ;
wire \us22/_0712_ ;
wire \us22/_0713_ ;
wire \us22/_0714_ ;
wire \us22/_0715_ ;
wire \us22/_0717_ ;
wire \us22/_0718_ ;
wire \us22/_0719_ ;
wire \us22/_0720_ ;
wire \us22/_0721_ ;
wire \us22/_0722_ ;
wire \us22/_0723_ ;
wire \us22/_0724_ ;
wire \us22/_0725_ ;
wire \us22/_0726_ ;
wire \us22/_0727_ ;
wire \us22/_0728_ ;
wire \us22/_0729_ ;
wire \us22/_0730_ ;
wire \us22/_0731_ ;
wire \us22/_0732_ ;
wire \us22/_0733_ ;
wire \us22/_0734_ ;
wire \us22/_0735_ ;
wire \us22/_0736_ ;
wire \us22/_0738_ ;
wire \us22/_0739_ ;
wire \us22/_0740_ ;
wire \us22/_0741_ ;
wire \us22/_0742_ ;
wire \us22/_0744_ ;
wire \us22/_0745_ ;
wire \us22/_0746_ ;
wire \us22/_0747_ ;
wire \us22/_0748_ ;
wire \us22/_0749_ ;
wire \us22/_0750_ ;
wire \us22/_0752_ ;
wire \us23/_0008_ ;
wire \us23/_0009_ ;
wire \us23/_0010_ ;
wire \us23/_0011_ ;
wire \us23/_0012_ ;
wire \us23/_0013_ ;
wire \us23/_0014_ ;
wire \us23/_0015_ ;
wire \us23/_0016_ ;
wire \us23/_0017_ ;
wire \us23/_0019_ ;
wire \us23/_0020_ ;
wire \us23/_0022_ ;
wire \us23/_0024_ ;
wire \us23/_0025_ ;
wire \us23/_0026_ ;
wire \us23/_0027_ ;
wire \us23/_0030_ ;
wire \us23/_0032_ ;
wire \us23/_0033_ ;
wire \us23/_0034_ ;
wire \us23/_0035_ ;
wire \us23/_0037_ ;
wire \us23/_0038_ ;
wire \us23/_0039_ ;
wire \us23/_0040_ ;
wire \us23/_0041_ ;
wire \us23/_0042_ ;
wire \us23/_0043_ ;
wire \us23/_0045_ ;
wire \us23/_0046_ ;
wire \us23/_0047_ ;
wire \us23/_0049_ ;
wire \us23/_0050_ ;
wire \us23/_0051_ ;
wire \us23/_0052_ ;
wire \us23/_0053_ ;
wire \us23/_0054_ ;
wire \us23/_0056_ ;
wire \us23/_0057_ ;
wire \us23/_0058_ ;
wire \us23/_0060_ ;
wire \us23/_0061_ ;
wire \us23/_0062_ ;
wire \us23/_0064_ ;
wire \us23/_0065_ ;
wire \us23/_0066_ ;
wire \us23/_0067_ ;
wire \us23/_0069_ ;
wire \us23/_0070_ ;
wire \us23/_0072_ ;
wire \us23/_0073_ ;
wire \us23/_0074_ ;
wire \us23/_0075_ ;
wire \us23/_0076_ ;
wire \us23/_0077_ ;
wire \us23/_0078_ ;
wire \us23/_0079_ ;
wire \us23/_0081_ ;
wire \us23/_0082_ ;
wire \us23/_0085_ ;
wire \us23/_0086_ ;
wire \us23/_0087_ ;
wire \us23/_0088_ ;
wire \us23/_0089_ ;
wire \us23/_0090_ ;
wire \us23/_0091_ ;
wire \us23/_0092_ ;
wire \us23/_0093_ ;
wire \us23/_0094_ ;
wire \us23/_0095_ ;
wire \us23/_0096_ ;
wire \us23/_0097_ ;
wire \us23/_0098_ ;
wire \us23/_0099_ ;
wire \us23/_0100_ ;
wire \us23/_0101_ ;
wire \us23/_0102_ ;
wire \us23/_0103_ ;
wire \us23/_0104_ ;
wire \us23/_0105_ ;
wire \us23/_0106_ ;
wire \us23/_0108_ ;
wire \us23/_0109_ ;
wire \us23/_0110_ ;
wire \us23/_0111_ ;
wire \us23/_0113_ ;
wire \us23/_0114_ ;
wire \us23/_0115_ ;
wire \us23/_0116_ ;
wire \us23/_0117_ ;
wire \us23/_0118_ ;
wire \us23/_0119_ ;
wire \us23/_0120_ ;
wire \us23/_0121_ ;
wire \us23/_0122_ ;
wire \us23/_0123_ ;
wire \us23/_0124_ ;
wire \us23/_0126_ ;
wire \us23/_0127_ ;
wire \us23/_0128_ ;
wire \us23/_0129_ ;
wire \us23/_0130_ ;
wire \us23/_0132_ ;
wire \us23/_0133_ ;
wire \us23/_0134_ ;
wire \us23/_0135_ ;
wire \us23/_0136_ ;
wire \us23/_0137_ ;
wire \us23/_0139_ ;
wire \us23/_0140_ ;
wire \us23/_0141_ ;
wire \us23/_0142_ ;
wire \us23/_0144_ ;
wire \us23/_0145_ ;
wire \us23/_0146_ ;
wire \us23/_0147_ ;
wire \us23/_0148_ ;
wire \us23/_0149_ ;
wire \us23/_0150_ ;
wire \us23/_0151_ ;
wire \us23/_0153_ ;
wire \us23/_0154_ ;
wire \us23/_0155_ ;
wire \us23/_0156_ ;
wire \us23/_0157_ ;
wire \us23/_0158_ ;
wire \us23/_0159_ ;
wire \us23/_0161_ ;
wire \us23/_0162_ ;
wire \us23/_0163_ ;
wire \us23/_0164_ ;
wire \us23/_0165_ ;
wire \us23/_0166_ ;
wire \us23/_0167_ ;
wire \us23/_0168_ ;
wire \us23/_0169_ ;
wire \us23/_0170_ ;
wire \us23/_0171_ ;
wire \us23/_0172_ ;
wire \us23/_0174_ ;
wire \us23/_0175_ ;
wire \us23/_0176_ ;
wire \us23/_0177_ ;
wire \us23/_0178_ ;
wire \us23/_0179_ ;
wire \us23/_0180_ ;
wire \us23/_0181_ ;
wire \us23/_0182_ ;
wire \us23/_0183_ ;
wire \us23/_0184_ ;
wire \us23/_0185_ ;
wire \us23/_0186_ ;
wire \us23/_0187_ ;
wire \us23/_0188_ ;
wire \us23/_0189_ ;
wire \us23/_0190_ ;
wire \us23/_0191_ ;
wire \us23/_0192_ ;
wire \us23/_0193_ ;
wire \us23/_0194_ ;
wire \us23/_0195_ ;
wire \us23/_0196_ ;
wire \us23/_0197_ ;
wire \us23/_0198_ ;
wire \us23/_0199_ ;
wire \us23/_0200_ ;
wire \us23/_0201_ ;
wire \us23/_0202_ ;
wire \us23/_0203_ ;
wire \us23/_0204_ ;
wire \us23/_0205_ ;
wire \us23/_0206_ ;
wire \us23/_0207_ ;
wire \us23/_0208_ ;
wire \us23/_0209_ ;
wire \us23/_0210_ ;
wire \us23/_0211_ ;
wire \us23/_0212_ ;
wire \us23/_0213_ ;
wire \us23/_0214_ ;
wire \us23/_0215_ ;
wire \us23/_0217_ ;
wire \us23/_0218_ ;
wire \us23/_0219_ ;
wire \us23/_0220_ ;
wire \us23/_0221_ ;
wire \us23/_0222_ ;
wire \us23/_0223_ ;
wire \us23/_0224_ ;
wire \us23/_0225_ ;
wire \us23/_0226_ ;
wire \us23/_0227_ ;
wire \us23/_0228_ ;
wire \us23/_0229_ ;
wire \us23/_0230_ ;
wire \us23/_0231_ ;
wire \us23/_0232_ ;
wire \us23/_0233_ ;
wire \us23/_0234_ ;
wire \us23/_0235_ ;
wire \us23/_0236_ ;
wire \us23/_0237_ ;
wire \us23/_0238_ ;
wire \us23/_0239_ ;
wire \us23/_0240_ ;
wire \us23/_0241_ ;
wire \us23/_0242_ ;
wire \us23/_0243_ ;
wire \us23/_0244_ ;
wire \us23/_0245_ ;
wire \us23/_0246_ ;
wire \us23/_0247_ ;
wire \us23/_0248_ ;
wire \us23/_0249_ ;
wire \us23/_0250_ ;
wire \us23/_0251_ ;
wire \us23/_0252_ ;
wire \us23/_0253_ ;
wire \us23/_0254_ ;
wire \us23/_0255_ ;
wire \us23/_0256_ ;
wire \us23/_0257_ ;
wire \us23/_0258_ ;
wire \us23/_0259_ ;
wire \us23/_0260_ ;
wire \us23/_0261_ ;
wire \us23/_0263_ ;
wire \us23/_0264_ ;
wire \us23/_0265_ ;
wire \us23/_0266_ ;
wire \us23/_0267_ ;
wire \us23/_0268_ ;
wire \us23/_0269_ ;
wire \us23/_0270_ ;
wire \us23/_0271_ ;
wire \us23/_0272_ ;
wire \us23/_0273_ ;
wire \us23/_0274_ ;
wire \us23/_0275_ ;
wire \us23/_0276_ ;
wire \us23/_0277_ ;
wire \us23/_0278_ ;
wire \us23/_0279_ ;
wire \us23/_0280_ ;
wire \us23/_0281_ ;
wire \us23/_0283_ ;
wire \us23/_0284_ ;
wire \us23/_0285_ ;
wire \us23/_0286_ ;
wire \us23/_0287_ ;
wire \us23/_0288_ ;
wire \us23/_0289_ ;
wire \us23/_0290_ ;
wire \us23/_0291_ ;
wire \us23/_0293_ ;
wire \us23/_0294_ ;
wire \us23/_0295_ ;
wire \us23/_0296_ ;
wire \us23/_0297_ ;
wire \us23/_0298_ ;
wire \us23/_0299_ ;
wire \us23/_0300_ ;
wire \us23/_0301_ ;
wire \us23/_0302_ ;
wire \us23/_0303_ ;
wire \us23/_0304_ ;
wire \us23/_0305_ ;
wire \us23/_0306_ ;
wire \us23/_0307_ ;
wire \us23/_0308_ ;
wire \us23/_0309_ ;
wire \us23/_0310_ ;
wire \us23/_0311_ ;
wire \us23/_0312_ ;
wire \us23/_0313_ ;
wire \us23/_0314_ ;
wire \us23/_0315_ ;
wire \us23/_0316_ ;
wire \us23/_0317_ ;
wire \us23/_0318_ ;
wire \us23/_0319_ ;
wire \us23/_0320_ ;
wire \us23/_0321_ ;
wire \us23/_0322_ ;
wire \us23/_0323_ ;
wire \us23/_0324_ ;
wire \us23/_0325_ ;
wire \us23/_0326_ ;
wire \us23/_0327_ ;
wire \us23/_0328_ ;
wire \us23/_0329_ ;
wire \us23/_0330_ ;
wire \us23/_0331_ ;
wire \us23/_0332_ ;
wire \us23/_0333_ ;
wire \us23/_0334_ ;
wire \us23/_0335_ ;
wire \us23/_0337_ ;
wire \us23/_0338_ ;
wire \us23/_0339_ ;
wire \us23/_0340_ ;
wire \us23/_0341_ ;
wire \us23/_0342_ ;
wire \us23/_0343_ ;
wire \us23/_0344_ ;
wire \us23/_0345_ ;
wire \us23/_0347_ ;
wire \us23/_0348_ ;
wire \us23/_0349_ ;
wire \us23/_0350_ ;
wire \us23/_0351_ ;
wire \us23/_0352_ ;
wire \us23/_0353_ ;
wire \us23/_0354_ ;
wire \us23/_0355_ ;
wire \us23/_0356_ ;
wire \us23/_0357_ ;
wire \us23/_0358_ ;
wire \us23/_0359_ ;
wire \us23/_0360_ ;
wire \us23/_0361_ ;
wire \us23/_0362_ ;
wire \us23/_0363_ ;
wire \us23/_0365_ ;
wire \us23/_0366_ ;
wire \us23/_0367_ ;
wire \us23/_0368_ ;
wire \us23/_0370_ ;
wire \us23/_0371_ ;
wire \us23/_0372_ ;
wire \us23/_0373_ ;
wire \us23/_0374_ ;
wire \us23/_0375_ ;
wire \us23/_0376_ ;
wire \us23/_0377_ ;
wire \us23/_0378_ ;
wire \us23/_0379_ ;
wire \us23/_0380_ ;
wire \us23/_0381_ ;
wire \us23/_0382_ ;
wire \us23/_0383_ ;
wire \us23/_0384_ ;
wire \us23/_0385_ ;
wire \us23/_0386_ ;
wire \us23/_0387_ ;
wire \us23/_0388_ ;
wire \us23/_0389_ ;
wire \us23/_0390_ ;
wire \us23/_0391_ ;
wire \us23/_0392_ ;
wire \us23/_0393_ ;
wire \us23/_0394_ ;
wire \us23/_0395_ ;
wire \us23/_0396_ ;
wire \us23/_0397_ ;
wire \us23/_0398_ ;
wire \us23/_0399_ ;
wire \us23/_0400_ ;
wire \us23/_0401_ ;
wire \us23/_0402_ ;
wire \us23/_0403_ ;
wire \us23/_0404_ ;
wire \us23/_0405_ ;
wire \us23/_0406_ ;
wire \us23/_0407_ ;
wire \us23/_0408_ ;
wire \us23/_0409_ ;
wire \us23/_0410_ ;
wire \us23/_0411_ ;
wire \us23/_0412_ ;
wire \us23/_0413_ ;
wire \us23/_0414_ ;
wire \us23/_0415_ ;
wire \us23/_0416_ ;
wire \us23/_0417_ ;
wire \us23/_0418_ ;
wire \us23/_0419_ ;
wire \us23/_0420_ ;
wire \us23/_0421_ ;
wire \us23/_0422_ ;
wire \us23/_0423_ ;
wire \us23/_0424_ ;
wire \us23/_0425_ ;
wire \us23/_0426_ ;
wire \us23/_0427_ ;
wire \us23/_0428_ ;
wire \us23/_0429_ ;
wire \us23/_0430_ ;
wire \us23/_0431_ ;
wire \us23/_0432_ ;
wire \us23/_0433_ ;
wire \us23/_0434_ ;
wire \us23/_0435_ ;
wire \us23/_0436_ ;
wire \us23/_0437_ ;
wire \us23/_0438_ ;
wire \us23/_0439_ ;
wire \us23/_0440_ ;
wire \us23/_0441_ ;
wire \us23/_0442_ ;
wire \us23/_0443_ ;
wire \us23/_0444_ ;
wire \us23/_0446_ ;
wire \us23/_0447_ ;
wire \us23/_0448_ ;
wire \us23/_0449_ ;
wire \us23/_0450_ ;
wire \us23/_0451_ ;
wire \us23/_0452_ ;
wire \us23/_0453_ ;
wire \us23/_0454_ ;
wire \us23/_0455_ ;
wire \us23/_0457_ ;
wire \us23/_0458_ ;
wire \us23/_0459_ ;
wire \us23/_0460_ ;
wire \us23/_0461_ ;
wire \us23/_0462_ ;
wire \us23/_0463_ ;
wire \us23/_0464_ ;
wire \us23/_0465_ ;
wire \us23/_0466_ ;
wire \us23/_0467_ ;
wire \us23/_0468_ ;
wire \us23/_0469_ ;
wire \us23/_0470_ ;
wire \us23/_0471_ ;
wire \us23/_0472_ ;
wire \us23/_0473_ ;
wire \us23/_0474_ ;
wire \us23/_0475_ ;
wire \us23/_0476_ ;
wire \us23/_0477_ ;
wire \us23/_0478_ ;
wire \us23/_0479_ ;
wire \us23/_0480_ ;
wire \us23/_0481_ ;
wire \us23/_0482_ ;
wire \us23/_0483_ ;
wire \us23/_0484_ ;
wire \us23/_0485_ ;
wire \us23/_0486_ ;
wire \us23/_0487_ ;
wire \us23/_0488_ ;
wire \us23/_0490_ ;
wire \us23/_0491_ ;
wire \us23/_0492_ ;
wire \us23/_0493_ ;
wire \us23/_0494_ ;
wire \us23/_0495_ ;
wire \us23/_0496_ ;
wire \us23/_0497_ ;
wire \us23/_0498_ ;
wire \us23/_0500_ ;
wire \us23/_0501_ ;
wire \us23/_0502_ ;
wire \us23/_0503_ ;
wire \us23/_0504_ ;
wire \us23/_0505_ ;
wire \us23/_0506_ ;
wire \us23/_0507_ ;
wire \us23/_0508_ ;
wire \us23/_0509_ ;
wire \us23/_0510_ ;
wire \us23/_0511_ ;
wire \us23/_0512_ ;
wire \us23/_0513_ ;
wire \us23/_0514_ ;
wire \us23/_0515_ ;
wire \us23/_0516_ ;
wire \us23/_0517_ ;
wire \us23/_0518_ ;
wire \us23/_0519_ ;
wire \us23/_0520_ ;
wire \us23/_0521_ ;
wire \us23/_0522_ ;
wire \us23/_0523_ ;
wire \us23/_0524_ ;
wire \us23/_0525_ ;
wire \us23/_0526_ ;
wire \us23/_0527_ ;
wire \us23/_0528_ ;
wire \us23/_0529_ ;
wire \us23/_0530_ ;
wire \us23/_0531_ ;
wire \us23/_0532_ ;
wire \us23/_0533_ ;
wire \us23/_0534_ ;
wire \us23/_0535_ ;
wire \us23/_0536_ ;
wire \us23/_0537_ ;
wire \us23/_0538_ ;
wire \us23/_0539_ ;
wire \us23/_0540_ ;
wire \us23/_0541_ ;
wire \us23/_0542_ ;
wire \us23/_0543_ ;
wire \us23/_0544_ ;
wire \us23/_0545_ ;
wire \us23/_0546_ ;
wire \us23/_0547_ ;
wire \us23/_0548_ ;
wire \us23/_0549_ ;
wire \us23/_0550_ ;
wire \us23/_0551_ ;
wire \us23/_0552_ ;
wire \us23/_0553_ ;
wire \us23/_0554_ ;
wire \us23/_0555_ ;
wire \us23/_0556_ ;
wire \us23/_0557_ ;
wire \us23/_0558_ ;
wire \us23/_0559_ ;
wire \us23/_0560_ ;
wire \us23/_0561_ ;
wire \us23/_0562_ ;
wire \us23/_0563_ ;
wire \us23/_0565_ ;
wire \us23/_0566_ ;
wire \us23/_0567_ ;
wire \us23/_0568_ ;
wire \us23/_0569_ ;
wire \us23/_0570_ ;
wire \us23/_0571_ ;
wire \us23/_0572_ ;
wire \us23/_0573_ ;
wire \us23/_0574_ ;
wire \us23/_0575_ ;
wire \us23/_0576_ ;
wire \us23/_0577_ ;
wire \us23/_0578_ ;
wire \us23/_0579_ ;
wire \us23/_0580_ ;
wire \us23/_0581_ ;
wire \us23/_0582_ ;
wire \us23/_0583_ ;
wire \us23/_0584_ ;
wire \us23/_0585_ ;
wire \us23/_0586_ ;
wire \us23/_0587_ ;
wire \us23/_0588_ ;
wire \us23/_0589_ ;
wire \us23/_0590_ ;
wire \us23/_0591_ ;
wire \us23/_0592_ ;
wire \us23/_0593_ ;
wire \us23/_0594_ ;
wire \us23/_0595_ ;
wire \us23/_0596_ ;
wire \us23/_0598_ ;
wire \us23/_0599_ ;
wire \us23/_0600_ ;
wire \us23/_0601_ ;
wire \us23/_0602_ ;
wire \us23/_0603_ ;
wire \us23/_0604_ ;
wire \us23/_0605_ ;
wire \us23/_0606_ ;
wire \us23/_0607_ ;
wire \us23/_0608_ ;
wire \us23/_0609_ ;
wire \us23/_0610_ ;
wire \us23/_0611_ ;
wire \us23/_0612_ ;
wire \us23/_0613_ ;
wire \us23/_0614_ ;
wire \us23/_0615_ ;
wire \us23/_0616_ ;
wire \us23/_0617_ ;
wire \us23/_0618_ ;
wire \us23/_0619_ ;
wire \us23/_0620_ ;
wire \us23/_0621_ ;
wire \us23/_0622_ ;
wire \us23/_0623_ ;
wire \us23/_0624_ ;
wire \us23/_0625_ ;
wire \us23/_0626_ ;
wire \us23/_0627_ ;
wire \us23/_0628_ ;
wire \us23/_0629_ ;
wire \us23/_0630_ ;
wire \us23/_0631_ ;
wire \us23/_0632_ ;
wire \us23/_0633_ ;
wire \us23/_0634_ ;
wire \us23/_0635_ ;
wire \us23/_0636_ ;
wire \us23/_0637_ ;
wire \us23/_0638_ ;
wire \us23/_0639_ ;
wire \us23/_0640_ ;
wire \us23/_0641_ ;
wire \us23/_0642_ ;
wire \us23/_0643_ ;
wire \us23/_0644_ ;
wire \us23/_0645_ ;
wire \us23/_0646_ ;
wire \us23/_0647_ ;
wire \us23/_0648_ ;
wire \us23/_0649_ ;
wire \us23/_0650_ ;
wire \us23/_0652_ ;
wire \us23/_0653_ ;
wire \us23/_0654_ ;
wire \us23/_0655_ ;
wire \us23/_0656_ ;
wire \us23/_0657_ ;
wire \us23/_0658_ ;
wire \us23/_0659_ ;
wire \us23/_0660_ ;
wire \us23/_0661_ ;
wire \us23/_0662_ ;
wire \us23/_0663_ ;
wire \us23/_0664_ ;
wire \us23/_0665_ ;
wire \us23/_0666_ ;
wire \us23/_0667_ ;
wire \us23/_0668_ ;
wire \us23/_0669_ ;
wire \us23/_0670_ ;
wire \us23/_0671_ ;
wire \us23/_0673_ ;
wire \us23/_0674_ ;
wire \us23/_0675_ ;
wire \us23/_0676_ ;
wire \us23/_0677_ ;
wire \us23/_0678_ ;
wire \us23/_0679_ ;
wire \us23/_0680_ ;
wire \us23/_0681_ ;
wire \us23/_0682_ ;
wire \us23/_0683_ ;
wire \us23/_0684_ ;
wire \us23/_0685_ ;
wire \us23/_0686_ ;
wire \us23/_0687_ ;
wire \us23/_0688_ ;
wire \us23/_0689_ ;
wire \us23/_0690_ ;
wire \us23/_0691_ ;
wire \us23/_0692_ ;
wire \us23/_0693_ ;
wire \us23/_0694_ ;
wire \us23/_0695_ ;
wire \us23/_0696_ ;
wire \us23/_0697_ ;
wire \us23/_0698_ ;
wire \us23/_0699_ ;
wire \us23/_0700_ ;
wire \us23/_0701_ ;
wire \us23/_0702_ ;
wire \us23/_0703_ ;
wire \us23/_0704_ ;
wire \us23/_0705_ ;
wire \us23/_0706_ ;
wire \us23/_0707_ ;
wire \us23/_0708_ ;
wire \us23/_0709_ ;
wire \us23/_0710_ ;
wire \us23/_0711_ ;
wire \us23/_0712_ ;
wire \us23/_0713_ ;
wire \us23/_0714_ ;
wire \us23/_0715_ ;
wire \us23/_0717_ ;
wire \us23/_0718_ ;
wire \us23/_0719_ ;
wire \us23/_0720_ ;
wire \us23/_0721_ ;
wire \us23/_0722_ ;
wire \us23/_0723_ ;
wire \us23/_0724_ ;
wire \us23/_0725_ ;
wire \us23/_0726_ ;
wire \us23/_0727_ ;
wire \us23/_0728_ ;
wire \us23/_0729_ ;
wire \us23/_0730_ ;
wire \us23/_0731_ ;
wire \us23/_0733_ ;
wire \us23/_0734_ ;
wire \us23/_0735_ ;
wire \us23/_0736_ ;
wire \us23/_0738_ ;
wire \us23/_0739_ ;
wire \us23/_0740_ ;
wire \us23/_0741_ ;
wire \us23/_0742_ ;
wire \us23/_0744_ ;
wire \us23/_0745_ ;
wire \us23/_0746_ ;
wire \us23/_0748_ ;
wire \us23/_0749_ ;
wire \us23/_0750_ ;
wire \us23/_0752_ ;
wire \us30/_0008_ ;
wire \us30/_0009_ ;
wire \us30/_0010_ ;
wire \us30/_0011_ ;
wire \us30/_0012_ ;
wire \us30/_0013_ ;
wire \us30/_0014_ ;
wire \us30/_0015_ ;
wire \us30/_0016_ ;
wire \us30/_0017_ ;
wire \us30/_0019_ ;
wire \us30/_0020_ ;
wire \us30/_0022_ ;
wire \us30/_0024_ ;
wire \us30/_0025_ ;
wire \us30/_0026_ ;
wire \us30/_0027_ ;
wire \us30/_0030_ ;
wire \us30/_0032_ ;
wire \us30/_0033_ ;
wire \us30/_0034_ ;
wire \us30/_0035_ ;
wire \us30/_0037_ ;
wire \us30/_0038_ ;
wire \us30/_0039_ ;
wire \us30/_0040_ ;
wire \us30/_0041_ ;
wire \us30/_0042_ ;
wire \us30/_0043_ ;
wire \us30/_0045_ ;
wire \us30/_0046_ ;
wire \us30/_0047_ ;
wire \us30/_0049_ ;
wire \us30/_0050_ ;
wire \us30/_0051_ ;
wire \us30/_0052_ ;
wire \us30/_0053_ ;
wire \us30/_0054_ ;
wire \us30/_0057_ ;
wire \us30/_0058_ ;
wire \us30/_0060_ ;
wire \us30/_0061_ ;
wire \us30/_0062_ ;
wire \us30/_0064_ ;
wire \us30/_0065_ ;
wire \us30/_0066_ ;
wire \us30/_0067_ ;
wire \us30/_0069_ ;
wire \us30/_0070_ ;
wire \us30/_0072_ ;
wire \us30/_0073_ ;
wire \us30/_0074_ ;
wire \us30/_0075_ ;
wire \us30/_0076_ ;
wire \us30/_0077_ ;
wire \us30/_0078_ ;
wire \us30/_0079_ ;
wire \us30/_0081_ ;
wire \us30/_0082_ ;
wire \us30/_0085_ ;
wire \us30/_0086_ ;
wire \us30/_0087_ ;
wire \us30/_0088_ ;
wire \us30/_0089_ ;
wire \us30/_0090_ ;
wire \us30/_0091_ ;
wire \us30/_0092_ ;
wire \us30/_0093_ ;
wire \us30/_0094_ ;
wire \us30/_0095_ ;
wire \us30/_0096_ ;
wire \us30/_0097_ ;
wire \us30/_0098_ ;
wire \us30/_0099_ ;
wire \us30/_0100_ ;
wire \us30/_0101_ ;
wire \us30/_0102_ ;
wire \us30/_0103_ ;
wire \us30/_0104_ ;
wire \us30/_0105_ ;
wire \us30/_0106_ ;
wire \us30/_0108_ ;
wire \us30/_0109_ ;
wire \us30/_0110_ ;
wire \us30/_0111_ ;
wire \us30/_0113_ ;
wire \us30/_0114_ ;
wire \us30/_0115_ ;
wire \us30/_0116_ ;
wire \us30/_0117_ ;
wire \us30/_0118_ ;
wire \us30/_0119_ ;
wire \us30/_0120_ ;
wire \us30/_0121_ ;
wire \us30/_0122_ ;
wire \us30/_0123_ ;
wire \us30/_0124_ ;
wire \us30/_0126_ ;
wire \us30/_0127_ ;
wire \us30/_0128_ ;
wire \us30/_0129_ ;
wire \us30/_0130_ ;
wire \us30/_0132_ ;
wire \us30/_0133_ ;
wire \us30/_0134_ ;
wire \us30/_0135_ ;
wire \us30/_0136_ ;
wire \us30/_0137_ ;
wire \us30/_0139_ ;
wire \us30/_0140_ ;
wire \us30/_0141_ ;
wire \us30/_0142_ ;
wire \us30/_0144_ ;
wire \us30/_0145_ ;
wire \us30/_0146_ ;
wire \us30/_0147_ ;
wire \us30/_0148_ ;
wire \us30/_0149_ ;
wire \us30/_0150_ ;
wire \us30/_0151_ ;
wire \us30/_0153_ ;
wire \us30/_0154_ ;
wire \us30/_0155_ ;
wire \us30/_0156_ ;
wire \us30/_0157_ ;
wire \us30/_0158_ ;
wire \us30/_0159_ ;
wire \us30/_0161_ ;
wire \us30/_0162_ ;
wire \us30/_0163_ ;
wire \us30/_0164_ ;
wire \us30/_0165_ ;
wire \us30/_0166_ ;
wire \us30/_0167_ ;
wire \us30/_0168_ ;
wire \us30/_0169_ ;
wire \us30/_0170_ ;
wire \us30/_0171_ ;
wire \us30/_0172_ ;
wire \us30/_0174_ ;
wire \us30/_0175_ ;
wire \us30/_0176_ ;
wire \us30/_0177_ ;
wire \us30/_0178_ ;
wire \us30/_0179_ ;
wire \us30/_0180_ ;
wire \us30/_0181_ ;
wire \us30/_0182_ ;
wire \us30/_0183_ ;
wire \us30/_0184_ ;
wire \us30/_0185_ ;
wire \us30/_0186_ ;
wire \us30/_0187_ ;
wire \us30/_0188_ ;
wire \us30/_0189_ ;
wire \us30/_0190_ ;
wire \us30/_0191_ ;
wire \us30/_0192_ ;
wire \us30/_0193_ ;
wire \us30/_0194_ ;
wire \us30/_0195_ ;
wire \us30/_0196_ ;
wire \us30/_0197_ ;
wire \us30/_0198_ ;
wire \us30/_0199_ ;
wire \us30/_0200_ ;
wire \us30/_0201_ ;
wire \us30/_0202_ ;
wire \us30/_0203_ ;
wire \us30/_0204_ ;
wire \us30/_0205_ ;
wire \us30/_0206_ ;
wire \us30/_0207_ ;
wire \us30/_0208_ ;
wire \us30/_0209_ ;
wire \us30/_0210_ ;
wire \us30/_0211_ ;
wire \us30/_0212_ ;
wire \us30/_0213_ ;
wire \us30/_0214_ ;
wire \us30/_0215_ ;
wire \us30/_0217_ ;
wire \us30/_0219_ ;
wire \us30/_0220_ ;
wire \us30/_0221_ ;
wire \us30/_0222_ ;
wire \us30/_0223_ ;
wire \us30/_0224_ ;
wire \us30/_0225_ ;
wire \us30/_0226_ ;
wire \us30/_0227_ ;
wire \us30/_0228_ ;
wire \us30/_0229_ ;
wire \us30/_0230_ ;
wire \us30/_0231_ ;
wire \us30/_0232_ ;
wire \us30/_0233_ ;
wire \us30/_0234_ ;
wire \us30/_0235_ ;
wire \us30/_0236_ ;
wire \us30/_0237_ ;
wire \us30/_0238_ ;
wire \us30/_0239_ ;
wire \us30/_0240_ ;
wire \us30/_0241_ ;
wire \us30/_0242_ ;
wire \us30/_0243_ ;
wire \us30/_0244_ ;
wire \us30/_0245_ ;
wire \us30/_0246_ ;
wire \us30/_0247_ ;
wire \us30/_0248_ ;
wire \us30/_0249_ ;
wire \us30/_0250_ ;
wire \us30/_0251_ ;
wire \us30/_0252_ ;
wire \us30/_0253_ ;
wire \us30/_0254_ ;
wire \us30/_0255_ ;
wire \us30/_0256_ ;
wire \us30/_0257_ ;
wire \us30/_0258_ ;
wire \us30/_0259_ ;
wire \us30/_0260_ ;
wire \us30/_0261_ ;
wire \us30/_0263_ ;
wire \us30/_0264_ ;
wire \us30/_0265_ ;
wire \us30/_0266_ ;
wire \us30/_0267_ ;
wire \us30/_0268_ ;
wire \us30/_0269_ ;
wire \us30/_0270_ ;
wire \us30/_0271_ ;
wire \us30/_0272_ ;
wire \us30/_0273_ ;
wire \us30/_0274_ ;
wire \us30/_0275_ ;
wire \us30/_0276_ ;
wire \us30/_0277_ ;
wire \us30/_0278_ ;
wire \us30/_0279_ ;
wire \us30/_0280_ ;
wire \us30/_0281_ ;
wire \us30/_0283_ ;
wire \us30/_0284_ ;
wire \us30/_0285_ ;
wire \us30/_0286_ ;
wire \us30/_0287_ ;
wire \us30/_0288_ ;
wire \us30/_0289_ ;
wire \us30/_0290_ ;
wire \us30/_0291_ ;
wire \us30/_0292_ ;
wire \us30/_0293_ ;
wire \us30/_0294_ ;
wire \us30/_0295_ ;
wire \us30/_0296_ ;
wire \us30/_0297_ ;
wire \us30/_0298_ ;
wire \us30/_0299_ ;
wire \us30/_0300_ ;
wire \us30/_0301_ ;
wire \us30/_0302_ ;
wire \us30/_0303_ ;
wire \us30/_0304_ ;
wire \us30/_0305_ ;
wire \us30/_0306_ ;
wire \us30/_0307_ ;
wire \us30/_0308_ ;
wire \us30/_0309_ ;
wire \us30/_0310_ ;
wire \us30/_0311_ ;
wire \us30/_0312_ ;
wire \us30/_0313_ ;
wire \us30/_0314_ ;
wire \us30/_0315_ ;
wire \us30/_0316_ ;
wire \us30/_0317_ ;
wire \us30/_0318_ ;
wire \us30/_0319_ ;
wire \us30/_0320_ ;
wire \us30/_0321_ ;
wire \us30/_0322_ ;
wire \us30/_0323_ ;
wire \us30/_0324_ ;
wire \us30/_0325_ ;
wire \us30/_0326_ ;
wire \us30/_0327_ ;
wire \us30/_0328_ ;
wire \us30/_0329_ ;
wire \us30/_0330_ ;
wire \us30/_0331_ ;
wire \us30/_0332_ ;
wire \us30/_0333_ ;
wire \us30/_0334_ ;
wire \us30/_0335_ ;
wire \us30/_0337_ ;
wire \us30/_0338_ ;
wire \us30/_0339_ ;
wire \us30/_0340_ ;
wire \us30/_0341_ ;
wire \us30/_0342_ ;
wire \us30/_0343_ ;
wire \us30/_0344_ ;
wire \us30/_0345_ ;
wire \us30/_0347_ ;
wire \us30/_0348_ ;
wire \us30/_0349_ ;
wire \us30/_0350_ ;
wire \us30/_0351_ ;
wire \us30/_0352_ ;
wire \us30/_0353_ ;
wire \us30/_0354_ ;
wire \us30/_0355_ ;
wire \us30/_0356_ ;
wire \us30/_0357_ ;
wire \us30/_0358_ ;
wire \us30/_0359_ ;
wire \us30/_0360_ ;
wire \us30/_0361_ ;
wire \us30/_0362_ ;
wire \us30/_0363_ ;
wire \us30/_0365_ ;
wire \us30/_0366_ ;
wire \us30/_0367_ ;
wire \us30/_0368_ ;
wire \us30/_0370_ ;
wire \us30/_0371_ ;
wire \us30/_0372_ ;
wire \us30/_0373_ ;
wire \us30/_0374_ ;
wire \us30/_0375_ ;
wire \us30/_0376_ ;
wire \us30/_0377_ ;
wire \us30/_0378_ ;
wire \us30/_0379_ ;
wire \us30/_0380_ ;
wire \us30/_0381_ ;
wire \us30/_0382_ ;
wire \us30/_0383_ ;
wire \us30/_0384_ ;
wire \us30/_0385_ ;
wire \us30/_0386_ ;
wire \us30/_0387_ ;
wire \us30/_0388_ ;
wire \us30/_0389_ ;
wire \us30/_0390_ ;
wire \us30/_0391_ ;
wire \us30/_0392_ ;
wire \us30/_0393_ ;
wire \us30/_0394_ ;
wire \us30/_0395_ ;
wire \us30/_0396_ ;
wire \us30/_0397_ ;
wire \us30/_0398_ ;
wire \us30/_0399_ ;
wire \us30/_0400_ ;
wire \us30/_0401_ ;
wire \us30/_0402_ ;
wire \us30/_0403_ ;
wire \us30/_0404_ ;
wire \us30/_0405_ ;
wire \us30/_0406_ ;
wire \us30/_0407_ ;
wire \us30/_0408_ ;
wire \us30/_0409_ ;
wire \us30/_0410_ ;
wire \us30/_0411_ ;
wire \us30/_0412_ ;
wire \us30/_0413_ ;
wire \us30/_0414_ ;
wire \us30/_0415_ ;
wire \us30/_0416_ ;
wire \us30/_0417_ ;
wire \us30/_0418_ ;
wire \us30/_0419_ ;
wire \us30/_0420_ ;
wire \us30/_0421_ ;
wire \us30/_0422_ ;
wire \us30/_0424_ ;
wire \us30/_0425_ ;
wire \us30/_0426_ ;
wire \us30/_0427_ ;
wire \us30/_0428_ ;
wire \us30/_0429_ ;
wire \us30/_0430_ ;
wire \us30/_0431_ ;
wire \us30/_0432_ ;
wire \us30/_0433_ ;
wire \us30/_0434_ ;
wire \us30/_0435_ ;
wire \us30/_0436_ ;
wire \us30/_0437_ ;
wire \us30/_0438_ ;
wire \us30/_0439_ ;
wire \us30/_0440_ ;
wire \us30/_0441_ ;
wire \us30/_0442_ ;
wire \us30/_0443_ ;
wire \us30/_0444_ ;
wire \us30/_0446_ ;
wire \us30/_0447_ ;
wire \us30/_0448_ ;
wire \us30/_0449_ ;
wire \us30/_0450_ ;
wire \us30/_0451_ ;
wire \us30/_0452_ ;
wire \us30/_0453_ ;
wire \us30/_0454_ ;
wire \us30/_0455_ ;
wire \us30/_0457_ ;
wire \us30/_0458_ ;
wire \us30/_0459_ ;
wire \us30/_0460_ ;
wire \us30/_0461_ ;
wire \us30/_0462_ ;
wire \us30/_0463_ ;
wire \us30/_0464_ ;
wire \us30/_0465_ ;
wire \us30/_0466_ ;
wire \us30/_0467_ ;
wire \us30/_0468_ ;
wire \us30/_0469_ ;
wire \us30/_0470_ ;
wire \us30/_0471_ ;
wire \us30/_0472_ ;
wire \us30/_0473_ ;
wire \us30/_0474_ ;
wire \us30/_0475_ ;
wire \us30/_0476_ ;
wire \us30/_0477_ ;
wire \us30/_0478_ ;
wire \us30/_0479_ ;
wire \us30/_0480_ ;
wire \us30/_0481_ ;
wire \us30/_0482_ ;
wire \us30/_0483_ ;
wire \us30/_0484_ ;
wire \us30/_0485_ ;
wire \us30/_0486_ ;
wire \us30/_0487_ ;
wire \us30/_0488_ ;
wire \us30/_0490_ ;
wire \us30/_0491_ ;
wire \us30/_0492_ ;
wire \us30/_0493_ ;
wire \us30/_0494_ ;
wire \us30/_0495_ ;
wire \us30/_0496_ ;
wire \us30/_0497_ ;
wire \us30/_0498_ ;
wire \us30/_0499_ ;
wire \us30/_0500_ ;
wire \us30/_0501_ ;
wire \us30/_0502_ ;
wire \us30/_0503_ ;
wire \us30/_0504_ ;
wire \us30/_0505_ ;
wire \us30/_0506_ ;
wire \us30/_0507_ ;
wire \us30/_0508_ ;
wire \us30/_0509_ ;
wire \us30/_0510_ ;
wire \us30/_0511_ ;
wire \us30/_0512_ ;
wire \us30/_0513_ ;
wire \us30/_0514_ ;
wire \us30/_0515_ ;
wire \us30/_0516_ ;
wire \us30/_0517_ ;
wire \us30/_0518_ ;
wire \us30/_0519_ ;
wire \us30/_0520_ ;
wire \us30/_0521_ ;
wire \us30/_0522_ ;
wire \us30/_0523_ ;
wire \us30/_0524_ ;
wire \us30/_0525_ ;
wire \us30/_0526_ ;
wire \us30/_0527_ ;
wire \us30/_0528_ ;
wire \us30/_0529_ ;
wire \us30/_0530_ ;
wire \us30/_0531_ ;
wire \us30/_0532_ ;
wire \us30/_0533_ ;
wire \us30/_0534_ ;
wire \us30/_0535_ ;
wire \us30/_0536_ ;
wire \us30/_0537_ ;
wire \us30/_0538_ ;
wire \us30/_0539_ ;
wire \us30/_0540_ ;
wire \us30/_0541_ ;
wire \us30/_0542_ ;
wire \us30/_0544_ ;
wire \us30/_0545_ ;
wire \us30/_0546_ ;
wire \us30/_0547_ ;
wire \us30/_0548_ ;
wire \us30/_0549_ ;
wire \us30/_0550_ ;
wire \us30/_0551_ ;
wire \us30/_0552_ ;
wire \us30/_0553_ ;
wire \us30/_0554_ ;
wire \us30/_0555_ ;
wire \us30/_0556_ ;
wire \us30/_0557_ ;
wire \us30/_0558_ ;
wire \us30/_0559_ ;
wire \us30/_0560_ ;
wire \us30/_0561_ ;
wire \us30/_0562_ ;
wire \us30/_0563_ ;
wire \us30/_0565_ ;
wire \us30/_0566_ ;
wire \us30/_0567_ ;
wire \us30/_0568_ ;
wire \us30/_0569_ ;
wire \us30/_0570_ ;
wire \us30/_0571_ ;
wire \us30/_0572_ ;
wire \us30/_0573_ ;
wire \us30/_0574_ ;
wire \us30/_0575_ ;
wire \us30/_0576_ ;
wire \us30/_0577_ ;
wire \us30/_0578_ ;
wire \us30/_0579_ ;
wire \us30/_0580_ ;
wire \us30/_0581_ ;
wire \us30/_0582_ ;
wire \us30/_0583_ ;
wire \us30/_0584_ ;
wire \us30/_0585_ ;
wire \us30/_0586_ ;
wire \us30/_0587_ ;
wire \us30/_0588_ ;
wire \us30/_0589_ ;
wire \us30/_0590_ ;
wire \us30/_0591_ ;
wire \us30/_0592_ ;
wire \us30/_0593_ ;
wire \us30/_0594_ ;
wire \us30/_0595_ ;
wire \us30/_0596_ ;
wire \us30/_0598_ ;
wire \us30/_0599_ ;
wire \us30/_0600_ ;
wire \us30/_0601_ ;
wire \us30/_0602_ ;
wire \us30/_0603_ ;
wire \us30/_0604_ ;
wire \us30/_0605_ ;
wire \us30/_0606_ ;
wire \us30/_0607_ ;
wire \us30/_0608_ ;
wire \us30/_0609_ ;
wire \us30/_0610_ ;
wire \us30/_0611_ ;
wire \us30/_0612_ ;
wire \us30/_0613_ ;
wire \us30/_0614_ ;
wire \us30/_0615_ ;
wire \us30/_0616_ ;
wire \us30/_0617_ ;
wire \us30/_0618_ ;
wire \us30/_0619_ ;
wire \us30/_0620_ ;
wire \us30/_0621_ ;
wire \us30/_0622_ ;
wire \us30/_0623_ ;
wire \us30/_0624_ ;
wire \us30/_0625_ ;
wire \us30/_0626_ ;
wire \us30/_0627_ ;
wire \us30/_0628_ ;
wire \us30/_0629_ ;
wire \us30/_0630_ ;
wire \us30/_0631_ ;
wire \us30/_0632_ ;
wire \us30/_0633_ ;
wire \us30/_0634_ ;
wire \us30/_0635_ ;
wire \us30/_0636_ ;
wire \us30/_0637_ ;
wire \us30/_0638_ ;
wire \us30/_0639_ ;
wire \us30/_0640_ ;
wire \us30/_0641_ ;
wire \us30/_0642_ ;
wire \us30/_0643_ ;
wire \us30/_0644_ ;
wire \us30/_0645_ ;
wire \us30/_0646_ ;
wire \us30/_0647_ ;
wire \us30/_0648_ ;
wire \us30/_0649_ ;
wire \us30/_0650_ ;
wire \us30/_0652_ ;
wire \us30/_0653_ ;
wire \us30/_0654_ ;
wire \us30/_0655_ ;
wire \us30/_0656_ ;
wire \us30/_0657_ ;
wire \us30/_0658_ ;
wire \us30/_0659_ ;
wire \us30/_0660_ ;
wire \us30/_0661_ ;
wire \us30/_0662_ ;
wire \us30/_0663_ ;
wire \us30/_0664_ ;
wire \us30/_0665_ ;
wire \us30/_0666_ ;
wire \us30/_0667_ ;
wire \us30/_0668_ ;
wire \us30/_0669_ ;
wire \us30/_0670_ ;
wire \us30/_0671_ ;
wire \us30/_0673_ ;
wire \us30/_0674_ ;
wire \us30/_0675_ ;
wire \us30/_0676_ ;
wire \us30/_0677_ ;
wire \us30/_0678_ ;
wire \us30/_0679_ ;
wire \us30/_0680_ ;
wire \us30/_0681_ ;
wire \us30/_0682_ ;
wire \us30/_0683_ ;
wire \us30/_0684_ ;
wire \us30/_0685_ ;
wire \us30/_0686_ ;
wire \us30/_0687_ ;
wire \us30/_0688_ ;
wire \us30/_0689_ ;
wire \us30/_0690_ ;
wire \us30/_0691_ ;
wire \us30/_0692_ ;
wire \us30/_0693_ ;
wire \us30/_0694_ ;
wire \us30/_0695_ ;
wire \us30/_0696_ ;
wire \us30/_0697_ ;
wire \us30/_0698_ ;
wire \us30/_0699_ ;
wire \us30/_0700_ ;
wire \us30/_0701_ ;
wire \us30/_0702_ ;
wire \us30/_0703_ ;
wire \us30/_0704_ ;
wire \us30/_0705_ ;
wire \us30/_0706_ ;
wire \us30/_0707_ ;
wire \us30/_0708_ ;
wire \us30/_0709_ ;
wire \us30/_0710_ ;
wire \us30/_0711_ ;
wire \us30/_0712_ ;
wire \us30/_0713_ ;
wire \us30/_0714_ ;
wire \us30/_0715_ ;
wire \us30/_0717_ ;
wire \us30/_0718_ ;
wire \us30/_0719_ ;
wire \us30/_0720_ ;
wire \us30/_0721_ ;
wire \us30/_0722_ ;
wire \us30/_0723_ ;
wire \us30/_0724_ ;
wire \us30/_0725_ ;
wire \us30/_0726_ ;
wire \us30/_0727_ ;
wire \us30/_0728_ ;
wire \us30/_0729_ ;
wire \us30/_0730_ ;
wire \us30/_0731_ ;
wire \us30/_0733_ ;
wire \us30/_0734_ ;
wire \us30/_0735_ ;
wire \us30/_0736_ ;
wire \us30/_0738_ ;
wire \us30/_0739_ ;
wire \us30/_0740_ ;
wire \us30/_0741_ ;
wire \us30/_0742_ ;
wire \us30/_0744_ ;
wire \us30/_0745_ ;
wire \us30/_0746_ ;
wire \us30/_0748_ ;
wire \us30/_0749_ ;
wire \us30/_0750_ ;
wire \us30/_0752_ ;
wire \us31/_0008_ ;
wire \us31/_0009_ ;
wire \us31/_0010_ ;
wire \us31/_0011_ ;
wire \us31/_0012_ ;
wire \us31/_0013_ ;
wire \us31/_0014_ ;
wire \us31/_0015_ ;
wire \us31/_0016_ ;
wire \us31/_0017_ ;
wire \us31/_0019_ ;
wire \us31/_0020_ ;
wire \us31/_0022_ ;
wire \us31/_0024_ ;
wire \us31/_0025_ ;
wire \us31/_0026_ ;
wire \us31/_0027_ ;
wire \us31/_0030_ ;
wire \us31/_0032_ ;
wire \us31/_0033_ ;
wire \us31/_0034_ ;
wire \us31/_0035_ ;
wire \us31/_0037_ ;
wire \us31/_0038_ ;
wire \us31/_0039_ ;
wire \us31/_0040_ ;
wire \us31/_0041_ ;
wire \us31/_0042_ ;
wire \us31/_0043_ ;
wire \us31/_0045_ ;
wire \us31/_0046_ ;
wire \us31/_0047_ ;
wire \us31/_0049_ ;
wire \us31/_0050_ ;
wire \us31/_0051_ ;
wire \us31/_0052_ ;
wire \us31/_0053_ ;
wire \us31/_0054_ ;
wire \us31/_0057_ ;
wire \us31/_0058_ ;
wire \us31/_0060_ ;
wire \us31/_0061_ ;
wire \us31/_0062_ ;
wire \us31/_0064_ ;
wire \us31/_0065_ ;
wire \us31/_0066_ ;
wire \us31/_0067_ ;
wire \us31/_0069_ ;
wire \us31/_0070_ ;
wire \us31/_0072_ ;
wire \us31/_0073_ ;
wire \us31/_0074_ ;
wire \us31/_0075_ ;
wire \us31/_0076_ ;
wire \us31/_0077_ ;
wire \us31/_0078_ ;
wire \us31/_0079_ ;
wire \us31/_0081_ ;
wire \us31/_0082_ ;
wire \us31/_0084_ ;
wire \us31/_0085_ ;
wire \us31/_0086_ ;
wire \us31/_0087_ ;
wire \us31/_0088_ ;
wire \us31/_0089_ ;
wire \us31/_0090_ ;
wire \us31/_0091_ ;
wire \us31/_0092_ ;
wire \us31/_0093_ ;
wire \us31/_0094_ ;
wire \us31/_0095_ ;
wire \us31/_0096_ ;
wire \us31/_0097_ ;
wire \us31/_0098_ ;
wire \us31/_0099_ ;
wire \us31/_0100_ ;
wire \us31/_0101_ ;
wire \us31/_0102_ ;
wire \us31/_0103_ ;
wire \us31/_0104_ ;
wire \us31/_0105_ ;
wire \us31/_0106_ ;
wire \us31/_0108_ ;
wire \us31/_0109_ ;
wire \us31/_0110_ ;
wire \us31/_0111_ ;
wire \us31/_0113_ ;
wire \us31/_0114_ ;
wire \us31/_0115_ ;
wire \us31/_0116_ ;
wire \us31/_0117_ ;
wire \us31/_0118_ ;
wire \us31/_0119_ ;
wire \us31/_0120_ ;
wire \us31/_0121_ ;
wire \us31/_0122_ ;
wire \us31/_0123_ ;
wire \us31/_0124_ ;
wire \us31/_0126_ ;
wire \us31/_0127_ ;
wire \us31/_0128_ ;
wire \us31/_0129_ ;
wire \us31/_0130_ ;
wire \us31/_0132_ ;
wire \us31/_0133_ ;
wire \us31/_0134_ ;
wire \us31/_0135_ ;
wire \us31/_0136_ ;
wire \us31/_0137_ ;
wire \us31/_0139_ ;
wire \us31/_0140_ ;
wire \us31/_0141_ ;
wire \us31/_0142_ ;
wire \us31/_0144_ ;
wire \us31/_0145_ ;
wire \us31/_0146_ ;
wire \us31/_0147_ ;
wire \us31/_0148_ ;
wire \us31/_0149_ ;
wire \us31/_0150_ ;
wire \us31/_0151_ ;
wire \us31/_0153_ ;
wire \us31/_0154_ ;
wire \us31/_0155_ ;
wire \us31/_0156_ ;
wire \us31/_0157_ ;
wire \us31/_0158_ ;
wire \us31/_0159_ ;
wire \us31/_0161_ ;
wire \us31/_0162_ ;
wire \us31/_0163_ ;
wire \us31/_0164_ ;
wire \us31/_0165_ ;
wire \us31/_0166_ ;
wire \us31/_0167_ ;
wire \us31/_0168_ ;
wire \us31/_0169_ ;
wire \us31/_0170_ ;
wire \us31/_0171_ ;
wire \us31/_0172_ ;
wire \us31/_0174_ ;
wire \us31/_0175_ ;
wire \us31/_0176_ ;
wire \us31/_0177_ ;
wire \us31/_0178_ ;
wire \us31/_0179_ ;
wire \us31/_0180_ ;
wire \us31/_0181_ ;
wire \us31/_0182_ ;
wire \us31/_0183_ ;
wire \us31/_0184_ ;
wire \us31/_0185_ ;
wire \us31/_0186_ ;
wire \us31/_0187_ ;
wire \us31/_0188_ ;
wire \us31/_0189_ ;
wire \us31/_0190_ ;
wire \us31/_0191_ ;
wire \us31/_0192_ ;
wire \us31/_0193_ ;
wire \us31/_0194_ ;
wire \us31/_0195_ ;
wire \us31/_0196_ ;
wire \us31/_0197_ ;
wire \us31/_0198_ ;
wire \us31/_0199_ ;
wire \us31/_0200_ ;
wire \us31/_0201_ ;
wire \us31/_0202_ ;
wire \us31/_0203_ ;
wire \us31/_0204_ ;
wire \us31/_0205_ ;
wire \us31/_0206_ ;
wire \us31/_0207_ ;
wire \us31/_0208_ ;
wire \us31/_0209_ ;
wire \us31/_0210_ ;
wire \us31/_0211_ ;
wire \us31/_0212_ ;
wire \us31/_0213_ ;
wire \us31/_0214_ ;
wire \us31/_0215_ ;
wire \us31/_0217_ ;
wire \us31/_0218_ ;
wire \us31/_0219_ ;
wire \us31/_0220_ ;
wire \us31/_0221_ ;
wire \us31/_0222_ ;
wire \us31/_0223_ ;
wire \us31/_0224_ ;
wire \us31/_0225_ ;
wire \us31/_0226_ ;
wire \us31/_0227_ ;
wire \us31/_0228_ ;
wire \us31/_0229_ ;
wire \us31/_0230_ ;
wire \us31/_0231_ ;
wire \us31/_0232_ ;
wire \us31/_0233_ ;
wire \us31/_0234_ ;
wire \us31/_0235_ ;
wire \us31/_0236_ ;
wire \us31/_0237_ ;
wire \us31/_0238_ ;
wire \us31/_0239_ ;
wire \us31/_0240_ ;
wire \us31/_0241_ ;
wire \us31/_0242_ ;
wire \us31/_0243_ ;
wire \us31/_0244_ ;
wire \us31/_0245_ ;
wire \us31/_0246_ ;
wire \us31/_0247_ ;
wire \us31/_0248_ ;
wire \us31/_0249_ ;
wire \us31/_0250_ ;
wire \us31/_0251_ ;
wire \us31/_0252_ ;
wire \us31/_0253_ ;
wire \us31/_0254_ ;
wire \us31/_0255_ ;
wire \us31/_0256_ ;
wire \us31/_0257_ ;
wire \us31/_0258_ ;
wire \us31/_0259_ ;
wire \us31/_0260_ ;
wire \us31/_0261_ ;
wire \us31/_0263_ ;
wire \us31/_0264_ ;
wire \us31/_0265_ ;
wire \us31/_0266_ ;
wire \us31/_0267_ ;
wire \us31/_0268_ ;
wire \us31/_0269_ ;
wire \us31/_0270_ ;
wire \us31/_0271_ ;
wire \us31/_0272_ ;
wire \us31/_0273_ ;
wire \us31/_0274_ ;
wire \us31/_0275_ ;
wire \us31/_0276_ ;
wire \us31/_0277_ ;
wire \us31/_0278_ ;
wire \us31/_0279_ ;
wire \us31/_0281_ ;
wire \us31/_0283_ ;
wire \us31/_0284_ ;
wire \us31/_0285_ ;
wire \us31/_0286_ ;
wire \us31/_0287_ ;
wire \us31/_0288_ ;
wire \us31/_0289_ ;
wire \us31/_0290_ ;
wire \us31/_0291_ ;
wire \us31/_0292_ ;
wire \us31/_0293_ ;
wire \us31/_0294_ ;
wire \us31/_0295_ ;
wire \us31/_0296_ ;
wire \us31/_0297_ ;
wire \us31/_0298_ ;
wire \us31/_0299_ ;
wire \us31/_0300_ ;
wire \us31/_0301_ ;
wire \us31/_0302_ ;
wire \us31/_0303_ ;
wire \us31/_0304_ ;
wire \us31/_0305_ ;
wire \us31/_0306_ ;
wire \us31/_0307_ ;
wire \us31/_0308_ ;
wire \us31/_0309_ ;
wire \us31/_0310_ ;
wire \us31/_0311_ ;
wire \us31/_0312_ ;
wire \us31/_0313_ ;
wire \us31/_0314_ ;
wire \us31/_0315_ ;
wire \us31/_0316_ ;
wire \us31/_0317_ ;
wire \us31/_0318_ ;
wire \us31/_0319_ ;
wire \us31/_0320_ ;
wire \us31/_0321_ ;
wire \us31/_0322_ ;
wire \us31/_0323_ ;
wire \us31/_0324_ ;
wire \us31/_0325_ ;
wire \us31/_0326_ ;
wire \us31/_0327_ ;
wire \us31/_0328_ ;
wire \us31/_0329_ ;
wire \us31/_0330_ ;
wire \us31/_0331_ ;
wire \us31/_0332_ ;
wire \us31/_0333_ ;
wire \us31/_0334_ ;
wire \us31/_0335_ ;
wire \us31/_0337_ ;
wire \us31/_0338_ ;
wire \us31/_0339_ ;
wire \us31/_0340_ ;
wire \us31/_0341_ ;
wire \us31/_0342_ ;
wire \us31/_0343_ ;
wire \us31/_0344_ ;
wire \us31/_0345_ ;
wire \us31/_0347_ ;
wire \us31/_0348_ ;
wire \us31/_0349_ ;
wire \us31/_0350_ ;
wire \us31/_0351_ ;
wire \us31/_0352_ ;
wire \us31/_0353_ ;
wire \us31/_0354_ ;
wire \us31/_0355_ ;
wire \us31/_0356_ ;
wire \us31/_0357_ ;
wire \us31/_0358_ ;
wire \us31/_0359_ ;
wire \us31/_0360_ ;
wire \us31/_0361_ ;
wire \us31/_0362_ ;
wire \us31/_0363_ ;
wire \us31/_0365_ ;
wire \us31/_0366_ ;
wire \us31/_0367_ ;
wire \us31/_0368_ ;
wire \us31/_0370_ ;
wire \us31/_0371_ ;
wire \us31/_0372_ ;
wire \us31/_0373_ ;
wire \us31/_0374_ ;
wire \us31/_0375_ ;
wire \us31/_0376_ ;
wire \us31/_0377_ ;
wire \us31/_0378_ ;
wire \us31/_0379_ ;
wire \us31/_0380_ ;
wire \us31/_0381_ ;
wire \us31/_0382_ ;
wire \us31/_0383_ ;
wire \us31/_0384_ ;
wire \us31/_0385_ ;
wire \us31/_0386_ ;
wire \us31/_0387_ ;
wire \us31/_0388_ ;
wire \us31/_0389_ ;
wire \us31/_0390_ ;
wire \us31/_0391_ ;
wire \us31/_0392_ ;
wire \us31/_0393_ ;
wire \us31/_0394_ ;
wire \us31/_0395_ ;
wire \us31/_0396_ ;
wire \us31/_0397_ ;
wire \us31/_0398_ ;
wire \us31/_0399_ ;
wire \us31/_0400_ ;
wire \us31/_0401_ ;
wire \us31/_0402_ ;
wire \us31/_0403_ ;
wire \us31/_0404_ ;
wire \us31/_0405_ ;
wire \us31/_0406_ ;
wire \us31/_0407_ ;
wire \us31/_0408_ ;
wire \us31/_0409_ ;
wire \us31/_0410_ ;
wire \us31/_0411_ ;
wire \us31/_0412_ ;
wire \us31/_0413_ ;
wire \us31/_0414_ ;
wire \us31/_0415_ ;
wire \us31/_0416_ ;
wire \us31/_0417_ ;
wire \us31/_0418_ ;
wire \us31/_0419_ ;
wire \us31/_0420_ ;
wire \us31/_0421_ ;
wire \us31/_0422_ ;
wire \us31/_0423_ ;
wire \us31/_0424_ ;
wire \us31/_0425_ ;
wire \us31/_0426_ ;
wire \us31/_0427_ ;
wire \us31/_0428_ ;
wire \us31/_0429_ ;
wire \us31/_0430_ ;
wire \us31/_0431_ ;
wire \us31/_0432_ ;
wire \us31/_0433_ ;
wire \us31/_0434_ ;
wire \us31/_0435_ ;
wire \us31/_0436_ ;
wire \us31/_0437_ ;
wire \us31/_0438_ ;
wire \us31/_0439_ ;
wire \us31/_0440_ ;
wire \us31/_0441_ ;
wire \us31/_0442_ ;
wire \us31/_0443_ ;
wire \us31/_0444_ ;
wire \us31/_0446_ ;
wire \us31/_0447_ ;
wire \us31/_0448_ ;
wire \us31/_0449_ ;
wire \us31/_0450_ ;
wire \us31/_0451_ ;
wire \us31/_0452_ ;
wire \us31/_0453_ ;
wire \us31/_0454_ ;
wire \us31/_0455_ ;
wire \us31/_0457_ ;
wire \us31/_0458_ ;
wire \us31/_0459_ ;
wire \us31/_0460_ ;
wire \us31/_0461_ ;
wire \us31/_0462_ ;
wire \us31/_0463_ ;
wire \us31/_0464_ ;
wire \us31/_0465_ ;
wire \us31/_0466_ ;
wire \us31/_0467_ ;
wire \us31/_0468_ ;
wire \us31/_0469_ ;
wire \us31/_0470_ ;
wire \us31/_0471_ ;
wire \us31/_0472_ ;
wire \us31/_0473_ ;
wire \us31/_0474_ ;
wire \us31/_0475_ ;
wire \us31/_0476_ ;
wire \us31/_0477_ ;
wire \us31/_0478_ ;
wire \us31/_0479_ ;
wire \us31/_0480_ ;
wire \us31/_0481_ ;
wire \us31/_0482_ ;
wire \us31/_0483_ ;
wire \us31/_0484_ ;
wire \us31/_0485_ ;
wire \us31/_0486_ ;
wire \us31/_0487_ ;
wire \us31/_0488_ ;
wire \us31/_0490_ ;
wire \us31/_0491_ ;
wire \us31/_0492_ ;
wire \us31/_0493_ ;
wire \us31/_0494_ ;
wire \us31/_0495_ ;
wire \us31/_0496_ ;
wire \us31/_0497_ ;
wire \us31/_0498_ ;
wire \us31/_0500_ ;
wire \us31/_0501_ ;
wire \us31/_0502_ ;
wire \us31/_0503_ ;
wire \us31/_0504_ ;
wire \us31/_0505_ ;
wire \us31/_0506_ ;
wire \us31/_0507_ ;
wire \us31/_0508_ ;
wire \us31/_0509_ ;
wire \us31/_0510_ ;
wire \us31/_0511_ ;
wire \us31/_0512_ ;
wire \us31/_0513_ ;
wire \us31/_0514_ ;
wire \us31/_0515_ ;
wire \us31/_0516_ ;
wire \us31/_0517_ ;
wire \us31/_0518_ ;
wire \us31/_0519_ ;
wire \us31/_0520_ ;
wire \us31/_0521_ ;
wire \us31/_0522_ ;
wire \us31/_0523_ ;
wire \us31/_0524_ ;
wire \us31/_0525_ ;
wire \us31/_0526_ ;
wire \us31/_0527_ ;
wire \us31/_0528_ ;
wire \us31/_0529_ ;
wire \us31/_0530_ ;
wire \us31/_0531_ ;
wire \us31/_0532_ ;
wire \us31/_0533_ ;
wire \us31/_0534_ ;
wire \us31/_0535_ ;
wire \us31/_0536_ ;
wire \us31/_0537_ ;
wire \us31/_0538_ ;
wire \us31/_0539_ ;
wire \us31/_0540_ ;
wire \us31/_0541_ ;
wire \us31/_0542_ ;
wire \us31/_0543_ ;
wire \us31/_0544_ ;
wire \us31/_0545_ ;
wire \us31/_0546_ ;
wire \us31/_0547_ ;
wire \us31/_0548_ ;
wire \us31/_0549_ ;
wire \us31/_0550_ ;
wire \us31/_0551_ ;
wire \us31/_0552_ ;
wire \us31/_0553_ ;
wire \us31/_0554_ ;
wire \us31/_0555_ ;
wire \us31/_0556_ ;
wire \us31/_0557_ ;
wire \us31/_0558_ ;
wire \us31/_0559_ ;
wire \us31/_0560_ ;
wire \us31/_0561_ ;
wire \us31/_0562_ ;
wire \us31/_0563_ ;
wire \us31/_0565_ ;
wire \us31/_0566_ ;
wire \us31/_0567_ ;
wire \us31/_0568_ ;
wire \us31/_0569_ ;
wire \us31/_0570_ ;
wire \us31/_0571_ ;
wire \us31/_0572_ ;
wire \us31/_0573_ ;
wire \us31/_0574_ ;
wire \us31/_0575_ ;
wire \us31/_0576_ ;
wire \us31/_0577_ ;
wire \us31/_0578_ ;
wire \us31/_0579_ ;
wire \us31/_0580_ ;
wire \us31/_0581_ ;
wire \us31/_0582_ ;
wire \us31/_0583_ ;
wire \us31/_0584_ ;
wire \us31/_0585_ ;
wire \us31/_0586_ ;
wire \us31/_0587_ ;
wire \us31/_0588_ ;
wire \us31/_0589_ ;
wire \us31/_0590_ ;
wire \us31/_0591_ ;
wire \us31/_0592_ ;
wire \us31/_0593_ ;
wire \us31/_0594_ ;
wire \us31/_0595_ ;
wire \us31/_0596_ ;
wire \us31/_0598_ ;
wire \us31/_0599_ ;
wire \us31/_0600_ ;
wire \us31/_0601_ ;
wire \us31/_0602_ ;
wire \us31/_0603_ ;
wire \us31/_0604_ ;
wire \us31/_0605_ ;
wire \us31/_0606_ ;
wire \us31/_0607_ ;
wire \us31/_0608_ ;
wire \us31/_0609_ ;
wire \us31/_0610_ ;
wire \us31/_0611_ ;
wire \us31/_0612_ ;
wire \us31/_0613_ ;
wire \us31/_0614_ ;
wire \us31/_0615_ ;
wire \us31/_0616_ ;
wire \us31/_0617_ ;
wire \us31/_0618_ ;
wire \us31/_0619_ ;
wire \us31/_0620_ ;
wire \us31/_0621_ ;
wire \us31/_0622_ ;
wire \us31/_0623_ ;
wire \us31/_0624_ ;
wire \us31/_0625_ ;
wire \us31/_0626_ ;
wire \us31/_0627_ ;
wire \us31/_0628_ ;
wire \us31/_0629_ ;
wire \us31/_0630_ ;
wire \us31/_0631_ ;
wire \us31/_0632_ ;
wire \us31/_0633_ ;
wire \us31/_0634_ ;
wire \us31/_0635_ ;
wire \us31/_0636_ ;
wire \us31/_0637_ ;
wire \us31/_0638_ ;
wire \us31/_0639_ ;
wire \us31/_0640_ ;
wire \us31/_0641_ ;
wire \us31/_0642_ ;
wire \us31/_0643_ ;
wire \us31/_0644_ ;
wire \us31/_0645_ ;
wire \us31/_0646_ ;
wire \us31/_0647_ ;
wire \us31/_0648_ ;
wire \us31/_0649_ ;
wire \us31/_0650_ ;
wire \us31/_0652_ ;
wire \us31/_0653_ ;
wire \us31/_0654_ ;
wire \us31/_0655_ ;
wire \us31/_0656_ ;
wire \us31/_0657_ ;
wire \us31/_0658_ ;
wire \us31/_0659_ ;
wire \us31/_0660_ ;
wire \us31/_0661_ ;
wire \us31/_0662_ ;
wire \us31/_0663_ ;
wire \us31/_0664_ ;
wire \us31/_0665_ ;
wire \us31/_0666_ ;
wire \us31/_0667_ ;
wire \us31/_0668_ ;
wire \us31/_0669_ ;
wire \us31/_0670_ ;
wire \us31/_0671_ ;
wire \us31/_0673_ ;
wire \us31/_0674_ ;
wire \us31/_0675_ ;
wire \us31/_0676_ ;
wire \us31/_0677_ ;
wire \us31/_0678_ ;
wire \us31/_0679_ ;
wire \us31/_0680_ ;
wire \us31/_0681_ ;
wire \us31/_0682_ ;
wire \us31/_0683_ ;
wire \us31/_0684_ ;
wire \us31/_0685_ ;
wire \us31/_0686_ ;
wire \us31/_0687_ ;
wire \us31/_0688_ ;
wire \us31/_0689_ ;
wire \us31/_0690_ ;
wire \us31/_0691_ ;
wire \us31/_0692_ ;
wire \us31/_0693_ ;
wire \us31/_0694_ ;
wire \us31/_0695_ ;
wire \us31/_0696_ ;
wire \us31/_0697_ ;
wire \us31/_0698_ ;
wire \us31/_0699_ ;
wire \us31/_0700_ ;
wire \us31/_0701_ ;
wire \us31/_0702_ ;
wire \us31/_0703_ ;
wire \us31/_0704_ ;
wire \us31/_0705_ ;
wire \us31/_0706_ ;
wire \us31/_0707_ ;
wire \us31/_0708_ ;
wire \us31/_0709_ ;
wire \us31/_0710_ ;
wire \us31/_0711_ ;
wire \us31/_0712_ ;
wire \us31/_0713_ ;
wire \us31/_0714_ ;
wire \us31/_0715_ ;
wire \us31/_0717_ ;
wire \us31/_0718_ ;
wire \us31/_0719_ ;
wire \us31/_0720_ ;
wire \us31/_0721_ ;
wire \us31/_0722_ ;
wire \us31/_0723_ ;
wire \us31/_0724_ ;
wire \us31/_0725_ ;
wire \us31/_0726_ ;
wire \us31/_0727_ ;
wire \us31/_0728_ ;
wire \us31/_0729_ ;
wire \us31/_0730_ ;
wire \us31/_0731_ ;
wire \us31/_0733_ ;
wire \us31/_0734_ ;
wire \us31/_0735_ ;
wire \us31/_0736_ ;
wire \us31/_0738_ ;
wire \us31/_0739_ ;
wire \us31/_0740_ ;
wire \us31/_0741_ ;
wire \us31/_0742_ ;
wire \us31/_0744_ ;
wire \us31/_0745_ ;
wire \us31/_0746_ ;
wire \us31/_0748_ ;
wire \us31/_0749_ ;
wire \us31/_0750_ ;
wire \us31/_0752_ ;
wire \us32/_0008_ ;
wire \us32/_0009_ ;
wire \us32/_0010_ ;
wire \us32/_0011_ ;
wire \us32/_0012_ ;
wire \us32/_0013_ ;
wire \us32/_0014_ ;
wire \us32/_0015_ ;
wire \us32/_0016_ ;
wire \us32/_0017_ ;
wire \us32/_0019_ ;
wire \us32/_0020_ ;
wire \us32/_0022_ ;
wire \us32/_0024_ ;
wire \us32/_0025_ ;
wire \us32/_0026_ ;
wire \us32/_0027_ ;
wire \us32/_0030_ ;
wire \us32/_0032_ ;
wire \us32/_0033_ ;
wire \us32/_0034_ ;
wire \us32/_0035_ ;
wire \us32/_0037_ ;
wire \us32/_0038_ ;
wire \us32/_0039_ ;
wire \us32/_0040_ ;
wire \us32/_0041_ ;
wire \us32/_0042_ ;
wire \us32/_0043_ ;
wire \us32/_0045_ ;
wire \us32/_0046_ ;
wire \us32/_0047_ ;
wire \us32/_0049_ ;
wire \us32/_0050_ ;
wire \us32/_0051_ ;
wire \us32/_0052_ ;
wire \us32/_0053_ ;
wire \us32/_0054_ ;
wire \us32/_0056_ ;
wire \us32/_0057_ ;
wire \us32/_0058_ ;
wire \us32/_0060_ ;
wire \us32/_0061_ ;
wire \us32/_0062_ ;
wire \us32/_0064_ ;
wire \us32/_0065_ ;
wire \us32/_0066_ ;
wire \us32/_0067_ ;
wire \us32/_0069_ ;
wire \us32/_0070_ ;
wire \us32/_0072_ ;
wire \us32/_0073_ ;
wire \us32/_0074_ ;
wire \us32/_0075_ ;
wire \us32/_0076_ ;
wire \us32/_0077_ ;
wire \us32/_0078_ ;
wire \us32/_0079_ ;
wire \us32/_0081_ ;
wire \us32/_0082_ ;
wire \us32/_0085_ ;
wire \us32/_0086_ ;
wire \us32/_0087_ ;
wire \us32/_0088_ ;
wire \us32/_0089_ ;
wire \us32/_0090_ ;
wire \us32/_0091_ ;
wire \us32/_0092_ ;
wire \us32/_0093_ ;
wire \us32/_0094_ ;
wire \us32/_0095_ ;
wire \us32/_0096_ ;
wire \us32/_0097_ ;
wire \us32/_0098_ ;
wire \us32/_0099_ ;
wire \us32/_0100_ ;
wire \us32/_0101_ ;
wire \us32/_0102_ ;
wire \us32/_0103_ ;
wire \us32/_0104_ ;
wire \us32/_0105_ ;
wire \us32/_0106_ ;
wire \us32/_0108_ ;
wire \us32/_0109_ ;
wire \us32/_0110_ ;
wire \us32/_0111_ ;
wire \us32/_0113_ ;
wire \us32/_0114_ ;
wire \us32/_0115_ ;
wire \us32/_0116_ ;
wire \us32/_0117_ ;
wire \us32/_0118_ ;
wire \us32/_0119_ ;
wire \us32/_0120_ ;
wire \us32/_0121_ ;
wire \us32/_0122_ ;
wire \us32/_0123_ ;
wire \us32/_0124_ ;
wire \us32/_0126_ ;
wire \us32/_0127_ ;
wire \us32/_0128_ ;
wire \us32/_0129_ ;
wire \us32/_0130_ ;
wire \us32/_0132_ ;
wire \us32/_0133_ ;
wire \us32/_0134_ ;
wire \us32/_0135_ ;
wire \us32/_0136_ ;
wire \us32/_0137_ ;
wire \us32/_0139_ ;
wire \us32/_0140_ ;
wire \us32/_0141_ ;
wire \us32/_0142_ ;
wire \us32/_0144_ ;
wire \us32/_0145_ ;
wire \us32/_0146_ ;
wire \us32/_0147_ ;
wire \us32/_0148_ ;
wire \us32/_0149_ ;
wire \us32/_0150_ ;
wire \us32/_0151_ ;
wire \us32/_0153_ ;
wire \us32/_0154_ ;
wire \us32/_0155_ ;
wire \us32/_0156_ ;
wire \us32/_0157_ ;
wire \us32/_0158_ ;
wire \us32/_0159_ ;
wire \us32/_0161_ ;
wire \us32/_0162_ ;
wire \us32/_0163_ ;
wire \us32/_0164_ ;
wire \us32/_0165_ ;
wire \us32/_0166_ ;
wire \us32/_0167_ ;
wire \us32/_0168_ ;
wire \us32/_0169_ ;
wire \us32/_0170_ ;
wire \us32/_0171_ ;
wire \us32/_0172_ ;
wire \us32/_0174_ ;
wire \us32/_0175_ ;
wire \us32/_0176_ ;
wire \us32/_0177_ ;
wire \us32/_0178_ ;
wire \us32/_0179_ ;
wire \us32/_0180_ ;
wire \us32/_0181_ ;
wire \us32/_0182_ ;
wire \us32/_0183_ ;
wire \us32/_0184_ ;
wire \us32/_0185_ ;
wire \us32/_0186_ ;
wire \us32/_0187_ ;
wire \us32/_0188_ ;
wire \us32/_0189_ ;
wire \us32/_0190_ ;
wire \us32/_0191_ ;
wire \us32/_0192_ ;
wire \us32/_0193_ ;
wire \us32/_0194_ ;
wire \us32/_0195_ ;
wire \us32/_0196_ ;
wire \us32/_0197_ ;
wire \us32/_0198_ ;
wire \us32/_0199_ ;
wire \us32/_0200_ ;
wire \us32/_0201_ ;
wire \us32/_0202_ ;
wire \us32/_0203_ ;
wire \us32/_0204_ ;
wire \us32/_0205_ ;
wire \us32/_0206_ ;
wire \us32/_0207_ ;
wire \us32/_0208_ ;
wire \us32/_0209_ ;
wire \us32/_0210_ ;
wire \us32/_0211_ ;
wire \us32/_0212_ ;
wire \us32/_0213_ ;
wire \us32/_0214_ ;
wire \us32/_0215_ ;
wire \us32/_0217_ ;
wire \us32/_0219_ ;
wire \us32/_0220_ ;
wire \us32/_0221_ ;
wire \us32/_0222_ ;
wire \us32/_0223_ ;
wire \us32/_0224_ ;
wire \us32/_0225_ ;
wire \us32/_0226_ ;
wire \us32/_0227_ ;
wire \us32/_0228_ ;
wire \us32/_0229_ ;
wire \us32/_0230_ ;
wire \us32/_0231_ ;
wire \us32/_0232_ ;
wire \us32/_0233_ ;
wire \us32/_0234_ ;
wire \us32/_0235_ ;
wire \us32/_0236_ ;
wire \us32/_0237_ ;
wire \us32/_0238_ ;
wire \us32/_0239_ ;
wire \us32/_0240_ ;
wire \us32/_0241_ ;
wire \us32/_0242_ ;
wire \us32/_0243_ ;
wire \us32/_0244_ ;
wire \us32/_0245_ ;
wire \us32/_0246_ ;
wire \us32/_0247_ ;
wire \us32/_0248_ ;
wire \us32/_0249_ ;
wire \us32/_0250_ ;
wire \us32/_0251_ ;
wire \us32/_0252_ ;
wire \us32/_0253_ ;
wire \us32/_0254_ ;
wire \us32/_0255_ ;
wire \us32/_0256_ ;
wire \us32/_0257_ ;
wire \us32/_0258_ ;
wire \us32/_0259_ ;
wire \us32/_0260_ ;
wire \us32/_0261_ ;
wire \us32/_0263_ ;
wire \us32/_0264_ ;
wire \us32/_0265_ ;
wire \us32/_0266_ ;
wire \us32/_0267_ ;
wire \us32/_0268_ ;
wire \us32/_0269_ ;
wire \us32/_0270_ ;
wire \us32/_0271_ ;
wire \us32/_0272_ ;
wire \us32/_0273_ ;
wire \us32/_0274_ ;
wire \us32/_0275_ ;
wire \us32/_0276_ ;
wire \us32/_0277_ ;
wire \us32/_0278_ ;
wire \us32/_0279_ ;
wire \us32/_0280_ ;
wire \us32/_0281_ ;
wire \us32/_0283_ ;
wire \us32/_0284_ ;
wire \us32/_0285_ ;
wire \us32/_0286_ ;
wire \us32/_0287_ ;
wire \us32/_0288_ ;
wire \us32/_0289_ ;
wire \us32/_0290_ ;
wire \us32/_0291_ ;
wire \us32/_0293_ ;
wire \us32/_0294_ ;
wire \us32/_0295_ ;
wire \us32/_0296_ ;
wire \us32/_0297_ ;
wire \us32/_0298_ ;
wire \us32/_0299_ ;
wire \us32/_0300_ ;
wire \us32/_0301_ ;
wire \us32/_0302_ ;
wire \us32/_0303_ ;
wire \us32/_0304_ ;
wire \us32/_0305_ ;
wire \us32/_0306_ ;
wire \us32/_0307_ ;
wire \us32/_0308_ ;
wire \us32/_0309_ ;
wire \us32/_0310_ ;
wire \us32/_0311_ ;
wire \us32/_0312_ ;
wire \us32/_0313_ ;
wire \us32/_0314_ ;
wire \us32/_0315_ ;
wire \us32/_0316_ ;
wire \us32/_0317_ ;
wire \us32/_0318_ ;
wire \us32/_0319_ ;
wire \us32/_0320_ ;
wire \us32/_0321_ ;
wire \us32/_0322_ ;
wire \us32/_0323_ ;
wire \us32/_0324_ ;
wire \us32/_0325_ ;
wire \us32/_0326_ ;
wire \us32/_0327_ ;
wire \us32/_0328_ ;
wire \us32/_0329_ ;
wire \us32/_0330_ ;
wire \us32/_0331_ ;
wire \us32/_0332_ ;
wire \us32/_0333_ ;
wire \us32/_0334_ ;
wire \us32/_0335_ ;
wire \us32/_0337_ ;
wire \us32/_0338_ ;
wire \us32/_0339_ ;
wire \us32/_0340_ ;
wire \us32/_0341_ ;
wire \us32/_0342_ ;
wire \us32/_0343_ ;
wire \us32/_0344_ ;
wire \us32/_0345_ ;
wire \us32/_0347_ ;
wire \us32/_0348_ ;
wire \us32/_0349_ ;
wire \us32/_0350_ ;
wire \us32/_0351_ ;
wire \us32/_0352_ ;
wire \us32/_0353_ ;
wire \us32/_0354_ ;
wire \us32/_0355_ ;
wire \us32/_0356_ ;
wire \us32/_0357_ ;
wire \us32/_0358_ ;
wire \us32/_0359_ ;
wire \us32/_0360_ ;
wire \us32/_0361_ ;
wire \us32/_0362_ ;
wire \us32/_0363_ ;
wire \us32/_0365_ ;
wire \us32/_0366_ ;
wire \us32/_0367_ ;
wire \us32/_0368_ ;
wire \us32/_0370_ ;
wire \us32/_0371_ ;
wire \us32/_0372_ ;
wire \us32/_0373_ ;
wire \us32/_0374_ ;
wire \us32/_0375_ ;
wire \us32/_0376_ ;
wire \us32/_0377_ ;
wire \us32/_0378_ ;
wire \us32/_0379_ ;
wire \us32/_0380_ ;
wire \us32/_0381_ ;
wire \us32/_0382_ ;
wire \us32/_0383_ ;
wire \us32/_0384_ ;
wire \us32/_0385_ ;
wire \us32/_0386_ ;
wire \us32/_0387_ ;
wire \us32/_0388_ ;
wire \us32/_0389_ ;
wire \us32/_0390_ ;
wire \us32/_0391_ ;
wire \us32/_0392_ ;
wire \us32/_0393_ ;
wire \us32/_0394_ ;
wire \us32/_0395_ ;
wire \us32/_0396_ ;
wire \us32/_0397_ ;
wire \us32/_0398_ ;
wire \us32/_0399_ ;
wire \us32/_0400_ ;
wire \us32/_0401_ ;
wire \us32/_0402_ ;
wire \us32/_0403_ ;
wire \us32/_0404_ ;
wire \us32/_0405_ ;
wire \us32/_0406_ ;
wire \us32/_0407_ ;
wire \us32/_0408_ ;
wire \us32/_0409_ ;
wire \us32/_0410_ ;
wire \us32/_0411_ ;
wire \us32/_0412_ ;
wire \us32/_0413_ ;
wire \us32/_0414_ ;
wire \us32/_0415_ ;
wire \us32/_0416_ ;
wire \us32/_0417_ ;
wire \us32/_0418_ ;
wire \us32/_0419_ ;
wire \us32/_0420_ ;
wire \us32/_0421_ ;
wire \us32/_0422_ ;
wire \us32/_0424_ ;
wire \us32/_0425_ ;
wire \us32/_0426_ ;
wire \us32/_0427_ ;
wire \us32/_0428_ ;
wire \us32/_0429_ ;
wire \us32/_0430_ ;
wire \us32/_0431_ ;
wire \us32/_0432_ ;
wire \us32/_0433_ ;
wire \us32/_0434_ ;
wire \us32/_0435_ ;
wire \us32/_0436_ ;
wire \us32/_0437_ ;
wire \us32/_0438_ ;
wire \us32/_0439_ ;
wire \us32/_0440_ ;
wire \us32/_0441_ ;
wire \us32/_0442_ ;
wire \us32/_0443_ ;
wire \us32/_0444_ ;
wire \us32/_0446_ ;
wire \us32/_0447_ ;
wire \us32/_0448_ ;
wire \us32/_0449_ ;
wire \us32/_0450_ ;
wire \us32/_0451_ ;
wire \us32/_0452_ ;
wire \us32/_0453_ ;
wire \us32/_0454_ ;
wire \us32/_0455_ ;
wire \us32/_0457_ ;
wire \us32/_0458_ ;
wire \us32/_0459_ ;
wire \us32/_0460_ ;
wire \us32/_0461_ ;
wire \us32/_0462_ ;
wire \us32/_0463_ ;
wire \us32/_0464_ ;
wire \us32/_0465_ ;
wire \us32/_0466_ ;
wire \us32/_0467_ ;
wire \us32/_0468_ ;
wire \us32/_0469_ ;
wire \us32/_0470_ ;
wire \us32/_0471_ ;
wire \us32/_0472_ ;
wire \us32/_0473_ ;
wire \us32/_0474_ ;
wire \us32/_0475_ ;
wire \us32/_0476_ ;
wire \us32/_0477_ ;
wire \us32/_0478_ ;
wire \us32/_0479_ ;
wire \us32/_0480_ ;
wire \us32/_0481_ ;
wire \us32/_0482_ ;
wire \us32/_0483_ ;
wire \us32/_0484_ ;
wire \us32/_0485_ ;
wire \us32/_0486_ ;
wire \us32/_0487_ ;
wire \us32/_0488_ ;
wire \us32/_0490_ ;
wire \us32/_0491_ ;
wire \us32/_0492_ ;
wire \us32/_0493_ ;
wire \us32/_0494_ ;
wire \us32/_0495_ ;
wire \us32/_0496_ ;
wire \us32/_0497_ ;
wire \us32/_0498_ ;
wire \us32/_0499_ ;
wire \us32/_0500_ ;
wire \us32/_0501_ ;
wire \us32/_0502_ ;
wire \us32/_0503_ ;
wire \us32/_0504_ ;
wire \us32/_0505_ ;
wire \us32/_0506_ ;
wire \us32/_0507_ ;
wire \us32/_0508_ ;
wire \us32/_0509_ ;
wire \us32/_0510_ ;
wire \us32/_0511_ ;
wire \us32/_0512_ ;
wire \us32/_0513_ ;
wire \us32/_0514_ ;
wire \us32/_0515_ ;
wire \us32/_0516_ ;
wire \us32/_0517_ ;
wire \us32/_0518_ ;
wire \us32/_0519_ ;
wire \us32/_0520_ ;
wire \us32/_0521_ ;
wire \us32/_0522_ ;
wire \us32/_0523_ ;
wire \us32/_0524_ ;
wire \us32/_0525_ ;
wire \us32/_0526_ ;
wire \us32/_0527_ ;
wire \us32/_0528_ ;
wire \us32/_0529_ ;
wire \us32/_0530_ ;
wire \us32/_0531_ ;
wire \us32/_0532_ ;
wire \us32/_0533_ ;
wire \us32/_0534_ ;
wire \us32/_0535_ ;
wire \us32/_0536_ ;
wire \us32/_0537_ ;
wire \us32/_0538_ ;
wire \us32/_0539_ ;
wire \us32/_0540_ ;
wire \us32/_0541_ ;
wire \us32/_0542_ ;
wire \us32/_0544_ ;
wire \us32/_0545_ ;
wire \us32/_0546_ ;
wire \us32/_0547_ ;
wire \us32/_0548_ ;
wire \us32/_0549_ ;
wire \us32/_0550_ ;
wire \us32/_0551_ ;
wire \us32/_0552_ ;
wire \us32/_0553_ ;
wire \us32/_0554_ ;
wire \us32/_0555_ ;
wire \us32/_0556_ ;
wire \us32/_0557_ ;
wire \us32/_0558_ ;
wire \us32/_0559_ ;
wire \us32/_0560_ ;
wire \us32/_0561_ ;
wire \us32/_0562_ ;
wire \us32/_0563_ ;
wire \us32/_0565_ ;
wire \us32/_0566_ ;
wire \us32/_0567_ ;
wire \us32/_0568_ ;
wire \us32/_0569_ ;
wire \us32/_0570_ ;
wire \us32/_0571_ ;
wire \us32/_0572_ ;
wire \us32/_0573_ ;
wire \us32/_0574_ ;
wire \us32/_0575_ ;
wire \us32/_0576_ ;
wire \us32/_0577_ ;
wire \us32/_0578_ ;
wire \us32/_0579_ ;
wire \us32/_0580_ ;
wire \us32/_0581_ ;
wire \us32/_0582_ ;
wire \us32/_0583_ ;
wire \us32/_0584_ ;
wire \us32/_0585_ ;
wire \us32/_0586_ ;
wire \us32/_0587_ ;
wire \us32/_0588_ ;
wire \us32/_0589_ ;
wire \us32/_0590_ ;
wire \us32/_0591_ ;
wire \us32/_0592_ ;
wire \us32/_0593_ ;
wire \us32/_0594_ ;
wire \us32/_0595_ ;
wire \us32/_0596_ ;
wire \us32/_0598_ ;
wire \us32/_0599_ ;
wire \us32/_0600_ ;
wire \us32/_0601_ ;
wire \us32/_0602_ ;
wire \us32/_0603_ ;
wire \us32/_0604_ ;
wire \us32/_0605_ ;
wire \us32/_0606_ ;
wire \us32/_0607_ ;
wire \us32/_0608_ ;
wire \us32/_0609_ ;
wire \us32/_0610_ ;
wire \us32/_0611_ ;
wire \us32/_0612_ ;
wire \us32/_0613_ ;
wire \us32/_0614_ ;
wire \us32/_0615_ ;
wire \us32/_0616_ ;
wire \us32/_0617_ ;
wire \us32/_0618_ ;
wire \us32/_0619_ ;
wire \us32/_0620_ ;
wire \us32/_0621_ ;
wire \us32/_0622_ ;
wire \us32/_0623_ ;
wire \us32/_0624_ ;
wire \us32/_0625_ ;
wire \us32/_0626_ ;
wire \us32/_0627_ ;
wire \us32/_0628_ ;
wire \us32/_0629_ ;
wire \us32/_0630_ ;
wire \us32/_0631_ ;
wire \us32/_0632_ ;
wire \us32/_0633_ ;
wire \us32/_0634_ ;
wire \us32/_0635_ ;
wire \us32/_0636_ ;
wire \us32/_0637_ ;
wire \us32/_0638_ ;
wire \us32/_0639_ ;
wire \us32/_0640_ ;
wire \us32/_0641_ ;
wire \us32/_0642_ ;
wire \us32/_0643_ ;
wire \us32/_0644_ ;
wire \us32/_0645_ ;
wire \us32/_0646_ ;
wire \us32/_0647_ ;
wire \us32/_0648_ ;
wire \us32/_0649_ ;
wire \us32/_0650_ ;
wire \us32/_0652_ ;
wire \us32/_0653_ ;
wire \us32/_0654_ ;
wire \us32/_0655_ ;
wire \us32/_0656_ ;
wire \us32/_0657_ ;
wire \us32/_0658_ ;
wire \us32/_0659_ ;
wire \us32/_0660_ ;
wire \us32/_0661_ ;
wire \us32/_0662_ ;
wire \us32/_0663_ ;
wire \us32/_0664_ ;
wire \us32/_0665_ ;
wire \us32/_0666_ ;
wire \us32/_0667_ ;
wire \us32/_0668_ ;
wire \us32/_0669_ ;
wire \us32/_0670_ ;
wire \us32/_0671_ ;
wire \us32/_0673_ ;
wire \us32/_0674_ ;
wire \us32/_0675_ ;
wire \us32/_0676_ ;
wire \us32/_0677_ ;
wire \us32/_0678_ ;
wire \us32/_0679_ ;
wire \us32/_0680_ ;
wire \us32/_0681_ ;
wire \us32/_0682_ ;
wire \us32/_0683_ ;
wire \us32/_0684_ ;
wire \us32/_0685_ ;
wire \us32/_0686_ ;
wire \us32/_0687_ ;
wire \us32/_0688_ ;
wire \us32/_0689_ ;
wire \us32/_0690_ ;
wire \us32/_0691_ ;
wire \us32/_0692_ ;
wire \us32/_0693_ ;
wire \us32/_0694_ ;
wire \us32/_0695_ ;
wire \us32/_0696_ ;
wire \us32/_0697_ ;
wire \us32/_0698_ ;
wire \us32/_0699_ ;
wire \us32/_0700_ ;
wire \us32/_0701_ ;
wire \us32/_0702_ ;
wire \us32/_0703_ ;
wire \us32/_0704_ ;
wire \us32/_0705_ ;
wire \us32/_0706_ ;
wire \us32/_0707_ ;
wire \us32/_0708_ ;
wire \us32/_0709_ ;
wire \us32/_0710_ ;
wire \us32/_0711_ ;
wire \us32/_0712_ ;
wire \us32/_0713_ ;
wire \us32/_0714_ ;
wire \us32/_0715_ ;
wire \us32/_0717_ ;
wire \us32/_0718_ ;
wire \us32/_0719_ ;
wire \us32/_0720_ ;
wire \us32/_0721_ ;
wire \us32/_0722_ ;
wire \us32/_0723_ ;
wire \us32/_0724_ ;
wire \us32/_0725_ ;
wire \us32/_0726_ ;
wire \us32/_0727_ ;
wire \us32/_0728_ ;
wire \us32/_0729_ ;
wire \us32/_0730_ ;
wire \us32/_0731_ ;
wire \us32/_0733_ ;
wire \us32/_0734_ ;
wire \us32/_0735_ ;
wire \us32/_0736_ ;
wire \us32/_0738_ ;
wire \us32/_0739_ ;
wire \us32/_0740_ ;
wire \us32/_0741_ ;
wire \us32/_0742_ ;
wire \us32/_0744_ ;
wire \us32/_0745_ ;
wire \us32/_0746_ ;
wire \us32/_0748_ ;
wire \us32/_0749_ ;
wire \us32/_0750_ ;
wire \us32/_0752_ ;
wire \us33/_0008_ ;
wire \us33/_0009_ ;
wire \us33/_0010_ ;
wire \us33/_0011_ ;
wire \us33/_0012_ ;
wire \us33/_0013_ ;
wire \us33/_0014_ ;
wire \us33/_0015_ ;
wire \us33/_0016_ ;
wire \us33/_0017_ ;
wire \us33/_0019_ ;
wire \us33/_0020_ ;
wire \us33/_0022_ ;
wire \us33/_0024_ ;
wire \us33/_0025_ ;
wire \us33/_0026_ ;
wire \us33/_0027_ ;
wire \us33/_0030_ ;
wire \us33/_0032_ ;
wire \us33/_0033_ ;
wire \us33/_0034_ ;
wire \us33/_0035_ ;
wire \us33/_0037_ ;
wire \us33/_0038_ ;
wire \us33/_0039_ ;
wire \us33/_0040_ ;
wire \us33/_0041_ ;
wire \us33/_0042_ ;
wire \us33/_0043_ ;
wire \us33/_0045_ ;
wire \us33/_0046_ ;
wire \us33/_0047_ ;
wire \us33/_0049_ ;
wire \us33/_0050_ ;
wire \us33/_0051_ ;
wire \us33/_0052_ ;
wire \us33/_0053_ ;
wire \us33/_0054_ ;
wire \us33/_0057_ ;
wire \us33/_0058_ ;
wire \us33/_0060_ ;
wire \us33/_0061_ ;
wire \us33/_0062_ ;
wire \us33/_0064_ ;
wire \us33/_0065_ ;
wire \us33/_0066_ ;
wire \us33/_0067_ ;
wire \us33/_0069_ ;
wire \us33/_0070_ ;
wire \us33/_0072_ ;
wire \us33/_0073_ ;
wire \us33/_0074_ ;
wire \us33/_0075_ ;
wire \us33/_0076_ ;
wire \us33/_0077_ ;
wire \us33/_0078_ ;
wire \us33/_0079_ ;
wire \us33/_0081_ ;
wire \us33/_0082_ ;
wire \us33/_0085_ ;
wire \us33/_0086_ ;
wire \us33/_0087_ ;
wire \us33/_0088_ ;
wire \us33/_0089_ ;
wire \us33/_0090_ ;
wire \us33/_0091_ ;
wire \us33/_0092_ ;
wire \us33/_0093_ ;
wire \us33/_0094_ ;
wire \us33/_0095_ ;
wire \us33/_0096_ ;
wire \us33/_0097_ ;
wire \us33/_0098_ ;
wire \us33/_0099_ ;
wire \us33/_0100_ ;
wire \us33/_0101_ ;
wire \us33/_0102_ ;
wire \us33/_0103_ ;
wire \us33/_0104_ ;
wire \us33/_0105_ ;
wire \us33/_0106_ ;
wire \us33/_0108_ ;
wire \us33/_0109_ ;
wire \us33/_0110_ ;
wire \us33/_0111_ ;
wire \us33/_0113_ ;
wire \us33/_0114_ ;
wire \us33/_0115_ ;
wire \us33/_0116_ ;
wire \us33/_0117_ ;
wire \us33/_0118_ ;
wire \us33/_0119_ ;
wire \us33/_0120_ ;
wire \us33/_0121_ ;
wire \us33/_0122_ ;
wire \us33/_0123_ ;
wire \us33/_0124_ ;
wire \us33/_0126_ ;
wire \us33/_0127_ ;
wire \us33/_0128_ ;
wire \us33/_0129_ ;
wire \us33/_0130_ ;
wire \us33/_0132_ ;
wire \us33/_0133_ ;
wire \us33/_0134_ ;
wire \us33/_0135_ ;
wire \us33/_0136_ ;
wire \us33/_0137_ ;
wire \us33/_0139_ ;
wire \us33/_0140_ ;
wire \us33/_0141_ ;
wire \us33/_0142_ ;
wire \us33/_0144_ ;
wire \us33/_0145_ ;
wire \us33/_0146_ ;
wire \us33/_0147_ ;
wire \us33/_0148_ ;
wire \us33/_0149_ ;
wire \us33/_0150_ ;
wire \us33/_0151_ ;
wire \us33/_0153_ ;
wire \us33/_0154_ ;
wire \us33/_0155_ ;
wire \us33/_0156_ ;
wire \us33/_0157_ ;
wire \us33/_0158_ ;
wire \us33/_0159_ ;
wire \us33/_0161_ ;
wire \us33/_0162_ ;
wire \us33/_0163_ ;
wire \us33/_0164_ ;
wire \us33/_0165_ ;
wire \us33/_0166_ ;
wire \us33/_0167_ ;
wire \us33/_0168_ ;
wire \us33/_0169_ ;
wire \us33/_0170_ ;
wire \us33/_0171_ ;
wire \us33/_0172_ ;
wire \us33/_0174_ ;
wire \us33/_0175_ ;
wire \us33/_0176_ ;
wire \us33/_0177_ ;
wire \us33/_0178_ ;
wire \us33/_0179_ ;
wire \us33/_0180_ ;
wire \us33/_0181_ ;
wire \us33/_0182_ ;
wire \us33/_0183_ ;
wire \us33/_0184_ ;
wire \us33/_0185_ ;
wire \us33/_0186_ ;
wire \us33/_0187_ ;
wire \us33/_0188_ ;
wire \us33/_0189_ ;
wire \us33/_0190_ ;
wire \us33/_0191_ ;
wire \us33/_0192_ ;
wire \us33/_0193_ ;
wire \us33/_0194_ ;
wire \us33/_0195_ ;
wire \us33/_0196_ ;
wire \us33/_0197_ ;
wire \us33/_0198_ ;
wire \us33/_0199_ ;
wire \us33/_0200_ ;
wire \us33/_0201_ ;
wire \us33/_0202_ ;
wire \us33/_0203_ ;
wire \us33/_0204_ ;
wire \us33/_0205_ ;
wire \us33/_0206_ ;
wire \us33/_0207_ ;
wire \us33/_0208_ ;
wire \us33/_0209_ ;
wire \us33/_0210_ ;
wire \us33/_0211_ ;
wire \us33/_0212_ ;
wire \us33/_0213_ ;
wire \us33/_0214_ ;
wire \us33/_0215_ ;
wire \us33/_0217_ ;
wire \us33/_0219_ ;
wire \us33/_0220_ ;
wire \us33/_0221_ ;
wire \us33/_0222_ ;
wire \us33/_0223_ ;
wire \us33/_0224_ ;
wire \us33/_0225_ ;
wire \us33/_0226_ ;
wire \us33/_0227_ ;
wire \us33/_0228_ ;
wire \us33/_0229_ ;
wire \us33/_0230_ ;
wire \us33/_0231_ ;
wire \us33/_0232_ ;
wire \us33/_0233_ ;
wire \us33/_0234_ ;
wire \us33/_0235_ ;
wire \us33/_0236_ ;
wire \us33/_0237_ ;
wire \us33/_0238_ ;
wire \us33/_0239_ ;
wire \us33/_0240_ ;
wire \us33/_0241_ ;
wire \us33/_0242_ ;
wire \us33/_0243_ ;
wire \us33/_0244_ ;
wire \us33/_0245_ ;
wire \us33/_0246_ ;
wire \us33/_0247_ ;
wire \us33/_0248_ ;
wire \us33/_0249_ ;
wire \us33/_0250_ ;
wire \us33/_0251_ ;
wire \us33/_0252_ ;
wire \us33/_0253_ ;
wire \us33/_0254_ ;
wire \us33/_0255_ ;
wire \us33/_0256_ ;
wire \us33/_0257_ ;
wire \us33/_0258_ ;
wire \us33/_0259_ ;
wire \us33/_0260_ ;
wire \us33/_0261_ ;
wire \us33/_0263_ ;
wire \us33/_0264_ ;
wire \us33/_0265_ ;
wire \us33/_0266_ ;
wire \us33/_0267_ ;
wire \us33/_0268_ ;
wire \us33/_0269_ ;
wire \us33/_0270_ ;
wire \us33/_0271_ ;
wire \us33/_0272_ ;
wire \us33/_0273_ ;
wire \us33/_0274_ ;
wire \us33/_0275_ ;
wire \us33/_0276_ ;
wire \us33/_0277_ ;
wire \us33/_0278_ ;
wire \us33/_0279_ ;
wire \us33/_0280_ ;
wire \us33/_0281_ ;
wire \us33/_0283_ ;
wire \us33/_0284_ ;
wire \us33/_0285_ ;
wire \us33/_0286_ ;
wire \us33/_0287_ ;
wire \us33/_0288_ ;
wire \us33/_0289_ ;
wire \us33/_0290_ ;
wire \us33/_0291_ ;
wire \us33/_0292_ ;
wire \us33/_0293_ ;
wire \us33/_0294_ ;
wire \us33/_0295_ ;
wire \us33/_0296_ ;
wire \us33/_0297_ ;
wire \us33/_0298_ ;
wire \us33/_0299_ ;
wire \us33/_0300_ ;
wire \us33/_0301_ ;
wire \us33/_0302_ ;
wire \us33/_0303_ ;
wire \us33/_0304_ ;
wire \us33/_0305_ ;
wire \us33/_0306_ ;
wire \us33/_0307_ ;
wire \us33/_0308_ ;
wire \us33/_0309_ ;
wire \us33/_0310_ ;
wire \us33/_0311_ ;
wire \us33/_0312_ ;
wire \us33/_0313_ ;
wire \us33/_0314_ ;
wire \us33/_0315_ ;
wire \us33/_0316_ ;
wire \us33/_0317_ ;
wire \us33/_0318_ ;
wire \us33/_0319_ ;
wire \us33/_0320_ ;
wire \us33/_0321_ ;
wire \us33/_0322_ ;
wire \us33/_0323_ ;
wire \us33/_0324_ ;
wire \us33/_0325_ ;
wire \us33/_0326_ ;
wire \us33/_0327_ ;
wire \us33/_0328_ ;
wire \us33/_0329_ ;
wire \us33/_0330_ ;
wire \us33/_0331_ ;
wire \us33/_0332_ ;
wire \us33/_0333_ ;
wire \us33/_0334_ ;
wire \us33/_0335_ ;
wire \us33/_0337_ ;
wire \us33/_0338_ ;
wire \us33/_0339_ ;
wire \us33/_0340_ ;
wire \us33/_0341_ ;
wire \us33/_0342_ ;
wire \us33/_0343_ ;
wire \us33/_0344_ ;
wire \us33/_0345_ ;
wire \us33/_0347_ ;
wire \us33/_0348_ ;
wire \us33/_0349_ ;
wire \us33/_0350_ ;
wire \us33/_0351_ ;
wire \us33/_0352_ ;
wire \us33/_0353_ ;
wire \us33/_0354_ ;
wire \us33/_0355_ ;
wire \us33/_0356_ ;
wire \us33/_0357_ ;
wire \us33/_0358_ ;
wire \us33/_0359_ ;
wire \us33/_0360_ ;
wire \us33/_0361_ ;
wire \us33/_0362_ ;
wire \us33/_0363_ ;
wire \us33/_0365_ ;
wire \us33/_0366_ ;
wire \us33/_0367_ ;
wire \us33/_0368_ ;
wire \us33/_0370_ ;
wire \us33/_0371_ ;
wire \us33/_0372_ ;
wire \us33/_0373_ ;
wire \us33/_0374_ ;
wire \us33/_0375_ ;
wire \us33/_0376_ ;
wire \us33/_0377_ ;
wire \us33/_0378_ ;
wire \us33/_0379_ ;
wire \us33/_0380_ ;
wire \us33/_0381_ ;
wire \us33/_0382_ ;
wire \us33/_0383_ ;
wire \us33/_0384_ ;
wire \us33/_0385_ ;
wire \us33/_0386_ ;
wire \us33/_0387_ ;
wire \us33/_0388_ ;
wire \us33/_0389_ ;
wire \us33/_0390_ ;
wire \us33/_0391_ ;
wire \us33/_0392_ ;
wire \us33/_0393_ ;
wire \us33/_0394_ ;
wire \us33/_0395_ ;
wire \us33/_0396_ ;
wire \us33/_0397_ ;
wire \us33/_0398_ ;
wire \us33/_0399_ ;
wire \us33/_0400_ ;
wire \us33/_0401_ ;
wire \us33/_0402_ ;
wire \us33/_0403_ ;
wire \us33/_0404_ ;
wire \us33/_0405_ ;
wire \us33/_0406_ ;
wire \us33/_0407_ ;
wire \us33/_0408_ ;
wire \us33/_0409_ ;
wire \us33/_0410_ ;
wire \us33/_0411_ ;
wire \us33/_0412_ ;
wire \us33/_0413_ ;
wire \us33/_0414_ ;
wire \us33/_0415_ ;
wire \us33/_0416_ ;
wire \us33/_0417_ ;
wire \us33/_0418_ ;
wire \us33/_0419_ ;
wire \us33/_0420_ ;
wire \us33/_0421_ ;
wire \us33/_0422_ ;
wire \us33/_0424_ ;
wire \us33/_0425_ ;
wire \us33/_0426_ ;
wire \us33/_0427_ ;
wire \us33/_0428_ ;
wire \us33/_0429_ ;
wire \us33/_0430_ ;
wire \us33/_0431_ ;
wire \us33/_0432_ ;
wire \us33/_0433_ ;
wire \us33/_0434_ ;
wire \us33/_0435_ ;
wire \us33/_0436_ ;
wire \us33/_0437_ ;
wire \us33/_0438_ ;
wire \us33/_0439_ ;
wire \us33/_0440_ ;
wire \us33/_0441_ ;
wire \us33/_0442_ ;
wire \us33/_0443_ ;
wire \us33/_0444_ ;
wire \us33/_0446_ ;
wire \us33/_0447_ ;
wire \us33/_0448_ ;
wire \us33/_0449_ ;
wire \us33/_0450_ ;
wire \us33/_0451_ ;
wire \us33/_0452_ ;
wire \us33/_0453_ ;
wire \us33/_0454_ ;
wire \us33/_0455_ ;
wire \us33/_0457_ ;
wire \us33/_0458_ ;
wire \us33/_0459_ ;
wire \us33/_0460_ ;
wire \us33/_0461_ ;
wire \us33/_0462_ ;
wire \us33/_0463_ ;
wire \us33/_0464_ ;
wire \us33/_0465_ ;
wire \us33/_0466_ ;
wire \us33/_0467_ ;
wire \us33/_0468_ ;
wire \us33/_0469_ ;
wire \us33/_0470_ ;
wire \us33/_0471_ ;
wire \us33/_0472_ ;
wire \us33/_0473_ ;
wire \us33/_0474_ ;
wire \us33/_0475_ ;
wire \us33/_0476_ ;
wire \us33/_0477_ ;
wire \us33/_0478_ ;
wire \us33/_0479_ ;
wire \us33/_0480_ ;
wire \us33/_0481_ ;
wire \us33/_0482_ ;
wire \us33/_0483_ ;
wire \us33/_0484_ ;
wire \us33/_0485_ ;
wire \us33/_0486_ ;
wire \us33/_0487_ ;
wire \us33/_0488_ ;
wire \us33/_0490_ ;
wire \us33/_0491_ ;
wire \us33/_0492_ ;
wire \us33/_0493_ ;
wire \us33/_0494_ ;
wire \us33/_0495_ ;
wire \us33/_0496_ ;
wire \us33/_0497_ ;
wire \us33/_0498_ ;
wire \us33/_0499_ ;
wire \us33/_0500_ ;
wire \us33/_0501_ ;
wire \us33/_0502_ ;
wire \us33/_0503_ ;
wire \us33/_0504_ ;
wire \us33/_0505_ ;
wire \us33/_0506_ ;
wire \us33/_0507_ ;
wire \us33/_0508_ ;
wire \us33/_0509_ ;
wire \us33/_0510_ ;
wire \us33/_0511_ ;
wire \us33/_0512_ ;
wire \us33/_0513_ ;
wire \us33/_0514_ ;
wire \us33/_0515_ ;
wire \us33/_0516_ ;
wire \us33/_0517_ ;
wire \us33/_0518_ ;
wire \us33/_0519_ ;
wire \us33/_0520_ ;
wire \us33/_0521_ ;
wire \us33/_0522_ ;
wire \us33/_0523_ ;
wire \us33/_0524_ ;
wire \us33/_0525_ ;
wire \us33/_0526_ ;
wire \us33/_0527_ ;
wire \us33/_0528_ ;
wire \us33/_0529_ ;
wire \us33/_0530_ ;
wire \us33/_0531_ ;
wire \us33/_0532_ ;
wire \us33/_0533_ ;
wire \us33/_0534_ ;
wire \us33/_0535_ ;
wire \us33/_0536_ ;
wire \us33/_0537_ ;
wire \us33/_0538_ ;
wire \us33/_0539_ ;
wire \us33/_0540_ ;
wire \us33/_0541_ ;
wire \us33/_0542_ ;
wire \us33/_0544_ ;
wire \us33/_0545_ ;
wire \us33/_0546_ ;
wire \us33/_0547_ ;
wire \us33/_0548_ ;
wire \us33/_0549_ ;
wire \us33/_0550_ ;
wire \us33/_0551_ ;
wire \us33/_0552_ ;
wire \us33/_0553_ ;
wire \us33/_0554_ ;
wire \us33/_0555_ ;
wire \us33/_0556_ ;
wire \us33/_0557_ ;
wire \us33/_0558_ ;
wire \us33/_0559_ ;
wire \us33/_0560_ ;
wire \us33/_0561_ ;
wire \us33/_0562_ ;
wire \us33/_0563_ ;
wire \us33/_0565_ ;
wire \us33/_0566_ ;
wire \us33/_0567_ ;
wire \us33/_0568_ ;
wire \us33/_0569_ ;
wire \us33/_0570_ ;
wire \us33/_0571_ ;
wire \us33/_0572_ ;
wire \us33/_0573_ ;
wire \us33/_0574_ ;
wire \us33/_0575_ ;
wire \us33/_0576_ ;
wire \us33/_0577_ ;
wire \us33/_0578_ ;
wire \us33/_0579_ ;
wire \us33/_0580_ ;
wire \us33/_0581_ ;
wire \us33/_0582_ ;
wire \us33/_0583_ ;
wire \us33/_0584_ ;
wire \us33/_0585_ ;
wire \us33/_0586_ ;
wire \us33/_0587_ ;
wire \us33/_0588_ ;
wire \us33/_0589_ ;
wire \us33/_0590_ ;
wire \us33/_0591_ ;
wire \us33/_0592_ ;
wire \us33/_0593_ ;
wire \us33/_0594_ ;
wire \us33/_0595_ ;
wire \us33/_0596_ ;
wire \us33/_0598_ ;
wire \us33/_0599_ ;
wire \us33/_0600_ ;
wire \us33/_0601_ ;
wire \us33/_0602_ ;
wire \us33/_0603_ ;
wire \us33/_0604_ ;
wire \us33/_0605_ ;
wire \us33/_0606_ ;
wire \us33/_0607_ ;
wire \us33/_0608_ ;
wire \us33/_0609_ ;
wire \us33/_0610_ ;
wire \us33/_0611_ ;
wire \us33/_0612_ ;
wire \us33/_0613_ ;
wire \us33/_0614_ ;
wire \us33/_0615_ ;
wire \us33/_0616_ ;
wire \us33/_0617_ ;
wire \us33/_0618_ ;
wire \us33/_0619_ ;
wire \us33/_0620_ ;
wire \us33/_0621_ ;
wire \us33/_0622_ ;
wire \us33/_0623_ ;
wire \us33/_0624_ ;
wire \us33/_0625_ ;
wire \us33/_0626_ ;
wire \us33/_0627_ ;
wire \us33/_0628_ ;
wire \us33/_0629_ ;
wire \us33/_0630_ ;
wire \us33/_0631_ ;
wire \us33/_0632_ ;
wire \us33/_0633_ ;
wire \us33/_0634_ ;
wire \us33/_0635_ ;
wire \us33/_0636_ ;
wire \us33/_0637_ ;
wire \us33/_0638_ ;
wire \us33/_0639_ ;
wire \us33/_0640_ ;
wire \us33/_0641_ ;
wire \us33/_0642_ ;
wire \us33/_0643_ ;
wire \us33/_0644_ ;
wire \us33/_0645_ ;
wire \us33/_0646_ ;
wire \us33/_0647_ ;
wire \us33/_0648_ ;
wire \us33/_0649_ ;
wire \us33/_0650_ ;
wire \us33/_0652_ ;
wire \us33/_0653_ ;
wire \us33/_0654_ ;
wire \us33/_0655_ ;
wire \us33/_0656_ ;
wire \us33/_0657_ ;
wire \us33/_0658_ ;
wire \us33/_0659_ ;
wire \us33/_0660_ ;
wire \us33/_0661_ ;
wire \us33/_0662_ ;
wire \us33/_0663_ ;
wire \us33/_0664_ ;
wire \us33/_0665_ ;
wire \us33/_0666_ ;
wire \us33/_0667_ ;
wire \us33/_0668_ ;
wire \us33/_0669_ ;
wire \us33/_0670_ ;
wire \us33/_0671_ ;
wire \us33/_0673_ ;
wire \us33/_0674_ ;
wire \us33/_0675_ ;
wire \us33/_0676_ ;
wire \us33/_0677_ ;
wire \us33/_0678_ ;
wire \us33/_0679_ ;
wire \us33/_0680_ ;
wire \us33/_0681_ ;
wire \us33/_0682_ ;
wire \us33/_0683_ ;
wire \us33/_0684_ ;
wire \us33/_0685_ ;
wire \us33/_0686_ ;
wire \us33/_0687_ ;
wire \us33/_0688_ ;
wire \us33/_0689_ ;
wire \us33/_0690_ ;
wire \us33/_0691_ ;
wire \us33/_0692_ ;
wire \us33/_0693_ ;
wire \us33/_0694_ ;
wire \us33/_0695_ ;
wire \us33/_0696_ ;
wire \us33/_0697_ ;
wire \us33/_0698_ ;
wire \us33/_0699_ ;
wire \us33/_0700_ ;
wire \us33/_0701_ ;
wire \us33/_0702_ ;
wire \us33/_0703_ ;
wire \us33/_0704_ ;
wire \us33/_0705_ ;
wire \us33/_0706_ ;
wire \us33/_0707_ ;
wire \us33/_0708_ ;
wire \us33/_0709_ ;
wire \us33/_0710_ ;
wire \us33/_0711_ ;
wire \us33/_0712_ ;
wire \us33/_0713_ ;
wire \us33/_0714_ ;
wire \us33/_0715_ ;
wire \us33/_0717_ ;
wire \us33/_0718_ ;
wire \us33/_0719_ ;
wire \us33/_0720_ ;
wire \us33/_0721_ ;
wire \us33/_0722_ ;
wire \us33/_0723_ ;
wire \us33/_0724_ ;
wire \us33/_0725_ ;
wire \us33/_0726_ ;
wire \us33/_0727_ ;
wire \us33/_0728_ ;
wire \us33/_0729_ ;
wire \us33/_0730_ ;
wire \us33/_0731_ ;
wire \us33/_0733_ ;
wire \us33/_0734_ ;
wire \us33/_0735_ ;
wire \us33/_0736_ ;
wire \us33/_0738_ ;
wire \us33/_0739_ ;
wire \us33/_0740_ ;
wire \us33/_0741_ ;
wire \us33/_0742_ ;
wire \us33/_0744_ ;
wire \us33/_0745_ ;
wire \us33/_0746_ ;
wire \us33/_0748_ ;
wire \us33/_0749_ ;
wire \us33/_0750_ ;
wire \us33/_0752_ ;
wire \w0[0] ;
wire \w0[10] ;
wire \w0[11] ;
wire \w0[12] ;
wire \w0[13] ;
wire \w0[14] ;
wire \w0[15] ;
wire \w0[16] ;
wire \w0[17] ;
wire \w0[18] ;
wire \w0[19] ;
wire \w0[1] ;
wire \w0[20] ;
wire \w0[21] ;
wire \w0[22] ;
wire \w0[23] ;
wire \w0[24] ;
wire \w0[25] ;
wire \w0[26] ;
wire \w0[27] ;
wire \w0[28] ;
wire \w0[29] ;
wire \w0[2] ;
wire \w0[30] ;
wire \w0[31] ;
wire \w0[3] ;
wire \w0[4] ;
wire \w0[5] ;
wire \w0[6] ;
wire \w0[7] ;
wire \w0[8] ;
wire \w0[9] ;
wire \w1[0] ;
wire \w1[10] ;
wire \w1[11] ;
wire \w1[12] ;
wire \w1[13] ;
wire \w1[14] ;
wire \w1[15] ;
wire \w1[16] ;
wire \w1[17] ;
wire \w1[18] ;
wire \w1[19] ;
wire \w1[1] ;
wire \w1[20] ;
wire \w1[21] ;
wire \w1[22] ;
wire \w1[23] ;
wire \w1[24] ;
wire \w1[25] ;
wire \w1[26] ;
wire \w1[27] ;
wire \w1[28] ;
wire \w1[29] ;
wire \w1[2] ;
wire \w1[30] ;
wire \w1[31] ;
wire \w1[3] ;
wire \w1[4] ;
wire \w1[5] ;
wire \w1[6] ;
wire \w1[7] ;
wire \w1[8] ;
wire \w1[9] ;
wire \w2[0] ;
wire \w2[10] ;
wire \w2[11] ;
wire \w2[12] ;
wire \w2[13] ;
wire \w2[14] ;
wire \w2[15] ;
wire \w2[16] ;
wire \w2[17] ;
wire \w2[18] ;
wire \w2[19] ;
wire \w2[1] ;
wire \w2[20] ;
wire \w2[21] ;
wire \w2[22] ;
wire \w2[23] ;
wire \w2[24] ;
wire \w2[25] ;
wire \w2[26] ;
wire \w2[27] ;
wire \w2[28] ;
wire \w2[29] ;
wire \w2[2] ;
wire \w2[30] ;
wire \w2[31] ;
wire \w2[3] ;
wire \w2[4] ;
wire \w2[5] ;
wire \w2[6] ;
wire \w2[7] ;
wire \w2[8] ;
wire \w2[9] ;
wire \w3[0] ;
wire \w3[10] ;
wire \w3[11] ;
wire \w3[12] ;
wire \w3[13] ;
wire \w3[14] ;
wire \w3[15] ;
wire \w3[16] ;
wire \w3[17] ;
wire \w3[18] ;
wire \w3[19] ;
wire \w3[1] ;
wire \w3[20] ;
wire \w3[21] ;
wire \w3[22] ;
wire \w3[23] ;
wire \w3[24] ;
wire \w3[25] ;
wire \w3[26] ;
wire \w3[27] ;
wire \w3[28] ;
wire \w3[29] ;
wire \w3[2] ;
wire \w3[30] ;
wire \w3[31] ;
wire \w3[3] ;
wire \w3[4] ;
wire \w3[5] ;
wire \w3[6] ;
wire \w3[7] ;
wire \w3[8] ;
wire \w3[9] ;
wire [127:0] key ;
wire [127:0] text_in ;
wire [127:0] text_out ;

sky130_fd_sc_hd__clkbuf_4 FE_OFC0_text_out_80 ( .A(FE_OFN0_text_out_80 ), .X(\text_out[80] ) );
sky130_fd_sc_hd__clkinv_8 CTS_ccl_a_inv_00081 ( .A(CTS_19 ), .Y(CTS_18 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00069 ( .A(CTS_19 ), .Y(CTS_21 ) );
sky130_fd_sc_hd__clkinv_8 CTS_ccl_a_inv_00065 ( .A(CTS_19 ), .Y(CTS_20 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00106 ( .A(CTS_22 ), .Y(CTS_19 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00083 ( .A(CTS_15 ), .Y(CTS_14 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00079 ( .A(CTS_15 ), .Y(CTS_17 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00077 ( .A(CTS_15 ), .Y(CTS_16 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00104 ( .A(CTS_22 ), .Y(CTS_15 ) );
sky130_fd_sc_hd__clkinv_8 CTS_ccl_a_inv_00113 ( .A(CTS_23 ), .Y(CTS_22 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00067 ( .A(CTS_10 ), .Y(CTS_9 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00059 ( .A(CTS_10 ), .Y(CTS_12 ) );
sky130_fd_sc_hd__clkinv_2 CTS_ccl_a_inv_00057 ( .A(CTS_10 ), .Y(CTS_11 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00102 ( .A(CTS_13 ), .Y(CTS_10 ) );
sky130_fd_sc_hd__clkinv_4 CTS_ccl_a_inv_00073 ( .A(CTS_6 ), .Y(CTS_5 ) );
sky130_fd_sc_hd__clkinv_8 CTS_ccl_a_inv_00071 ( .A(CTS_6 ), .Y(CTS_8 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00061 ( .A(CTS_6 ), .Y(CTS_7 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00100 ( .A(CTS_13 ), .Y(CTS_6 ) );
sky130_fd_sc_hd__clkinv_8 CTS_ccl_a_inv_00075 ( .A(CTS_2 ), .Y(CTS_1 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00063 ( .A(CTS_2 ), .Y(CTS_4 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00055 ( .A(CTS_2 ), .Y(CTS_3 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00098 ( .A(CTS_13 ), .Y(CTS_2 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00111 ( .A(CTS_23 ), .Y(CTS_13 ) );
sky130_fd_sc_hd__clkinv_16 CTS_ccl_a_inv_00118 ( .A(clk ), .Y(CTS_23 ) );
sky130_fd_sc_hd__fill_1 PHY_0 (  );
sky130_fd_sc_hd__fill_1 PHY_1 (  );
sky130_fd_sc_hd__fill_1 PHY_10 (  );
sky130_fd_sc_hd__fill_1 PHY_100 (  );
sky130_fd_sc_hd__fill_1 PHY_101 (  );
sky130_fd_sc_hd__fill_1 PHY_102 (  );
sky130_fd_sc_hd__fill_1 PHY_103 (  );
sky130_fd_sc_hd__fill_1 PHY_104 (  );
sky130_fd_sc_hd__fill_1 PHY_105 (  );
sky130_fd_sc_hd__fill_1 PHY_106 (  );
sky130_fd_sc_hd__fill_1 PHY_107 (  );
sky130_fd_sc_hd__fill_1 PHY_108 (  );
sky130_fd_sc_hd__fill_1 PHY_109 (  );
sky130_fd_sc_hd__fill_1 PHY_11 (  );
sky130_fd_sc_hd__fill_1 PHY_110 (  );
sky130_fd_sc_hd__fill_1 PHY_111 (  );
sky130_fd_sc_hd__fill_1 PHY_112 (  );
sky130_fd_sc_hd__fill_1 PHY_113 (  );
sky130_fd_sc_hd__fill_1 PHY_114 (  );
sky130_fd_sc_hd__fill_1 PHY_115 (  );
sky130_fd_sc_hd__fill_1 PHY_116 (  );
sky130_fd_sc_hd__fill_1 PHY_117 (  );
sky130_fd_sc_hd__fill_1 PHY_118 (  );
sky130_fd_sc_hd__fill_1 PHY_119 (  );
sky130_fd_sc_hd__fill_1 PHY_12 (  );
sky130_fd_sc_hd__fill_1 PHY_120 (  );
sky130_fd_sc_hd__fill_1 PHY_121 (  );
sky130_fd_sc_hd__fill_1 PHY_122 (  );
sky130_fd_sc_hd__fill_1 PHY_123 (  );
sky130_fd_sc_hd__fill_1 PHY_124 (  );
sky130_fd_sc_hd__fill_1 PHY_125 (  );
sky130_fd_sc_hd__fill_1 PHY_126 (  );
sky130_fd_sc_hd__fill_1 PHY_127 (  );
sky130_fd_sc_hd__fill_1 PHY_128 (  );
sky130_fd_sc_hd__fill_1 PHY_129 (  );
sky130_fd_sc_hd__fill_1 PHY_13 (  );
sky130_fd_sc_hd__fill_1 PHY_130 (  );
sky130_fd_sc_hd__fill_1 PHY_131 (  );
sky130_fd_sc_hd__fill_1 PHY_132 (  );
sky130_fd_sc_hd__fill_1 PHY_133 (  );
sky130_fd_sc_hd__fill_1 PHY_134 (  );
sky130_fd_sc_hd__fill_1 PHY_135 (  );
sky130_fd_sc_hd__fill_1 PHY_136 (  );
sky130_fd_sc_hd__fill_1 PHY_137 (  );
sky130_fd_sc_hd__fill_1 PHY_138 (  );
sky130_fd_sc_hd__fill_1 PHY_139 (  );
sky130_fd_sc_hd__fill_1 PHY_14 (  );
sky130_fd_sc_hd__fill_1 PHY_140 (  );
sky130_fd_sc_hd__fill_1 PHY_141 (  );
sky130_fd_sc_hd__fill_1 PHY_142 (  );
sky130_fd_sc_hd__fill_1 PHY_143 (  );
sky130_fd_sc_hd__fill_1 PHY_144 (  );
sky130_fd_sc_hd__fill_1 PHY_145 (  );
sky130_fd_sc_hd__fill_1 PHY_146 (  );
sky130_fd_sc_hd__fill_1 PHY_147 (  );
sky130_fd_sc_hd__fill_1 PHY_148 (  );
sky130_fd_sc_hd__fill_1 PHY_149 (  );
sky130_fd_sc_hd__fill_1 PHY_15 (  );
sky130_fd_sc_hd__fill_1 PHY_150 (  );
sky130_fd_sc_hd__fill_1 PHY_151 (  );
sky130_fd_sc_hd__fill_1 PHY_152 (  );
sky130_fd_sc_hd__fill_1 PHY_153 (  );
sky130_fd_sc_hd__fill_1 PHY_154 (  );
sky130_fd_sc_hd__fill_1 PHY_155 (  );
sky130_fd_sc_hd__fill_1 PHY_156 (  );
sky130_fd_sc_hd__fill_1 PHY_157 (  );
sky130_fd_sc_hd__fill_1 PHY_158 (  );
sky130_fd_sc_hd__fill_1 PHY_159 (  );
sky130_fd_sc_hd__fill_1 PHY_16 (  );
sky130_fd_sc_hd__fill_1 PHY_160 (  );
sky130_fd_sc_hd__fill_1 PHY_161 (  );
sky130_fd_sc_hd__fill_1 PHY_162 (  );
sky130_fd_sc_hd__fill_1 PHY_163 (  );
sky130_fd_sc_hd__fill_1 PHY_164 (  );
sky130_fd_sc_hd__fill_1 PHY_165 (  );
sky130_fd_sc_hd__fill_1 PHY_166 (  );
sky130_fd_sc_hd__fill_1 PHY_167 (  );
sky130_fd_sc_hd__fill_1 PHY_168 (  );
sky130_fd_sc_hd__fill_1 PHY_169 (  );
sky130_fd_sc_hd__fill_1 PHY_17 (  );
sky130_fd_sc_hd__fill_1 PHY_170 (  );
sky130_fd_sc_hd__fill_1 PHY_171 (  );
sky130_fd_sc_hd__fill_1 PHY_172 (  );
sky130_fd_sc_hd__fill_1 PHY_173 (  );
sky130_fd_sc_hd__fill_1 PHY_174 (  );
sky130_fd_sc_hd__fill_1 PHY_175 (  );
sky130_fd_sc_hd__fill_1 PHY_176 (  );
sky130_fd_sc_hd__fill_1 PHY_177 (  );
sky130_fd_sc_hd__fill_1 PHY_178 (  );
sky130_fd_sc_hd__fill_1 PHY_179 (  );
sky130_fd_sc_hd__fill_1 PHY_18 (  );
sky130_fd_sc_hd__fill_1 PHY_180 (  );
sky130_fd_sc_hd__fill_1 PHY_181 (  );
sky130_fd_sc_hd__fill_1 PHY_182 (  );
sky130_fd_sc_hd__fill_1 PHY_183 (  );
sky130_fd_sc_hd__fill_1 PHY_184 (  );
sky130_fd_sc_hd__fill_1 PHY_185 (  );
sky130_fd_sc_hd__fill_1 PHY_186 (  );
sky130_fd_sc_hd__fill_1 PHY_187 (  );
sky130_fd_sc_hd__fill_1 PHY_188 (  );
sky130_fd_sc_hd__fill_1 PHY_189 (  );
sky130_fd_sc_hd__fill_1 PHY_19 (  );
sky130_fd_sc_hd__fill_1 PHY_190 (  );
sky130_fd_sc_hd__fill_1 PHY_191 (  );
sky130_fd_sc_hd__fill_1 PHY_192 (  );
sky130_fd_sc_hd__fill_1 PHY_193 (  );
sky130_fd_sc_hd__fill_1 PHY_194 (  );
sky130_fd_sc_hd__fill_1 PHY_195 (  );
sky130_fd_sc_hd__fill_1 PHY_196 (  );
sky130_fd_sc_hd__fill_1 PHY_197 (  );
sky130_fd_sc_hd__fill_1 PHY_198 (  );
sky130_fd_sc_hd__fill_1 PHY_199 (  );
sky130_fd_sc_hd__fill_1 PHY_2 (  );
sky130_fd_sc_hd__fill_1 PHY_20 (  );
sky130_fd_sc_hd__fill_1 PHY_200 (  );
sky130_fd_sc_hd__fill_1 PHY_201 (  );
sky130_fd_sc_hd__fill_1 PHY_202 (  );
sky130_fd_sc_hd__fill_1 PHY_203 (  );
sky130_fd_sc_hd__fill_1 PHY_204 (  );
sky130_fd_sc_hd__fill_1 PHY_205 (  );
sky130_fd_sc_hd__fill_1 PHY_206 (  );
sky130_fd_sc_hd__fill_1 PHY_207 (  );
sky130_fd_sc_hd__fill_1 PHY_208 (  );
sky130_fd_sc_hd__fill_1 PHY_209 (  );
sky130_fd_sc_hd__fill_1 PHY_21 (  );
sky130_fd_sc_hd__fill_1 PHY_210 (  );
sky130_fd_sc_hd__fill_1 PHY_211 (  );
sky130_fd_sc_hd__fill_1 PHY_212 (  );
sky130_fd_sc_hd__fill_1 PHY_213 (  );
sky130_fd_sc_hd__fill_1 PHY_214 (  );
sky130_fd_sc_hd__fill_1 PHY_215 (  );
sky130_fd_sc_hd__fill_1 PHY_216 (  );
sky130_fd_sc_hd__fill_1 PHY_217 (  );
sky130_fd_sc_hd__fill_1 PHY_218 (  );
sky130_fd_sc_hd__fill_1 PHY_219 (  );
sky130_fd_sc_hd__fill_1 PHY_22 (  );
sky130_fd_sc_hd__fill_1 PHY_220 (  );
sky130_fd_sc_hd__fill_1 PHY_221 (  );
sky130_fd_sc_hd__fill_1 PHY_222 (  );
sky130_fd_sc_hd__fill_1 PHY_223 (  );
sky130_fd_sc_hd__fill_1 PHY_224 (  );
sky130_fd_sc_hd__fill_1 PHY_225 (  );
sky130_fd_sc_hd__fill_1 PHY_226 (  );
sky130_fd_sc_hd__fill_1 PHY_227 (  );
sky130_fd_sc_hd__fill_1 PHY_228 (  );
sky130_fd_sc_hd__fill_1 PHY_229 (  );
sky130_fd_sc_hd__fill_1 PHY_23 (  );
sky130_fd_sc_hd__fill_1 PHY_230 (  );
sky130_fd_sc_hd__fill_1 PHY_231 (  );
sky130_fd_sc_hd__fill_1 PHY_232 (  );
sky130_fd_sc_hd__fill_1 PHY_233 (  );
sky130_fd_sc_hd__fill_1 PHY_234 (  );
sky130_fd_sc_hd__fill_1 PHY_235 (  );
sky130_fd_sc_hd__fill_1 PHY_236 (  );
sky130_fd_sc_hd__fill_1 PHY_237 (  );
sky130_fd_sc_hd__fill_1 PHY_238 (  );
sky130_fd_sc_hd__fill_1 PHY_239 (  );
sky130_fd_sc_hd__fill_1 PHY_24 (  );
sky130_fd_sc_hd__fill_1 PHY_240 (  );
sky130_fd_sc_hd__fill_1 PHY_241 (  );
sky130_fd_sc_hd__fill_1 PHY_242 (  );
sky130_fd_sc_hd__fill_1 PHY_243 (  );
sky130_fd_sc_hd__fill_1 PHY_244 (  );
sky130_fd_sc_hd__fill_1 PHY_245 (  );
sky130_fd_sc_hd__fill_1 PHY_246 (  );
sky130_fd_sc_hd__fill_1 PHY_247 (  );
sky130_fd_sc_hd__fill_1 PHY_248 (  );
sky130_fd_sc_hd__fill_1 PHY_249 (  );
sky130_fd_sc_hd__fill_1 PHY_25 (  );
sky130_fd_sc_hd__fill_1 PHY_250 (  );
sky130_fd_sc_hd__fill_1 PHY_251 (  );
sky130_fd_sc_hd__fill_1 PHY_252 (  );
sky130_fd_sc_hd__fill_1 PHY_253 (  );
sky130_fd_sc_hd__fill_1 PHY_254 (  );
sky130_fd_sc_hd__fill_1 PHY_255 (  );
sky130_fd_sc_hd__fill_1 PHY_256 (  );
sky130_fd_sc_hd__fill_1 PHY_257 (  );
sky130_fd_sc_hd__fill_1 PHY_258 (  );
sky130_fd_sc_hd__fill_1 PHY_259 (  );
sky130_fd_sc_hd__fill_1 PHY_26 (  );
sky130_fd_sc_hd__fill_1 PHY_260 (  );
sky130_fd_sc_hd__fill_1 PHY_261 (  );
sky130_fd_sc_hd__fill_1 PHY_262 (  );
sky130_fd_sc_hd__fill_1 PHY_263 (  );
sky130_fd_sc_hd__fill_1 PHY_264 (  );
sky130_fd_sc_hd__fill_1 PHY_265 (  );
sky130_fd_sc_hd__fill_1 PHY_266 (  );
sky130_fd_sc_hd__fill_1 PHY_267 (  );
sky130_fd_sc_hd__fill_1 PHY_268 (  );
sky130_fd_sc_hd__fill_1 PHY_269 (  );
sky130_fd_sc_hd__fill_1 PHY_27 (  );
sky130_fd_sc_hd__fill_1 PHY_270 (  );
sky130_fd_sc_hd__fill_1 PHY_271 (  );
sky130_fd_sc_hd__fill_1 PHY_272 (  );
sky130_fd_sc_hd__fill_1 PHY_273 (  );
sky130_fd_sc_hd__fill_1 PHY_274 (  );
sky130_fd_sc_hd__fill_1 PHY_275 (  );
sky130_fd_sc_hd__fill_1 PHY_276 (  );
sky130_fd_sc_hd__fill_1 PHY_277 (  );
sky130_fd_sc_hd__fill_1 PHY_278 (  );
sky130_fd_sc_hd__fill_1 PHY_279 (  );
sky130_fd_sc_hd__fill_1 PHY_28 (  );
sky130_fd_sc_hd__fill_1 PHY_280 (  );
sky130_fd_sc_hd__fill_1 PHY_281 (  );
sky130_fd_sc_hd__fill_1 PHY_282 (  );
sky130_fd_sc_hd__fill_1 PHY_283 (  );
sky130_fd_sc_hd__fill_1 PHY_284 (  );
sky130_fd_sc_hd__fill_1 PHY_285 (  );
sky130_fd_sc_hd__fill_1 PHY_286 (  );
sky130_fd_sc_hd__fill_1 PHY_287 (  );
sky130_fd_sc_hd__fill_1 PHY_288 (  );
sky130_fd_sc_hd__fill_1 PHY_289 (  );
sky130_fd_sc_hd__fill_1 PHY_29 (  );
sky130_fd_sc_hd__fill_1 PHY_290 (  );
sky130_fd_sc_hd__fill_1 PHY_291 (  );
sky130_fd_sc_hd__fill_1 PHY_292 (  );
sky130_fd_sc_hd__fill_1 PHY_293 (  );
sky130_fd_sc_hd__fill_1 PHY_294 (  );
sky130_fd_sc_hd__fill_1 PHY_295 (  );
sky130_fd_sc_hd__fill_1 PHY_296 (  );
sky130_fd_sc_hd__fill_1 PHY_297 (  );
sky130_fd_sc_hd__fill_1 PHY_298 (  );
sky130_fd_sc_hd__fill_1 PHY_299 (  );
sky130_fd_sc_hd__fill_1 PHY_3 (  );
sky130_fd_sc_hd__fill_1 PHY_30 (  );
sky130_fd_sc_hd__fill_1 PHY_300 (  );
sky130_fd_sc_hd__fill_1 PHY_301 (  );
sky130_fd_sc_hd__fill_1 PHY_302 (  );
sky130_fd_sc_hd__fill_1 PHY_303 (  );
sky130_fd_sc_hd__fill_1 PHY_304 (  );
sky130_fd_sc_hd__fill_1 PHY_305 (  );
sky130_fd_sc_hd__fill_1 PHY_306 (  );
sky130_fd_sc_hd__fill_1 PHY_307 (  );
sky130_fd_sc_hd__fill_1 PHY_308 (  );
sky130_fd_sc_hd__fill_1 PHY_309 (  );
sky130_fd_sc_hd__fill_1 PHY_31 (  );
sky130_fd_sc_hd__fill_1 PHY_310 (  );
sky130_fd_sc_hd__fill_1 PHY_311 (  );
sky130_fd_sc_hd__fill_1 PHY_312 (  );
sky130_fd_sc_hd__fill_1 PHY_313 (  );
sky130_fd_sc_hd__fill_1 PHY_314 (  );
sky130_fd_sc_hd__fill_1 PHY_315 (  );
sky130_fd_sc_hd__fill_1 PHY_316 (  );
sky130_fd_sc_hd__fill_1 PHY_317 (  );
sky130_fd_sc_hd__fill_1 PHY_318 (  );
sky130_fd_sc_hd__fill_1 PHY_319 (  );
sky130_fd_sc_hd__fill_1 PHY_32 (  );
sky130_fd_sc_hd__fill_1 PHY_320 (  );
sky130_fd_sc_hd__fill_1 PHY_321 (  );
sky130_fd_sc_hd__fill_1 PHY_322 (  );
sky130_fd_sc_hd__fill_1 PHY_323 (  );
sky130_fd_sc_hd__fill_1 PHY_324 (  );
sky130_fd_sc_hd__fill_1 PHY_325 (  );
sky130_fd_sc_hd__fill_1 PHY_326 (  );
sky130_fd_sc_hd__fill_1 PHY_327 (  );
sky130_fd_sc_hd__fill_1 PHY_328 (  );
sky130_fd_sc_hd__fill_1 PHY_329 (  );
sky130_fd_sc_hd__fill_1 PHY_33 (  );
sky130_fd_sc_hd__fill_1 PHY_330 (  );
sky130_fd_sc_hd__fill_1 PHY_331 (  );
sky130_fd_sc_hd__fill_1 PHY_332 (  );
sky130_fd_sc_hd__fill_1 PHY_333 (  );
sky130_fd_sc_hd__fill_1 PHY_334 (  );
sky130_fd_sc_hd__fill_1 PHY_335 (  );
sky130_fd_sc_hd__fill_1 PHY_336 (  );
sky130_fd_sc_hd__fill_1 PHY_337 (  );
sky130_fd_sc_hd__fill_1 PHY_338 (  );
sky130_fd_sc_hd__fill_1 PHY_339 (  );
sky130_fd_sc_hd__fill_1 PHY_34 (  );
sky130_fd_sc_hd__fill_1 PHY_340 (  );
sky130_fd_sc_hd__fill_1 PHY_341 (  );
sky130_fd_sc_hd__fill_1 PHY_342 (  );
sky130_fd_sc_hd__fill_1 PHY_343 (  );
sky130_fd_sc_hd__fill_1 PHY_344 (  );
sky130_fd_sc_hd__fill_1 PHY_345 (  );
sky130_fd_sc_hd__fill_1 PHY_346 (  );
sky130_fd_sc_hd__fill_1 PHY_347 (  );
sky130_fd_sc_hd__fill_1 PHY_348 (  );
sky130_fd_sc_hd__fill_1 PHY_349 (  );
sky130_fd_sc_hd__fill_1 PHY_35 (  );
sky130_fd_sc_hd__fill_1 PHY_350 (  );
sky130_fd_sc_hd__fill_1 PHY_351 (  );
sky130_fd_sc_hd__fill_1 PHY_352 (  );
sky130_fd_sc_hd__fill_1 PHY_353 (  );
sky130_fd_sc_hd__fill_1 PHY_354 (  );
sky130_fd_sc_hd__fill_1 PHY_355 (  );
sky130_fd_sc_hd__fill_1 PHY_356 (  );
sky130_fd_sc_hd__fill_1 PHY_357 (  );
sky130_fd_sc_hd__fill_1 PHY_358 (  );
sky130_fd_sc_hd__fill_1 PHY_359 (  );
sky130_fd_sc_hd__fill_1 PHY_36 (  );
sky130_fd_sc_hd__fill_1 PHY_360 (  );
sky130_fd_sc_hd__fill_1 PHY_361 (  );
sky130_fd_sc_hd__fill_1 PHY_362 (  );
sky130_fd_sc_hd__fill_1 PHY_363 (  );
sky130_fd_sc_hd__fill_1 PHY_364 (  );
sky130_fd_sc_hd__fill_1 PHY_365 (  );
sky130_fd_sc_hd__fill_1 PHY_366 (  );
sky130_fd_sc_hd__fill_1 PHY_367 (  );
sky130_fd_sc_hd__fill_1 PHY_368 (  );
sky130_fd_sc_hd__fill_1 PHY_369 (  );
sky130_fd_sc_hd__fill_1 PHY_37 (  );
sky130_fd_sc_hd__fill_1 PHY_370 (  );
sky130_fd_sc_hd__fill_1 PHY_371 (  );
sky130_fd_sc_hd__fill_1 PHY_372 (  );
sky130_fd_sc_hd__fill_1 PHY_373 (  );
sky130_fd_sc_hd__fill_1 PHY_374 (  );
sky130_fd_sc_hd__fill_1 PHY_375 (  );
sky130_fd_sc_hd__fill_1 PHY_376 (  );
sky130_fd_sc_hd__fill_1 PHY_377 (  );
sky130_fd_sc_hd__fill_1 PHY_378 (  );
sky130_fd_sc_hd__fill_1 PHY_379 (  );
sky130_fd_sc_hd__fill_1 PHY_38 (  );
sky130_fd_sc_hd__fill_1 PHY_380 (  );
sky130_fd_sc_hd__fill_1 PHY_381 (  );
sky130_fd_sc_hd__fill_1 PHY_382 (  );
sky130_fd_sc_hd__fill_1 PHY_383 (  );
sky130_fd_sc_hd__fill_1 PHY_384 (  );
sky130_fd_sc_hd__fill_1 PHY_385 (  );
sky130_fd_sc_hd__fill_1 PHY_386 (  );
sky130_fd_sc_hd__fill_1 PHY_387 (  );
sky130_fd_sc_hd__fill_1 PHY_388 (  );
sky130_fd_sc_hd__fill_1 PHY_389 (  );
sky130_fd_sc_hd__fill_1 PHY_39 (  );
sky130_fd_sc_hd__fill_1 PHY_390 (  );
sky130_fd_sc_hd__fill_1 PHY_391 (  );
sky130_fd_sc_hd__fill_1 PHY_392 (  );
sky130_fd_sc_hd__fill_1 PHY_393 (  );
sky130_fd_sc_hd__fill_1 PHY_394 (  );
sky130_fd_sc_hd__fill_1 PHY_395 (  );
sky130_fd_sc_hd__fill_1 PHY_396 (  );
sky130_fd_sc_hd__fill_1 PHY_397 (  );
sky130_fd_sc_hd__fill_1 PHY_398 (  );
sky130_fd_sc_hd__fill_1 PHY_399 (  );
sky130_fd_sc_hd__fill_1 PHY_4 (  );
sky130_fd_sc_hd__fill_1 PHY_40 (  );
sky130_fd_sc_hd__fill_1 PHY_400 (  );
sky130_fd_sc_hd__fill_1 PHY_401 (  );
sky130_fd_sc_hd__fill_1 PHY_402 (  );
sky130_fd_sc_hd__fill_1 PHY_403 (  );
sky130_fd_sc_hd__fill_1 PHY_404 (  );
sky130_fd_sc_hd__fill_1 PHY_405 (  );
sky130_fd_sc_hd__fill_1 PHY_406 (  );
sky130_fd_sc_hd__fill_1 PHY_407 (  );
sky130_fd_sc_hd__fill_1 PHY_408 (  );
sky130_fd_sc_hd__fill_1 PHY_409 (  );
sky130_fd_sc_hd__fill_1 PHY_41 (  );
sky130_fd_sc_hd__fill_1 PHY_410 (  );
sky130_fd_sc_hd__fill_1 PHY_411 (  );
sky130_fd_sc_hd__fill_1 PHY_412 (  );
sky130_fd_sc_hd__fill_1 PHY_413 (  );
sky130_fd_sc_hd__fill_1 PHY_414 (  );
sky130_fd_sc_hd__fill_1 PHY_415 (  );
sky130_fd_sc_hd__fill_1 PHY_416 (  );
sky130_fd_sc_hd__fill_1 PHY_417 (  );
sky130_fd_sc_hd__fill_1 PHY_418 (  );
sky130_fd_sc_hd__fill_1 PHY_419 (  );
sky130_fd_sc_hd__fill_1 PHY_42 (  );
sky130_fd_sc_hd__fill_1 PHY_420 (  );
sky130_fd_sc_hd__fill_1 PHY_421 (  );
sky130_fd_sc_hd__fill_1 PHY_422 (  );
sky130_fd_sc_hd__fill_1 PHY_423 (  );
sky130_fd_sc_hd__fill_1 PHY_424 (  );
sky130_fd_sc_hd__fill_1 PHY_425 (  );
sky130_fd_sc_hd__fill_1 PHY_426 (  );
sky130_fd_sc_hd__fill_1 PHY_427 (  );
sky130_fd_sc_hd__fill_1 PHY_428 (  );
sky130_fd_sc_hd__fill_1 PHY_429 (  );
sky130_fd_sc_hd__fill_1 PHY_43 (  );
sky130_fd_sc_hd__fill_1 PHY_430 (  );
sky130_fd_sc_hd__fill_1 PHY_431 (  );
sky130_fd_sc_hd__fill_1 PHY_432 (  );
sky130_fd_sc_hd__fill_1 PHY_433 (  );
sky130_fd_sc_hd__fill_1 PHY_434 (  );
sky130_fd_sc_hd__fill_1 PHY_435 (  );
sky130_fd_sc_hd__fill_1 PHY_436 (  );
sky130_fd_sc_hd__fill_1 PHY_437 (  );
sky130_fd_sc_hd__fill_1 PHY_438 (  );
sky130_fd_sc_hd__fill_1 PHY_439 (  );
sky130_fd_sc_hd__fill_1 PHY_44 (  );
sky130_fd_sc_hd__fill_1 PHY_440 (  );
sky130_fd_sc_hd__fill_1 PHY_441 (  );
sky130_fd_sc_hd__fill_1 PHY_442 (  );
sky130_fd_sc_hd__fill_1 PHY_443 (  );
sky130_fd_sc_hd__fill_1 PHY_444 (  );
sky130_fd_sc_hd__fill_1 PHY_445 (  );
sky130_fd_sc_hd__fill_1 PHY_446 (  );
sky130_fd_sc_hd__fill_1 PHY_447 (  );
sky130_fd_sc_hd__fill_1 PHY_448 (  );
sky130_fd_sc_hd__fill_1 PHY_449 (  );
sky130_fd_sc_hd__fill_1 PHY_45 (  );
sky130_fd_sc_hd__fill_1 PHY_450 (  );
sky130_fd_sc_hd__fill_1 PHY_451 (  );
sky130_fd_sc_hd__fill_1 PHY_452 (  );
sky130_fd_sc_hd__fill_1 PHY_453 (  );
sky130_fd_sc_hd__fill_1 PHY_454 (  );
sky130_fd_sc_hd__fill_1 PHY_455 (  );
sky130_fd_sc_hd__fill_1 PHY_456 (  );
sky130_fd_sc_hd__fill_1 PHY_457 (  );
sky130_fd_sc_hd__fill_1 PHY_458 (  );
sky130_fd_sc_hd__fill_1 PHY_459 (  );
sky130_fd_sc_hd__fill_1 PHY_46 (  );
sky130_fd_sc_hd__fill_1 PHY_460 (  );
sky130_fd_sc_hd__fill_1 PHY_461 (  );
sky130_fd_sc_hd__fill_1 PHY_462 (  );
sky130_fd_sc_hd__fill_1 PHY_463 (  );
sky130_fd_sc_hd__fill_1 PHY_464 (  );
sky130_fd_sc_hd__fill_1 PHY_465 (  );
sky130_fd_sc_hd__fill_1 PHY_466 (  );
sky130_fd_sc_hd__fill_1 PHY_467 (  );
sky130_fd_sc_hd__fill_1 PHY_468 (  );
sky130_fd_sc_hd__fill_1 PHY_469 (  );
sky130_fd_sc_hd__fill_1 PHY_47 (  );
sky130_fd_sc_hd__fill_1 PHY_470 (  );
sky130_fd_sc_hd__fill_1 PHY_471 (  );
sky130_fd_sc_hd__fill_1 PHY_472 (  );
sky130_fd_sc_hd__fill_1 PHY_473 (  );
sky130_fd_sc_hd__fill_1 PHY_474 (  );
sky130_fd_sc_hd__fill_1 PHY_475 (  );
sky130_fd_sc_hd__fill_1 PHY_476 (  );
sky130_fd_sc_hd__fill_1 PHY_477 (  );
sky130_fd_sc_hd__fill_1 PHY_478 (  );
sky130_fd_sc_hd__fill_1 PHY_479 (  );
sky130_fd_sc_hd__fill_1 PHY_48 (  );
sky130_fd_sc_hd__fill_1 PHY_480 (  );
sky130_fd_sc_hd__fill_1 PHY_481 (  );
sky130_fd_sc_hd__fill_1 PHY_482 (  );
sky130_fd_sc_hd__fill_1 PHY_483 (  );
sky130_fd_sc_hd__fill_1 PHY_484 (  );
sky130_fd_sc_hd__fill_1 PHY_485 (  );
sky130_fd_sc_hd__fill_1 PHY_486 (  );
sky130_fd_sc_hd__fill_1 PHY_487 (  );
sky130_fd_sc_hd__fill_1 PHY_488 (  );
sky130_fd_sc_hd__fill_1 PHY_489 (  );
sky130_fd_sc_hd__fill_1 PHY_49 (  );
sky130_fd_sc_hd__fill_1 PHY_490 (  );
sky130_fd_sc_hd__fill_1 PHY_491 (  );
sky130_fd_sc_hd__fill_1 PHY_492 (  );
sky130_fd_sc_hd__fill_1 PHY_493 (  );
sky130_fd_sc_hd__fill_1 PHY_494 (  );
sky130_fd_sc_hd__fill_1 PHY_495 (  );
sky130_fd_sc_hd__fill_1 PHY_496 (  );
sky130_fd_sc_hd__fill_1 PHY_497 (  );
sky130_fd_sc_hd__fill_1 PHY_498 (  );
sky130_fd_sc_hd__fill_1 PHY_499 (  );
sky130_fd_sc_hd__fill_1 PHY_5 (  );
sky130_fd_sc_hd__fill_1 PHY_50 (  );
sky130_fd_sc_hd__fill_1 PHY_500 (  );
sky130_fd_sc_hd__fill_1 PHY_501 (  );
sky130_fd_sc_hd__fill_1 PHY_502 (  );
sky130_fd_sc_hd__fill_1 PHY_503 (  );
sky130_fd_sc_hd__fill_1 PHY_504 (  );
sky130_fd_sc_hd__fill_1 PHY_505 (  );
sky130_fd_sc_hd__fill_1 PHY_506 (  );
sky130_fd_sc_hd__fill_1 PHY_507 (  );
sky130_fd_sc_hd__fill_1 PHY_508 (  );
sky130_fd_sc_hd__fill_1 PHY_509 (  );
sky130_fd_sc_hd__fill_1 PHY_51 (  );
sky130_fd_sc_hd__fill_1 PHY_510 (  );
sky130_fd_sc_hd__fill_1 PHY_511 (  );
sky130_fd_sc_hd__fill_1 PHY_512 (  );
sky130_fd_sc_hd__fill_1 PHY_513 (  );
sky130_fd_sc_hd__fill_1 PHY_514 (  );
sky130_fd_sc_hd__fill_1 PHY_515 (  );
sky130_fd_sc_hd__fill_1 PHY_516 (  );
sky130_fd_sc_hd__fill_1 PHY_517 (  );
sky130_fd_sc_hd__fill_1 PHY_518 (  );
sky130_fd_sc_hd__fill_1 PHY_519 (  );
sky130_fd_sc_hd__fill_1 PHY_52 (  );
sky130_fd_sc_hd__fill_1 PHY_520 (  );
sky130_fd_sc_hd__fill_1 PHY_521 (  );
sky130_fd_sc_hd__fill_1 PHY_522 (  );
sky130_fd_sc_hd__fill_1 PHY_523 (  );
sky130_fd_sc_hd__fill_1 PHY_524 (  );
sky130_fd_sc_hd__fill_1 PHY_525 (  );
sky130_fd_sc_hd__fill_1 PHY_526 (  );
sky130_fd_sc_hd__fill_1 PHY_527 (  );
sky130_fd_sc_hd__fill_1 PHY_528 (  );
sky130_fd_sc_hd__fill_1 PHY_529 (  );
sky130_fd_sc_hd__fill_1 PHY_53 (  );
sky130_fd_sc_hd__fill_1 PHY_530 (  );
sky130_fd_sc_hd__fill_1 PHY_531 (  );
sky130_fd_sc_hd__fill_1 PHY_532 (  );
sky130_fd_sc_hd__fill_1 PHY_533 (  );
sky130_fd_sc_hd__fill_1 PHY_534 (  );
sky130_fd_sc_hd__fill_1 PHY_535 (  );
sky130_fd_sc_hd__fill_1 PHY_536 (  );
sky130_fd_sc_hd__fill_1 PHY_537 (  );
sky130_fd_sc_hd__fill_1 PHY_538 (  );
sky130_fd_sc_hd__fill_1 PHY_539 (  );
sky130_fd_sc_hd__fill_1 PHY_54 (  );
sky130_fd_sc_hd__fill_1 PHY_540 (  );
sky130_fd_sc_hd__fill_1 PHY_541 (  );
sky130_fd_sc_hd__fill_1 PHY_542 (  );
sky130_fd_sc_hd__fill_1 PHY_543 (  );
sky130_fd_sc_hd__fill_1 PHY_544 (  );
sky130_fd_sc_hd__fill_1 PHY_545 (  );
sky130_fd_sc_hd__fill_1 PHY_546 (  );
sky130_fd_sc_hd__fill_1 PHY_547 (  );
sky130_fd_sc_hd__fill_1 PHY_548 (  );
sky130_fd_sc_hd__fill_1 PHY_549 (  );
sky130_fd_sc_hd__fill_1 PHY_55 (  );
sky130_fd_sc_hd__fill_1 PHY_550 (  );
sky130_fd_sc_hd__fill_1 PHY_551 (  );
sky130_fd_sc_hd__fill_1 PHY_552 (  );
sky130_fd_sc_hd__fill_1 PHY_553 (  );
sky130_fd_sc_hd__fill_1 PHY_554 (  );
sky130_fd_sc_hd__fill_1 PHY_555 (  );
sky130_fd_sc_hd__fill_1 PHY_556 (  );
sky130_fd_sc_hd__fill_1 PHY_557 (  );
sky130_fd_sc_hd__fill_1 PHY_558 (  );
sky130_fd_sc_hd__fill_1 PHY_559 (  );
sky130_fd_sc_hd__fill_1 PHY_56 (  );
sky130_fd_sc_hd__fill_1 PHY_560 (  );
sky130_fd_sc_hd__fill_1 PHY_561 (  );
sky130_fd_sc_hd__fill_1 PHY_562 (  );
sky130_fd_sc_hd__fill_1 PHY_563 (  );
sky130_fd_sc_hd__fill_1 PHY_564 (  );
sky130_fd_sc_hd__fill_1 PHY_565 (  );
sky130_fd_sc_hd__fill_1 PHY_566 (  );
sky130_fd_sc_hd__fill_1 PHY_567 (  );
sky130_fd_sc_hd__fill_1 PHY_568 (  );
sky130_fd_sc_hd__fill_1 PHY_569 (  );
sky130_fd_sc_hd__fill_1 PHY_57 (  );
sky130_fd_sc_hd__fill_1 PHY_570 (  );
sky130_fd_sc_hd__fill_1 PHY_571 (  );
sky130_fd_sc_hd__fill_1 PHY_572 (  );
sky130_fd_sc_hd__fill_1 PHY_573 (  );
sky130_fd_sc_hd__fill_1 PHY_574 (  );
sky130_fd_sc_hd__fill_1 PHY_575 (  );
sky130_fd_sc_hd__fill_1 PHY_576 (  );
sky130_fd_sc_hd__fill_1 PHY_577 (  );
sky130_fd_sc_hd__fill_1 PHY_578 (  );
sky130_fd_sc_hd__fill_1 PHY_579 (  );
sky130_fd_sc_hd__fill_1 PHY_58 (  );
sky130_fd_sc_hd__fill_1 PHY_580 (  );
sky130_fd_sc_hd__fill_1 PHY_581 (  );
sky130_fd_sc_hd__fill_1 PHY_582 (  );
sky130_fd_sc_hd__fill_1 PHY_583 (  );
sky130_fd_sc_hd__fill_1 PHY_584 (  );
sky130_fd_sc_hd__fill_1 PHY_585 (  );
sky130_fd_sc_hd__fill_1 PHY_586 (  );
sky130_fd_sc_hd__fill_1 PHY_587 (  );
sky130_fd_sc_hd__fill_1 PHY_588 (  );
sky130_fd_sc_hd__fill_1 PHY_589 (  );
sky130_fd_sc_hd__fill_1 PHY_59 (  );
sky130_fd_sc_hd__fill_1 PHY_590 (  );
sky130_fd_sc_hd__fill_1 PHY_591 (  );
sky130_fd_sc_hd__fill_1 PHY_592 (  );
sky130_fd_sc_hd__fill_1 PHY_593 (  );
sky130_fd_sc_hd__fill_1 PHY_594 (  );
sky130_fd_sc_hd__fill_1 PHY_595 (  );
sky130_fd_sc_hd__fill_1 PHY_596 (  );
sky130_fd_sc_hd__fill_1 PHY_597 (  );
sky130_fd_sc_hd__fill_1 PHY_598 (  );
sky130_fd_sc_hd__fill_1 PHY_599 (  );
sky130_fd_sc_hd__fill_1 PHY_6 (  );
sky130_fd_sc_hd__fill_1 PHY_60 (  );
sky130_fd_sc_hd__fill_1 PHY_600 (  );
sky130_fd_sc_hd__fill_1 PHY_601 (  );
sky130_fd_sc_hd__fill_1 PHY_602 (  );
sky130_fd_sc_hd__fill_1 PHY_603 (  );
sky130_fd_sc_hd__fill_1 PHY_604 (  );
sky130_fd_sc_hd__fill_1 PHY_605 (  );
sky130_fd_sc_hd__fill_1 PHY_606 (  );
sky130_fd_sc_hd__fill_1 PHY_607 (  );
sky130_fd_sc_hd__fill_1 PHY_608 (  );
sky130_fd_sc_hd__fill_1 PHY_609 (  );
sky130_fd_sc_hd__fill_1 PHY_61 (  );
sky130_fd_sc_hd__fill_1 PHY_610 (  );
sky130_fd_sc_hd__fill_1 PHY_611 (  );
sky130_fd_sc_hd__fill_1 PHY_612 (  );
sky130_fd_sc_hd__fill_1 PHY_613 (  );
sky130_fd_sc_hd__fill_1 PHY_614 (  );
sky130_fd_sc_hd__fill_1 PHY_615 (  );
sky130_fd_sc_hd__fill_1 PHY_616 (  );
sky130_fd_sc_hd__fill_1 PHY_617 (  );
sky130_fd_sc_hd__fill_1 PHY_618 (  );
sky130_fd_sc_hd__fill_1 PHY_619 (  );
sky130_fd_sc_hd__fill_1 PHY_62 (  );
sky130_fd_sc_hd__fill_1 PHY_620 (  );
sky130_fd_sc_hd__fill_1 PHY_621 (  );
sky130_fd_sc_hd__fill_1 PHY_622 (  );
sky130_fd_sc_hd__fill_1 PHY_623 (  );
sky130_fd_sc_hd__fill_1 PHY_624 (  );
sky130_fd_sc_hd__fill_1 PHY_625 (  );
sky130_fd_sc_hd__fill_1 PHY_626 (  );
sky130_fd_sc_hd__fill_1 PHY_627 (  );
sky130_fd_sc_hd__fill_1 PHY_628 (  );
sky130_fd_sc_hd__fill_1 PHY_629 (  );
sky130_fd_sc_hd__fill_1 PHY_63 (  );
sky130_fd_sc_hd__fill_1 PHY_630 (  );
sky130_fd_sc_hd__fill_1 PHY_631 (  );
sky130_fd_sc_hd__fill_1 PHY_632 (  );
sky130_fd_sc_hd__fill_1 PHY_633 (  );
sky130_fd_sc_hd__fill_1 PHY_634 (  );
sky130_fd_sc_hd__fill_1 PHY_635 (  );
sky130_fd_sc_hd__fill_1 PHY_636 (  );
sky130_fd_sc_hd__fill_1 PHY_637 (  );
sky130_fd_sc_hd__fill_1 PHY_638 (  );
sky130_fd_sc_hd__fill_1 PHY_639 (  );
sky130_fd_sc_hd__fill_1 PHY_64 (  );
sky130_fd_sc_hd__fill_1 PHY_640 (  );
sky130_fd_sc_hd__fill_1 PHY_641 (  );
sky130_fd_sc_hd__fill_1 PHY_642 (  );
sky130_fd_sc_hd__fill_1 PHY_643 (  );
sky130_fd_sc_hd__fill_1 PHY_644 (  );
sky130_fd_sc_hd__fill_1 PHY_645 (  );
sky130_fd_sc_hd__fill_1 PHY_646 (  );
sky130_fd_sc_hd__fill_1 PHY_647 (  );
sky130_fd_sc_hd__fill_1 PHY_648 (  );
sky130_fd_sc_hd__fill_1 PHY_649 (  );
sky130_fd_sc_hd__fill_1 PHY_65 (  );
sky130_fd_sc_hd__fill_1 PHY_650 (  );
sky130_fd_sc_hd__fill_1 PHY_651 (  );
sky130_fd_sc_hd__fill_1 PHY_652 (  );
sky130_fd_sc_hd__fill_1 PHY_653 (  );
sky130_fd_sc_hd__fill_1 PHY_654 (  );
sky130_fd_sc_hd__fill_1 PHY_655 (  );
sky130_fd_sc_hd__fill_1 PHY_656 (  );
sky130_fd_sc_hd__fill_1 PHY_657 (  );
sky130_fd_sc_hd__fill_1 PHY_658 (  );
sky130_fd_sc_hd__fill_1 PHY_659 (  );
sky130_fd_sc_hd__fill_1 PHY_66 (  );
sky130_fd_sc_hd__fill_1 PHY_660 (  );
sky130_fd_sc_hd__fill_1 PHY_661 (  );
sky130_fd_sc_hd__fill_1 PHY_662 (  );
sky130_fd_sc_hd__fill_1 PHY_663 (  );
sky130_fd_sc_hd__fill_1 PHY_664 (  );
sky130_fd_sc_hd__fill_1 PHY_665 (  );
sky130_fd_sc_hd__fill_1 PHY_666 (  );
sky130_fd_sc_hd__fill_1 PHY_667 (  );
sky130_fd_sc_hd__fill_1 PHY_668 (  );
sky130_fd_sc_hd__fill_1 PHY_669 (  );
sky130_fd_sc_hd__fill_1 PHY_67 (  );
sky130_fd_sc_hd__fill_1 PHY_670 (  );
sky130_fd_sc_hd__fill_1 PHY_671 (  );
sky130_fd_sc_hd__fill_1 PHY_672 (  );
sky130_fd_sc_hd__fill_1 PHY_673 (  );
sky130_fd_sc_hd__fill_1 PHY_674 (  );
sky130_fd_sc_hd__fill_1 PHY_675 (  );
sky130_fd_sc_hd__fill_1 PHY_676 (  );
sky130_fd_sc_hd__fill_1 PHY_677 (  );
sky130_fd_sc_hd__fill_1 PHY_678 (  );
sky130_fd_sc_hd__fill_1 PHY_679 (  );
sky130_fd_sc_hd__fill_1 PHY_68 (  );
sky130_fd_sc_hd__fill_1 PHY_680 (  );
sky130_fd_sc_hd__fill_1 PHY_681 (  );
sky130_fd_sc_hd__fill_1 PHY_682 (  );
sky130_fd_sc_hd__fill_1 PHY_683 (  );
sky130_fd_sc_hd__fill_1 PHY_684 (  );
sky130_fd_sc_hd__fill_1 PHY_685 (  );
sky130_fd_sc_hd__fill_1 PHY_686 (  );
sky130_fd_sc_hd__fill_1 PHY_687 (  );
sky130_fd_sc_hd__fill_1 PHY_688 (  );
sky130_fd_sc_hd__fill_1 PHY_689 (  );
sky130_fd_sc_hd__fill_1 PHY_69 (  );
sky130_fd_sc_hd__fill_1 PHY_690 (  );
sky130_fd_sc_hd__fill_1 PHY_691 (  );
sky130_fd_sc_hd__fill_1 PHY_692 (  );
sky130_fd_sc_hd__fill_1 PHY_693 (  );
sky130_fd_sc_hd__fill_1 PHY_694 (  );
sky130_fd_sc_hd__fill_1 PHY_695 (  );
sky130_fd_sc_hd__fill_1 PHY_696 (  );
sky130_fd_sc_hd__fill_1 PHY_697 (  );
sky130_fd_sc_hd__fill_1 PHY_698 (  );
sky130_fd_sc_hd__fill_1 PHY_699 (  );
sky130_fd_sc_hd__fill_1 PHY_7 (  );
sky130_fd_sc_hd__fill_1 PHY_70 (  );
sky130_fd_sc_hd__fill_1 PHY_700 (  );
sky130_fd_sc_hd__fill_1 PHY_701 (  );
sky130_fd_sc_hd__fill_1 PHY_702 (  );
sky130_fd_sc_hd__fill_1 PHY_703 (  );
sky130_fd_sc_hd__fill_1 PHY_704 (  );
sky130_fd_sc_hd__fill_1 PHY_705 (  );
sky130_fd_sc_hd__fill_1 PHY_706 (  );
sky130_fd_sc_hd__fill_1 PHY_707 (  );
sky130_fd_sc_hd__fill_1 PHY_708 (  );
sky130_fd_sc_hd__fill_1 PHY_709 (  );
sky130_fd_sc_hd__fill_1 PHY_71 (  );
sky130_fd_sc_hd__fill_1 PHY_710 (  );
sky130_fd_sc_hd__fill_1 PHY_711 (  );
sky130_fd_sc_hd__fill_1 PHY_712 (  );
sky130_fd_sc_hd__fill_1 PHY_713 (  );
sky130_fd_sc_hd__fill_1 PHY_714 (  );
sky130_fd_sc_hd__fill_1 PHY_715 (  );
sky130_fd_sc_hd__fill_1 PHY_716 (  );
sky130_fd_sc_hd__fill_1 PHY_717 (  );
sky130_fd_sc_hd__fill_1 PHY_718 (  );
sky130_fd_sc_hd__fill_1 PHY_719 (  );
sky130_fd_sc_hd__fill_1 PHY_72 (  );
sky130_fd_sc_hd__fill_1 PHY_720 (  );
sky130_fd_sc_hd__fill_1 PHY_721 (  );
sky130_fd_sc_hd__fill_1 PHY_722 (  );
sky130_fd_sc_hd__fill_1 PHY_723 (  );
sky130_fd_sc_hd__fill_1 PHY_724 (  );
sky130_fd_sc_hd__fill_1 PHY_725 (  );
sky130_fd_sc_hd__fill_1 PHY_726 (  );
sky130_fd_sc_hd__fill_1 PHY_727 (  );
sky130_fd_sc_hd__fill_1 PHY_728 (  );
sky130_fd_sc_hd__fill_1 PHY_729 (  );
sky130_fd_sc_hd__fill_1 PHY_73 (  );
sky130_fd_sc_hd__fill_1 PHY_730 (  );
sky130_fd_sc_hd__fill_1 PHY_731 (  );
sky130_fd_sc_hd__fill_1 PHY_732 (  );
sky130_fd_sc_hd__fill_1 PHY_733 (  );
sky130_fd_sc_hd__fill_1 PHY_74 (  );
sky130_fd_sc_hd__fill_1 PHY_75 (  );
sky130_fd_sc_hd__fill_1 PHY_76 (  );
sky130_fd_sc_hd__fill_1 PHY_77 (  );
sky130_fd_sc_hd__fill_1 PHY_78 (  );
sky130_fd_sc_hd__fill_1 PHY_79 (  );
sky130_fd_sc_hd__fill_1 PHY_8 (  );
sky130_fd_sc_hd__fill_1 PHY_80 (  );
sky130_fd_sc_hd__fill_1 PHY_81 (  );
sky130_fd_sc_hd__fill_1 PHY_82 (  );
sky130_fd_sc_hd__fill_1 PHY_83 (  );
sky130_fd_sc_hd__fill_1 PHY_84 (  );
sky130_fd_sc_hd__fill_1 PHY_85 (  );
sky130_fd_sc_hd__fill_1 PHY_86 (  );
sky130_fd_sc_hd__fill_1 PHY_87 (  );
sky130_fd_sc_hd__fill_1 PHY_88 (  );
sky130_fd_sc_hd__fill_1 PHY_89 (  );
sky130_fd_sc_hd__fill_1 PHY_9 (  );
sky130_fd_sc_hd__fill_1 PHY_90 (  );
sky130_fd_sc_hd__fill_1 PHY_91 (  );
sky130_fd_sc_hd__fill_1 PHY_92 (  );
sky130_fd_sc_hd__fill_1 PHY_93 (  );
sky130_fd_sc_hd__fill_1 PHY_94 (  );
sky130_fd_sc_hd__fill_1 PHY_95 (  );
sky130_fd_sc_hd__fill_1 PHY_96 (  );
sky130_fd_sc_hd__fill_1 PHY_97 (  );
sky130_fd_sc_hd__fill_1 PHY_98 (  );
sky130_fd_sc_hd__fill_1 PHY_99 (  );
sky130_fd_sc_hd__tap_1 TAP_1000 (  );
sky130_fd_sc_hd__tap_1 TAP_10000 (  );
sky130_fd_sc_hd__tap_1 TAP_10001 (  );
sky130_fd_sc_hd__tap_1 TAP_10002 (  );
sky130_fd_sc_hd__tap_1 TAP_10003 (  );
sky130_fd_sc_hd__tap_1 TAP_10004 (  );
sky130_fd_sc_hd__tap_1 TAP_10005 (  );
sky130_fd_sc_hd__tap_1 TAP_10006 (  );
sky130_fd_sc_hd__tap_1 TAP_10007 (  );
sky130_fd_sc_hd__tap_1 TAP_10008 (  );
sky130_fd_sc_hd__tap_1 TAP_10009 (  );
sky130_fd_sc_hd__tap_1 TAP_1001 (  );
sky130_fd_sc_hd__tap_1 TAP_10010 (  );
sky130_fd_sc_hd__tap_1 TAP_10011 (  );
sky130_fd_sc_hd__tap_1 TAP_10012 (  );
sky130_fd_sc_hd__tap_1 TAP_10013 (  );
sky130_fd_sc_hd__tap_1 TAP_10014 (  );
sky130_fd_sc_hd__tap_1 TAP_10015 (  );
sky130_fd_sc_hd__tap_1 TAP_10016 (  );
sky130_fd_sc_hd__tap_1 TAP_10017 (  );
sky130_fd_sc_hd__tap_1 TAP_10018 (  );
sky130_fd_sc_hd__tap_1 TAP_10019 (  );
sky130_fd_sc_hd__tap_1 TAP_1002 (  );
sky130_fd_sc_hd__tap_1 TAP_10020 (  );
sky130_fd_sc_hd__tap_1 TAP_10021 (  );
sky130_fd_sc_hd__tap_1 TAP_10022 (  );
sky130_fd_sc_hd__tap_1 TAP_10023 (  );
sky130_fd_sc_hd__tap_1 TAP_10024 (  );
sky130_fd_sc_hd__tap_1 TAP_10025 (  );
sky130_fd_sc_hd__tap_1 TAP_10026 (  );
sky130_fd_sc_hd__tap_1 TAP_10027 (  );
sky130_fd_sc_hd__tap_1 TAP_10028 (  );
sky130_fd_sc_hd__tap_1 TAP_10029 (  );
sky130_fd_sc_hd__tap_1 TAP_1003 (  );
sky130_fd_sc_hd__tap_1 TAP_10030 (  );
sky130_fd_sc_hd__tap_1 TAP_10031 (  );
sky130_fd_sc_hd__tap_1 TAP_10032 (  );
sky130_fd_sc_hd__tap_1 TAP_10033 (  );
sky130_fd_sc_hd__tap_1 TAP_10034 (  );
sky130_fd_sc_hd__tap_1 TAP_10035 (  );
sky130_fd_sc_hd__tap_1 TAP_10036 (  );
sky130_fd_sc_hd__tap_1 TAP_10037 (  );
sky130_fd_sc_hd__tap_1 TAP_10038 (  );
sky130_fd_sc_hd__tap_1 TAP_10039 (  );
sky130_fd_sc_hd__tap_1 TAP_1004 (  );
sky130_fd_sc_hd__tap_1 TAP_10040 (  );
sky130_fd_sc_hd__tap_1 TAP_10041 (  );
sky130_fd_sc_hd__tap_1 TAP_10042 (  );
sky130_fd_sc_hd__tap_1 TAP_10043 (  );
sky130_fd_sc_hd__tap_1 TAP_10044 (  );
sky130_fd_sc_hd__tap_1 TAP_10045 (  );
sky130_fd_sc_hd__tap_1 TAP_10046 (  );
sky130_fd_sc_hd__tap_1 TAP_10047 (  );
sky130_fd_sc_hd__tap_1 TAP_10048 (  );
sky130_fd_sc_hd__tap_1 TAP_10049 (  );
sky130_fd_sc_hd__tap_1 TAP_1005 (  );
sky130_fd_sc_hd__tap_1 TAP_10050 (  );
sky130_fd_sc_hd__tap_1 TAP_10051 (  );
sky130_fd_sc_hd__tap_1 TAP_10052 (  );
sky130_fd_sc_hd__tap_1 TAP_10053 (  );
sky130_fd_sc_hd__tap_1 TAP_10054 (  );
sky130_fd_sc_hd__tap_1 TAP_10055 (  );
sky130_fd_sc_hd__tap_1 TAP_10056 (  );
sky130_fd_sc_hd__tap_1 TAP_10057 (  );
sky130_fd_sc_hd__tap_1 TAP_10058 (  );
sky130_fd_sc_hd__tap_1 TAP_10059 (  );
sky130_fd_sc_hd__tap_1 TAP_1006 (  );
sky130_fd_sc_hd__tap_1 TAP_10060 (  );
sky130_fd_sc_hd__tap_1 TAP_10061 (  );
sky130_fd_sc_hd__tap_1 TAP_10062 (  );
sky130_fd_sc_hd__tap_1 TAP_10063 (  );
sky130_fd_sc_hd__tap_1 TAP_10064 (  );
sky130_fd_sc_hd__tap_1 TAP_10065 (  );
sky130_fd_sc_hd__tap_1 TAP_10066 (  );
sky130_fd_sc_hd__tap_1 TAP_10067 (  );
sky130_fd_sc_hd__tap_1 TAP_10068 (  );
sky130_fd_sc_hd__tap_1 TAP_10069 (  );
sky130_fd_sc_hd__tap_1 TAP_1007 (  );
sky130_fd_sc_hd__tap_1 TAP_10070 (  );
sky130_fd_sc_hd__tap_1 TAP_10071 (  );
sky130_fd_sc_hd__tap_1 TAP_10072 (  );
sky130_fd_sc_hd__tap_1 TAP_10073 (  );
sky130_fd_sc_hd__tap_1 TAP_10074 (  );
sky130_fd_sc_hd__tap_1 TAP_10075 (  );
sky130_fd_sc_hd__tap_1 TAP_10076 (  );
sky130_fd_sc_hd__tap_1 TAP_10077 (  );
sky130_fd_sc_hd__tap_1 TAP_10078 (  );
sky130_fd_sc_hd__tap_1 TAP_10079 (  );
sky130_fd_sc_hd__tap_1 TAP_1008 (  );
sky130_fd_sc_hd__tap_1 TAP_10080 (  );
sky130_fd_sc_hd__tap_1 TAP_10081 (  );
sky130_fd_sc_hd__tap_1 TAP_10082 (  );
sky130_fd_sc_hd__tap_1 TAP_10083 (  );
sky130_fd_sc_hd__tap_1 TAP_10084 (  );
sky130_fd_sc_hd__tap_1 TAP_10085 (  );
sky130_fd_sc_hd__tap_1 TAP_10086 (  );
sky130_fd_sc_hd__tap_1 TAP_10087 (  );
sky130_fd_sc_hd__tap_1 TAP_10088 (  );
sky130_fd_sc_hd__tap_1 TAP_10089 (  );
sky130_fd_sc_hd__tap_1 TAP_1009 (  );
sky130_fd_sc_hd__tap_1 TAP_10090 (  );
sky130_fd_sc_hd__tap_1 TAP_10091 (  );
sky130_fd_sc_hd__tap_1 TAP_10092 (  );
sky130_fd_sc_hd__tap_1 TAP_10093 (  );
sky130_fd_sc_hd__tap_1 TAP_10094 (  );
sky130_fd_sc_hd__tap_1 TAP_10095 (  );
sky130_fd_sc_hd__tap_1 TAP_10096 (  );
sky130_fd_sc_hd__tap_1 TAP_10097 (  );
sky130_fd_sc_hd__tap_1 TAP_10098 (  );
sky130_fd_sc_hd__tap_1 TAP_10099 (  );
sky130_fd_sc_hd__tap_1 TAP_1010 (  );
sky130_fd_sc_hd__tap_1 TAP_10100 (  );
sky130_fd_sc_hd__tap_1 TAP_10101 (  );
sky130_fd_sc_hd__tap_1 TAP_10102 (  );
sky130_fd_sc_hd__tap_1 TAP_10103 (  );
sky130_fd_sc_hd__tap_1 TAP_10104 (  );
sky130_fd_sc_hd__tap_1 TAP_10105 (  );
sky130_fd_sc_hd__tap_1 TAP_10106 (  );
sky130_fd_sc_hd__tap_1 TAP_10107 (  );
sky130_fd_sc_hd__tap_1 TAP_10108 (  );
sky130_fd_sc_hd__tap_1 TAP_10109 (  );
sky130_fd_sc_hd__tap_1 TAP_1011 (  );
sky130_fd_sc_hd__tap_1 TAP_10110 (  );
sky130_fd_sc_hd__tap_1 TAP_10111 (  );
sky130_fd_sc_hd__tap_1 TAP_10112 (  );
sky130_fd_sc_hd__tap_1 TAP_10113 (  );
sky130_fd_sc_hd__tap_1 TAP_10114 (  );
sky130_fd_sc_hd__tap_1 TAP_10115 (  );
sky130_fd_sc_hd__tap_1 TAP_10116 (  );
sky130_fd_sc_hd__tap_1 TAP_10117 (  );
sky130_fd_sc_hd__tap_1 TAP_10118 (  );
sky130_fd_sc_hd__tap_1 TAP_10119 (  );
sky130_fd_sc_hd__tap_1 TAP_1012 (  );
sky130_fd_sc_hd__tap_1 TAP_10120 (  );
sky130_fd_sc_hd__tap_1 TAP_10121 (  );
sky130_fd_sc_hd__tap_1 TAP_10122 (  );
sky130_fd_sc_hd__tap_1 TAP_10123 (  );
sky130_fd_sc_hd__tap_1 TAP_10124 (  );
sky130_fd_sc_hd__tap_1 TAP_10125 (  );
sky130_fd_sc_hd__tap_1 TAP_10126 (  );
sky130_fd_sc_hd__tap_1 TAP_10127 (  );
sky130_fd_sc_hd__tap_1 TAP_10128 (  );
sky130_fd_sc_hd__tap_1 TAP_10129 (  );
sky130_fd_sc_hd__tap_1 TAP_1013 (  );
sky130_fd_sc_hd__tap_1 TAP_10130 (  );
sky130_fd_sc_hd__tap_1 TAP_10131 (  );
sky130_fd_sc_hd__tap_1 TAP_10132 (  );
sky130_fd_sc_hd__tap_1 TAP_10133 (  );
sky130_fd_sc_hd__tap_1 TAP_10134 (  );
sky130_fd_sc_hd__tap_1 TAP_10135 (  );
sky130_fd_sc_hd__tap_1 TAP_10136 (  );
sky130_fd_sc_hd__tap_1 TAP_10137 (  );
sky130_fd_sc_hd__tap_1 TAP_10138 (  );
sky130_fd_sc_hd__tap_1 TAP_10139 (  );
sky130_fd_sc_hd__tap_1 TAP_1014 (  );
sky130_fd_sc_hd__tap_1 TAP_10140 (  );
sky130_fd_sc_hd__tap_1 TAP_10141 (  );
sky130_fd_sc_hd__tap_1 TAP_10142 (  );
sky130_fd_sc_hd__tap_1 TAP_10143 (  );
sky130_fd_sc_hd__tap_1 TAP_10144 (  );
sky130_fd_sc_hd__tap_1 TAP_10145 (  );
sky130_fd_sc_hd__tap_1 TAP_10146 (  );
sky130_fd_sc_hd__tap_1 TAP_10147 (  );
sky130_fd_sc_hd__tap_1 TAP_10148 (  );
sky130_fd_sc_hd__tap_1 TAP_10149 (  );
sky130_fd_sc_hd__tap_1 TAP_1015 (  );
sky130_fd_sc_hd__tap_1 TAP_10150 (  );
sky130_fd_sc_hd__tap_1 TAP_10151 (  );
sky130_fd_sc_hd__tap_1 TAP_10152 (  );
sky130_fd_sc_hd__tap_1 TAP_10153 (  );
sky130_fd_sc_hd__tap_1 TAP_10154 (  );
sky130_fd_sc_hd__tap_1 TAP_10155 (  );
sky130_fd_sc_hd__tap_1 TAP_10156 (  );
sky130_fd_sc_hd__tap_1 TAP_10157 (  );
sky130_fd_sc_hd__tap_1 TAP_10158 (  );
sky130_fd_sc_hd__tap_1 TAP_10159 (  );
sky130_fd_sc_hd__tap_1 TAP_1016 (  );
sky130_fd_sc_hd__tap_1 TAP_10160 (  );
sky130_fd_sc_hd__tap_1 TAP_10161 (  );
sky130_fd_sc_hd__tap_1 TAP_10162 (  );
sky130_fd_sc_hd__tap_1 TAP_10163 (  );
sky130_fd_sc_hd__tap_1 TAP_10164 (  );
sky130_fd_sc_hd__tap_1 TAP_10165 (  );
sky130_fd_sc_hd__tap_1 TAP_10166 (  );
sky130_fd_sc_hd__tap_1 TAP_10167 (  );
sky130_fd_sc_hd__tap_1 TAP_10168 (  );
sky130_fd_sc_hd__tap_1 TAP_10169 (  );
sky130_fd_sc_hd__tap_1 TAP_1017 (  );
sky130_fd_sc_hd__tap_1 TAP_10170 (  );
sky130_fd_sc_hd__tap_1 TAP_10171 (  );
sky130_fd_sc_hd__tap_1 TAP_10172 (  );
sky130_fd_sc_hd__tap_1 TAP_10173 (  );
sky130_fd_sc_hd__tap_1 TAP_10174 (  );
sky130_fd_sc_hd__tap_1 TAP_10175 (  );
sky130_fd_sc_hd__tap_1 TAP_10176 (  );
sky130_fd_sc_hd__tap_1 TAP_10177 (  );
sky130_fd_sc_hd__tap_1 TAP_10178 (  );
sky130_fd_sc_hd__tap_1 TAP_10179 (  );
sky130_fd_sc_hd__tap_1 TAP_1018 (  );
sky130_fd_sc_hd__tap_1 TAP_10180 (  );
sky130_fd_sc_hd__tap_1 TAP_10181 (  );
sky130_fd_sc_hd__tap_1 TAP_10182 (  );
sky130_fd_sc_hd__tap_1 TAP_10183 (  );
sky130_fd_sc_hd__tap_1 TAP_10184 (  );
sky130_fd_sc_hd__tap_1 TAP_10185 (  );
sky130_fd_sc_hd__tap_1 TAP_10186 (  );
sky130_fd_sc_hd__tap_1 TAP_10187 (  );
sky130_fd_sc_hd__tap_1 TAP_10188 (  );
sky130_fd_sc_hd__tap_1 TAP_10189 (  );
sky130_fd_sc_hd__tap_1 TAP_1019 (  );
sky130_fd_sc_hd__tap_1 TAP_10190 (  );
sky130_fd_sc_hd__tap_1 TAP_10191 (  );
sky130_fd_sc_hd__tap_1 TAP_10192 (  );
sky130_fd_sc_hd__tap_1 TAP_10193 (  );
sky130_fd_sc_hd__tap_1 TAP_10194 (  );
sky130_fd_sc_hd__tap_1 TAP_10195 (  );
sky130_fd_sc_hd__tap_1 TAP_10196 (  );
sky130_fd_sc_hd__tap_1 TAP_10197 (  );
sky130_fd_sc_hd__tap_1 TAP_10198 (  );
sky130_fd_sc_hd__tap_1 TAP_10199 (  );
sky130_fd_sc_hd__tap_1 TAP_1020 (  );
sky130_fd_sc_hd__tap_1 TAP_10200 (  );
sky130_fd_sc_hd__tap_1 TAP_10201 (  );
sky130_fd_sc_hd__tap_1 TAP_10202 (  );
sky130_fd_sc_hd__tap_1 TAP_10203 (  );
sky130_fd_sc_hd__tap_1 TAP_10204 (  );
sky130_fd_sc_hd__tap_1 TAP_10205 (  );
sky130_fd_sc_hd__tap_1 TAP_10206 (  );
sky130_fd_sc_hd__tap_1 TAP_10207 (  );
sky130_fd_sc_hd__tap_1 TAP_10208 (  );
sky130_fd_sc_hd__tap_1 TAP_10209 (  );
sky130_fd_sc_hd__tap_1 TAP_1021 (  );
sky130_fd_sc_hd__tap_1 TAP_10210 (  );
sky130_fd_sc_hd__tap_1 TAP_10211 (  );
sky130_fd_sc_hd__tap_1 TAP_10212 (  );
sky130_fd_sc_hd__tap_1 TAP_10213 (  );
sky130_fd_sc_hd__tap_1 TAP_10214 (  );
sky130_fd_sc_hd__tap_1 TAP_10215 (  );
sky130_fd_sc_hd__tap_1 TAP_10216 (  );
sky130_fd_sc_hd__tap_1 TAP_10217 (  );
sky130_fd_sc_hd__tap_1 TAP_10218 (  );
sky130_fd_sc_hd__tap_1 TAP_10219 (  );
sky130_fd_sc_hd__tap_1 TAP_1022 (  );
sky130_fd_sc_hd__tap_1 TAP_10220 (  );
sky130_fd_sc_hd__tap_1 TAP_10221 (  );
sky130_fd_sc_hd__tap_1 TAP_10222 (  );
sky130_fd_sc_hd__tap_1 TAP_10223 (  );
sky130_fd_sc_hd__tap_1 TAP_10224 (  );
sky130_fd_sc_hd__tap_1 TAP_10225 (  );
sky130_fd_sc_hd__tap_1 TAP_10226 (  );
sky130_fd_sc_hd__tap_1 TAP_10227 (  );
sky130_fd_sc_hd__tap_1 TAP_10228 (  );
sky130_fd_sc_hd__tap_1 TAP_10229 (  );
sky130_fd_sc_hd__tap_1 TAP_1023 (  );
sky130_fd_sc_hd__tap_1 TAP_10230 (  );
sky130_fd_sc_hd__tap_1 TAP_10231 (  );
sky130_fd_sc_hd__tap_1 TAP_10232 (  );
sky130_fd_sc_hd__tap_1 TAP_10233 (  );
sky130_fd_sc_hd__tap_1 TAP_10234 (  );
sky130_fd_sc_hd__tap_1 TAP_10235 (  );
sky130_fd_sc_hd__tap_1 TAP_10236 (  );
sky130_fd_sc_hd__tap_1 TAP_10237 (  );
sky130_fd_sc_hd__tap_1 TAP_10238 (  );
sky130_fd_sc_hd__tap_1 TAP_10239 (  );
sky130_fd_sc_hd__tap_1 TAP_1024 (  );
sky130_fd_sc_hd__tap_1 TAP_10240 (  );
sky130_fd_sc_hd__tap_1 TAP_10241 (  );
sky130_fd_sc_hd__tap_1 TAP_10242 (  );
sky130_fd_sc_hd__tap_1 TAP_10243 (  );
sky130_fd_sc_hd__tap_1 TAP_10244 (  );
sky130_fd_sc_hd__tap_1 TAP_10245 (  );
sky130_fd_sc_hd__tap_1 TAP_10246 (  );
sky130_fd_sc_hd__tap_1 TAP_10247 (  );
sky130_fd_sc_hd__tap_1 TAP_10248 (  );
sky130_fd_sc_hd__tap_1 TAP_10249 (  );
sky130_fd_sc_hd__tap_1 TAP_1025 (  );
sky130_fd_sc_hd__tap_1 TAP_10250 (  );
sky130_fd_sc_hd__tap_1 TAP_10251 (  );
sky130_fd_sc_hd__tap_1 TAP_10252 (  );
sky130_fd_sc_hd__tap_1 TAP_10253 (  );
sky130_fd_sc_hd__tap_1 TAP_10254 (  );
sky130_fd_sc_hd__tap_1 TAP_10255 (  );
sky130_fd_sc_hd__tap_1 TAP_10256 (  );
sky130_fd_sc_hd__tap_1 TAP_10257 (  );
sky130_fd_sc_hd__tap_1 TAP_10258 (  );
sky130_fd_sc_hd__tap_1 TAP_10259 (  );
sky130_fd_sc_hd__tap_1 TAP_1026 (  );
sky130_fd_sc_hd__tap_1 TAP_10260 (  );
sky130_fd_sc_hd__tap_1 TAP_10261 (  );
sky130_fd_sc_hd__tap_1 TAP_10262 (  );
sky130_fd_sc_hd__tap_1 TAP_10263 (  );
sky130_fd_sc_hd__tap_1 TAP_10264 (  );
sky130_fd_sc_hd__tap_1 TAP_10265 (  );
sky130_fd_sc_hd__tap_1 TAP_10266 (  );
sky130_fd_sc_hd__tap_1 TAP_10267 (  );
sky130_fd_sc_hd__tap_1 TAP_10268 (  );
sky130_fd_sc_hd__tap_1 TAP_10269 (  );
sky130_fd_sc_hd__tap_1 TAP_1027 (  );
sky130_fd_sc_hd__tap_1 TAP_10270 (  );
sky130_fd_sc_hd__tap_1 TAP_10271 (  );
sky130_fd_sc_hd__tap_1 TAP_10272 (  );
sky130_fd_sc_hd__tap_1 TAP_10273 (  );
sky130_fd_sc_hd__tap_1 TAP_10274 (  );
sky130_fd_sc_hd__tap_1 TAP_10275 (  );
sky130_fd_sc_hd__tap_1 TAP_10276 (  );
sky130_fd_sc_hd__tap_1 TAP_10277 (  );
sky130_fd_sc_hd__tap_1 TAP_10278 (  );
sky130_fd_sc_hd__tap_1 TAP_10279 (  );
sky130_fd_sc_hd__tap_1 TAP_1028 (  );
sky130_fd_sc_hd__tap_1 TAP_10280 (  );
sky130_fd_sc_hd__tap_1 TAP_10281 (  );
sky130_fd_sc_hd__tap_1 TAP_10282 (  );
sky130_fd_sc_hd__tap_1 TAP_10283 (  );
sky130_fd_sc_hd__tap_1 TAP_10284 (  );
sky130_fd_sc_hd__tap_1 TAP_10285 (  );
sky130_fd_sc_hd__tap_1 TAP_10286 (  );
sky130_fd_sc_hd__tap_1 TAP_10287 (  );
sky130_fd_sc_hd__tap_1 TAP_10288 (  );
sky130_fd_sc_hd__tap_1 TAP_10289 (  );
sky130_fd_sc_hd__tap_1 TAP_1029 (  );
sky130_fd_sc_hd__tap_1 TAP_10290 (  );
sky130_fd_sc_hd__tap_1 TAP_10291 (  );
sky130_fd_sc_hd__tap_1 TAP_10292 (  );
sky130_fd_sc_hd__tap_1 TAP_10293 (  );
sky130_fd_sc_hd__tap_1 TAP_10294 (  );
sky130_fd_sc_hd__tap_1 TAP_10295 (  );
sky130_fd_sc_hd__tap_1 TAP_10296 (  );
sky130_fd_sc_hd__tap_1 TAP_10297 (  );
sky130_fd_sc_hd__tap_1 TAP_10298 (  );
sky130_fd_sc_hd__tap_1 TAP_10299 (  );
sky130_fd_sc_hd__tap_1 TAP_1030 (  );
sky130_fd_sc_hd__tap_1 TAP_10300 (  );
sky130_fd_sc_hd__tap_1 TAP_10301 (  );
sky130_fd_sc_hd__tap_1 TAP_10302 (  );
sky130_fd_sc_hd__tap_1 TAP_10303 (  );
sky130_fd_sc_hd__tap_1 TAP_10304 (  );
sky130_fd_sc_hd__tap_1 TAP_10305 (  );
sky130_fd_sc_hd__tap_1 TAP_10306 (  );
sky130_fd_sc_hd__tap_1 TAP_10307 (  );
sky130_fd_sc_hd__tap_1 TAP_10308 (  );
sky130_fd_sc_hd__tap_1 TAP_10309 (  );
sky130_fd_sc_hd__tap_1 TAP_1031 (  );
sky130_fd_sc_hd__tap_1 TAP_10310 (  );
sky130_fd_sc_hd__tap_1 TAP_10311 (  );
sky130_fd_sc_hd__tap_1 TAP_10312 (  );
sky130_fd_sc_hd__tap_1 TAP_10313 (  );
sky130_fd_sc_hd__tap_1 TAP_10314 (  );
sky130_fd_sc_hd__tap_1 TAP_10315 (  );
sky130_fd_sc_hd__tap_1 TAP_10316 (  );
sky130_fd_sc_hd__tap_1 TAP_10317 (  );
sky130_fd_sc_hd__tap_1 TAP_10318 (  );
sky130_fd_sc_hd__tap_1 TAP_10319 (  );
sky130_fd_sc_hd__tap_1 TAP_1032 (  );
sky130_fd_sc_hd__tap_1 TAP_10320 (  );
sky130_fd_sc_hd__tap_1 TAP_10321 (  );
sky130_fd_sc_hd__tap_1 TAP_10322 (  );
sky130_fd_sc_hd__tap_1 TAP_10323 (  );
sky130_fd_sc_hd__tap_1 TAP_10324 (  );
sky130_fd_sc_hd__tap_1 TAP_10325 (  );
sky130_fd_sc_hd__tap_1 TAP_10326 (  );
sky130_fd_sc_hd__tap_1 TAP_10327 (  );
sky130_fd_sc_hd__tap_1 TAP_10328 (  );
sky130_fd_sc_hd__tap_1 TAP_10329 (  );
sky130_fd_sc_hd__tap_1 TAP_1033 (  );
sky130_fd_sc_hd__tap_1 TAP_10330 (  );
sky130_fd_sc_hd__tap_1 TAP_10331 (  );
sky130_fd_sc_hd__tap_1 TAP_10332 (  );
sky130_fd_sc_hd__tap_1 TAP_10333 (  );
sky130_fd_sc_hd__tap_1 TAP_10334 (  );
sky130_fd_sc_hd__tap_1 TAP_10335 (  );
sky130_fd_sc_hd__tap_1 TAP_10336 (  );
sky130_fd_sc_hd__tap_1 TAP_10337 (  );
sky130_fd_sc_hd__tap_1 TAP_10338 (  );
sky130_fd_sc_hd__tap_1 TAP_10339 (  );
sky130_fd_sc_hd__tap_1 TAP_1034 (  );
sky130_fd_sc_hd__tap_1 TAP_10340 (  );
sky130_fd_sc_hd__tap_1 TAP_10341 (  );
sky130_fd_sc_hd__tap_1 TAP_10342 (  );
sky130_fd_sc_hd__tap_1 TAP_10343 (  );
sky130_fd_sc_hd__tap_1 TAP_10344 (  );
sky130_fd_sc_hd__tap_1 TAP_10345 (  );
sky130_fd_sc_hd__tap_1 TAP_10346 (  );
sky130_fd_sc_hd__tap_1 TAP_10347 (  );
sky130_fd_sc_hd__tap_1 TAP_10348 (  );
sky130_fd_sc_hd__tap_1 TAP_10349 (  );
sky130_fd_sc_hd__tap_1 TAP_1035 (  );
sky130_fd_sc_hd__tap_1 TAP_10350 (  );
sky130_fd_sc_hd__tap_1 TAP_10351 (  );
sky130_fd_sc_hd__tap_1 TAP_10352 (  );
sky130_fd_sc_hd__tap_1 TAP_10353 (  );
sky130_fd_sc_hd__tap_1 TAP_10354 (  );
sky130_fd_sc_hd__tap_1 TAP_10355 (  );
sky130_fd_sc_hd__tap_1 TAP_10356 (  );
sky130_fd_sc_hd__tap_1 TAP_10357 (  );
sky130_fd_sc_hd__tap_1 TAP_10358 (  );
sky130_fd_sc_hd__tap_1 TAP_10359 (  );
sky130_fd_sc_hd__tap_1 TAP_1036 (  );
sky130_fd_sc_hd__tap_1 TAP_10360 (  );
sky130_fd_sc_hd__tap_1 TAP_10361 (  );
sky130_fd_sc_hd__tap_1 TAP_10362 (  );
sky130_fd_sc_hd__tap_1 TAP_10363 (  );
sky130_fd_sc_hd__tap_1 TAP_10364 (  );
sky130_fd_sc_hd__tap_1 TAP_10365 (  );
sky130_fd_sc_hd__tap_1 TAP_10366 (  );
sky130_fd_sc_hd__tap_1 TAP_10367 (  );
sky130_fd_sc_hd__tap_1 TAP_10368 (  );
sky130_fd_sc_hd__tap_1 TAP_10369 (  );
sky130_fd_sc_hd__tap_1 TAP_1037 (  );
sky130_fd_sc_hd__tap_1 TAP_10370 (  );
sky130_fd_sc_hd__tap_1 TAP_10371 (  );
sky130_fd_sc_hd__tap_1 TAP_10372 (  );
sky130_fd_sc_hd__tap_1 TAP_10373 (  );
sky130_fd_sc_hd__tap_1 TAP_10374 (  );
sky130_fd_sc_hd__tap_1 TAP_10375 (  );
sky130_fd_sc_hd__tap_1 TAP_10376 (  );
sky130_fd_sc_hd__tap_1 TAP_10377 (  );
sky130_fd_sc_hd__tap_1 TAP_10378 (  );
sky130_fd_sc_hd__tap_1 TAP_10379 (  );
sky130_fd_sc_hd__tap_1 TAP_1038 (  );
sky130_fd_sc_hd__tap_1 TAP_10380 (  );
sky130_fd_sc_hd__tap_1 TAP_10381 (  );
sky130_fd_sc_hd__tap_1 TAP_10382 (  );
sky130_fd_sc_hd__tap_1 TAP_10383 (  );
sky130_fd_sc_hd__tap_1 TAP_10384 (  );
sky130_fd_sc_hd__tap_1 TAP_10385 (  );
sky130_fd_sc_hd__tap_1 TAP_10386 (  );
sky130_fd_sc_hd__tap_1 TAP_10387 (  );
sky130_fd_sc_hd__tap_1 TAP_10388 (  );
sky130_fd_sc_hd__tap_1 TAP_10389 (  );
sky130_fd_sc_hd__tap_1 TAP_1039 (  );
sky130_fd_sc_hd__tap_1 TAP_10390 (  );
sky130_fd_sc_hd__tap_1 TAP_10391 (  );
sky130_fd_sc_hd__tap_1 TAP_10392 (  );
sky130_fd_sc_hd__tap_1 TAP_10393 (  );
sky130_fd_sc_hd__tap_1 TAP_10394 (  );
sky130_fd_sc_hd__tap_1 TAP_10395 (  );
sky130_fd_sc_hd__tap_1 TAP_10396 (  );
sky130_fd_sc_hd__tap_1 TAP_10397 (  );
sky130_fd_sc_hd__tap_1 TAP_10398 (  );
sky130_fd_sc_hd__tap_1 TAP_10399 (  );
sky130_fd_sc_hd__tap_1 TAP_1040 (  );
sky130_fd_sc_hd__tap_1 TAP_10400 (  );
sky130_fd_sc_hd__tap_1 TAP_10401 (  );
sky130_fd_sc_hd__tap_1 TAP_10402 (  );
sky130_fd_sc_hd__tap_1 TAP_10403 (  );
sky130_fd_sc_hd__tap_1 TAP_10404 (  );
sky130_fd_sc_hd__tap_1 TAP_10405 (  );
sky130_fd_sc_hd__tap_1 TAP_10406 (  );
sky130_fd_sc_hd__tap_1 TAP_10407 (  );
sky130_fd_sc_hd__tap_1 TAP_10408 (  );
sky130_fd_sc_hd__tap_1 TAP_10409 (  );
sky130_fd_sc_hd__tap_1 TAP_1041 (  );
sky130_fd_sc_hd__tap_1 TAP_10410 (  );
sky130_fd_sc_hd__tap_1 TAP_10411 (  );
sky130_fd_sc_hd__tap_1 TAP_10412 (  );
sky130_fd_sc_hd__tap_1 TAP_10413 (  );
sky130_fd_sc_hd__tap_1 TAP_10414 (  );
sky130_fd_sc_hd__tap_1 TAP_10415 (  );
sky130_fd_sc_hd__tap_1 TAP_10416 (  );
sky130_fd_sc_hd__tap_1 TAP_10417 (  );
sky130_fd_sc_hd__tap_1 TAP_10418 (  );
sky130_fd_sc_hd__tap_1 TAP_10419 (  );
sky130_fd_sc_hd__tap_1 TAP_1042 (  );
sky130_fd_sc_hd__tap_1 TAP_10420 (  );
sky130_fd_sc_hd__tap_1 TAP_10421 (  );
sky130_fd_sc_hd__tap_1 TAP_10422 (  );
sky130_fd_sc_hd__tap_1 TAP_10423 (  );
sky130_fd_sc_hd__tap_1 TAP_10424 (  );
sky130_fd_sc_hd__tap_1 TAP_10425 (  );
sky130_fd_sc_hd__tap_1 TAP_10426 (  );
sky130_fd_sc_hd__tap_1 TAP_10427 (  );
sky130_fd_sc_hd__tap_1 TAP_10428 (  );
sky130_fd_sc_hd__tap_1 TAP_10429 (  );
sky130_fd_sc_hd__tap_1 TAP_1043 (  );
sky130_fd_sc_hd__tap_1 TAP_10430 (  );
sky130_fd_sc_hd__tap_1 TAP_10431 (  );
sky130_fd_sc_hd__tap_1 TAP_10432 (  );
sky130_fd_sc_hd__tap_1 TAP_10433 (  );
sky130_fd_sc_hd__tap_1 TAP_10434 (  );
sky130_fd_sc_hd__tap_1 TAP_10435 (  );
sky130_fd_sc_hd__tap_1 TAP_10436 (  );
sky130_fd_sc_hd__tap_1 TAP_10437 (  );
sky130_fd_sc_hd__tap_1 TAP_10438 (  );
sky130_fd_sc_hd__tap_1 TAP_10439 (  );
sky130_fd_sc_hd__tap_1 TAP_1044 (  );
sky130_fd_sc_hd__tap_1 TAP_10440 (  );
sky130_fd_sc_hd__tap_1 TAP_10441 (  );
sky130_fd_sc_hd__tap_1 TAP_10442 (  );
sky130_fd_sc_hd__tap_1 TAP_10443 (  );
sky130_fd_sc_hd__tap_1 TAP_10444 (  );
sky130_fd_sc_hd__tap_1 TAP_10445 (  );
sky130_fd_sc_hd__tap_1 TAP_10446 (  );
sky130_fd_sc_hd__tap_1 TAP_10447 (  );
sky130_fd_sc_hd__tap_1 TAP_10448 (  );
sky130_fd_sc_hd__tap_1 TAP_10449 (  );
sky130_fd_sc_hd__tap_1 TAP_1045 (  );
sky130_fd_sc_hd__tap_1 TAP_10450 (  );
sky130_fd_sc_hd__tap_1 TAP_10451 (  );
sky130_fd_sc_hd__tap_1 TAP_10452 (  );
sky130_fd_sc_hd__tap_1 TAP_10453 (  );
sky130_fd_sc_hd__tap_1 TAP_10454 (  );
sky130_fd_sc_hd__tap_1 TAP_10455 (  );
sky130_fd_sc_hd__tap_1 TAP_10456 (  );
sky130_fd_sc_hd__tap_1 TAP_10457 (  );
sky130_fd_sc_hd__tap_1 TAP_10458 (  );
sky130_fd_sc_hd__tap_1 TAP_10459 (  );
sky130_fd_sc_hd__tap_1 TAP_1046 (  );
sky130_fd_sc_hd__tap_1 TAP_10460 (  );
sky130_fd_sc_hd__tap_1 TAP_10461 (  );
sky130_fd_sc_hd__tap_1 TAP_10462 (  );
sky130_fd_sc_hd__tap_1 TAP_10463 (  );
sky130_fd_sc_hd__tap_1 TAP_10464 (  );
sky130_fd_sc_hd__tap_1 TAP_10465 (  );
sky130_fd_sc_hd__tap_1 TAP_10466 (  );
sky130_fd_sc_hd__tap_1 TAP_10467 (  );
sky130_fd_sc_hd__tap_1 TAP_10468 (  );
sky130_fd_sc_hd__tap_1 TAP_10469 (  );
sky130_fd_sc_hd__tap_1 TAP_1047 (  );
sky130_fd_sc_hd__tap_1 TAP_10470 (  );
sky130_fd_sc_hd__tap_1 TAP_10471 (  );
sky130_fd_sc_hd__tap_1 TAP_10472 (  );
sky130_fd_sc_hd__tap_1 TAP_10473 (  );
sky130_fd_sc_hd__tap_1 TAP_10474 (  );
sky130_fd_sc_hd__tap_1 TAP_10475 (  );
sky130_fd_sc_hd__tap_1 TAP_10476 (  );
sky130_fd_sc_hd__tap_1 TAP_10477 (  );
sky130_fd_sc_hd__tap_1 TAP_10478 (  );
sky130_fd_sc_hd__tap_1 TAP_10479 (  );
sky130_fd_sc_hd__tap_1 TAP_1048 (  );
sky130_fd_sc_hd__tap_1 TAP_10480 (  );
sky130_fd_sc_hd__tap_1 TAP_10481 (  );
sky130_fd_sc_hd__tap_1 TAP_10482 (  );
sky130_fd_sc_hd__tap_1 TAP_10483 (  );
sky130_fd_sc_hd__tap_1 TAP_10484 (  );
sky130_fd_sc_hd__tap_1 TAP_10485 (  );
sky130_fd_sc_hd__tap_1 TAP_10486 (  );
sky130_fd_sc_hd__tap_1 TAP_10487 (  );
sky130_fd_sc_hd__tap_1 TAP_10488 (  );
sky130_fd_sc_hd__tap_1 TAP_10489 (  );
sky130_fd_sc_hd__tap_1 TAP_1049 (  );
sky130_fd_sc_hd__tap_1 TAP_10490 (  );
sky130_fd_sc_hd__tap_1 TAP_10491 (  );
sky130_fd_sc_hd__tap_1 TAP_10492 (  );
sky130_fd_sc_hd__tap_1 TAP_10493 (  );
sky130_fd_sc_hd__tap_1 TAP_10494 (  );
sky130_fd_sc_hd__tap_1 TAP_10495 (  );
sky130_fd_sc_hd__tap_1 TAP_10496 (  );
sky130_fd_sc_hd__tap_1 TAP_10497 (  );
sky130_fd_sc_hd__tap_1 TAP_10498 (  );
sky130_fd_sc_hd__tap_1 TAP_10499 (  );
sky130_fd_sc_hd__tap_1 TAP_1050 (  );
sky130_fd_sc_hd__tap_1 TAP_10500 (  );
sky130_fd_sc_hd__tap_1 TAP_10501 (  );
sky130_fd_sc_hd__tap_1 TAP_10502 (  );
sky130_fd_sc_hd__tap_1 TAP_10503 (  );
sky130_fd_sc_hd__tap_1 TAP_10504 (  );
sky130_fd_sc_hd__tap_1 TAP_10505 (  );
sky130_fd_sc_hd__tap_1 TAP_10506 (  );
sky130_fd_sc_hd__tap_1 TAP_10507 (  );
sky130_fd_sc_hd__tap_1 TAP_10508 (  );
sky130_fd_sc_hd__tap_1 TAP_10509 (  );
sky130_fd_sc_hd__tap_1 TAP_1051 (  );
sky130_fd_sc_hd__tap_1 TAP_10510 (  );
sky130_fd_sc_hd__tap_1 TAP_10511 (  );
sky130_fd_sc_hd__tap_1 TAP_10512 (  );
sky130_fd_sc_hd__tap_1 TAP_10513 (  );
sky130_fd_sc_hd__tap_1 TAP_10514 (  );
sky130_fd_sc_hd__tap_1 TAP_10515 (  );
sky130_fd_sc_hd__tap_1 TAP_10516 (  );
sky130_fd_sc_hd__tap_1 TAP_10517 (  );
sky130_fd_sc_hd__tap_1 TAP_10518 (  );
sky130_fd_sc_hd__tap_1 TAP_10519 (  );
sky130_fd_sc_hd__tap_1 TAP_1052 (  );
sky130_fd_sc_hd__tap_1 TAP_10520 (  );
sky130_fd_sc_hd__tap_1 TAP_10521 (  );
sky130_fd_sc_hd__tap_1 TAP_10522 (  );
sky130_fd_sc_hd__tap_1 TAP_10523 (  );
sky130_fd_sc_hd__tap_1 TAP_10524 (  );
sky130_fd_sc_hd__tap_1 TAP_10525 (  );
sky130_fd_sc_hd__tap_1 TAP_10526 (  );
sky130_fd_sc_hd__tap_1 TAP_10527 (  );
sky130_fd_sc_hd__tap_1 TAP_10528 (  );
sky130_fd_sc_hd__tap_1 TAP_10529 (  );
sky130_fd_sc_hd__tap_1 TAP_1053 (  );
sky130_fd_sc_hd__tap_1 TAP_10530 (  );
sky130_fd_sc_hd__tap_1 TAP_10531 (  );
sky130_fd_sc_hd__tap_1 TAP_10532 (  );
sky130_fd_sc_hd__tap_1 TAP_10533 (  );
sky130_fd_sc_hd__tap_1 TAP_10534 (  );
sky130_fd_sc_hd__tap_1 TAP_10535 (  );
sky130_fd_sc_hd__tap_1 TAP_10536 (  );
sky130_fd_sc_hd__tap_1 TAP_10537 (  );
sky130_fd_sc_hd__tap_1 TAP_10538 (  );
sky130_fd_sc_hd__tap_1 TAP_10539 (  );
sky130_fd_sc_hd__tap_1 TAP_1054 (  );
sky130_fd_sc_hd__tap_1 TAP_10540 (  );
sky130_fd_sc_hd__tap_1 TAP_10541 (  );
sky130_fd_sc_hd__tap_1 TAP_10542 (  );
sky130_fd_sc_hd__tap_1 TAP_10543 (  );
sky130_fd_sc_hd__tap_1 TAP_10544 (  );
sky130_fd_sc_hd__tap_1 TAP_10545 (  );
sky130_fd_sc_hd__tap_1 TAP_10546 (  );
sky130_fd_sc_hd__tap_1 TAP_10547 (  );
sky130_fd_sc_hd__tap_1 TAP_10548 (  );
sky130_fd_sc_hd__tap_1 TAP_10549 (  );
sky130_fd_sc_hd__tap_1 TAP_1055 (  );
sky130_fd_sc_hd__tap_1 TAP_10550 (  );
sky130_fd_sc_hd__tap_1 TAP_10551 (  );
sky130_fd_sc_hd__tap_1 TAP_10552 (  );
sky130_fd_sc_hd__tap_1 TAP_10553 (  );
sky130_fd_sc_hd__tap_1 TAP_10554 (  );
sky130_fd_sc_hd__tap_1 TAP_10555 (  );
sky130_fd_sc_hd__tap_1 TAP_10556 (  );
sky130_fd_sc_hd__tap_1 TAP_10557 (  );
sky130_fd_sc_hd__tap_1 TAP_10558 (  );
sky130_fd_sc_hd__tap_1 TAP_10559 (  );
sky130_fd_sc_hd__tap_1 TAP_1056 (  );
sky130_fd_sc_hd__tap_1 TAP_10560 (  );
sky130_fd_sc_hd__tap_1 TAP_10561 (  );
sky130_fd_sc_hd__tap_1 TAP_10562 (  );
sky130_fd_sc_hd__tap_1 TAP_10563 (  );
sky130_fd_sc_hd__tap_1 TAP_10564 (  );
sky130_fd_sc_hd__tap_1 TAP_10565 (  );
sky130_fd_sc_hd__tap_1 TAP_10566 (  );
sky130_fd_sc_hd__tap_1 TAP_10567 (  );
sky130_fd_sc_hd__tap_1 TAP_10568 (  );
sky130_fd_sc_hd__tap_1 TAP_10569 (  );
sky130_fd_sc_hd__tap_1 TAP_1057 (  );
sky130_fd_sc_hd__tap_1 TAP_10570 (  );
sky130_fd_sc_hd__tap_1 TAP_10571 (  );
sky130_fd_sc_hd__tap_1 TAP_10572 (  );
sky130_fd_sc_hd__tap_1 TAP_10573 (  );
sky130_fd_sc_hd__tap_1 TAP_10574 (  );
sky130_fd_sc_hd__tap_1 TAP_10575 (  );
sky130_fd_sc_hd__tap_1 TAP_10576 (  );
sky130_fd_sc_hd__tap_1 TAP_10577 (  );
sky130_fd_sc_hd__tap_1 TAP_10578 (  );
sky130_fd_sc_hd__tap_1 TAP_10579 (  );
sky130_fd_sc_hd__tap_1 TAP_1058 (  );
sky130_fd_sc_hd__tap_1 TAP_10580 (  );
sky130_fd_sc_hd__tap_1 TAP_10581 (  );
sky130_fd_sc_hd__tap_1 TAP_10582 (  );
sky130_fd_sc_hd__tap_1 TAP_10583 (  );
sky130_fd_sc_hd__tap_1 TAP_10584 (  );
sky130_fd_sc_hd__tap_1 TAP_10585 (  );
sky130_fd_sc_hd__tap_1 TAP_10586 (  );
sky130_fd_sc_hd__tap_1 TAP_10587 (  );
sky130_fd_sc_hd__tap_1 TAP_10588 (  );
sky130_fd_sc_hd__tap_1 TAP_10589 (  );
sky130_fd_sc_hd__tap_1 TAP_1059 (  );
sky130_fd_sc_hd__tap_1 TAP_10590 (  );
sky130_fd_sc_hd__tap_1 TAP_10591 (  );
sky130_fd_sc_hd__tap_1 TAP_10592 (  );
sky130_fd_sc_hd__tap_1 TAP_10593 (  );
sky130_fd_sc_hd__tap_1 TAP_10594 (  );
sky130_fd_sc_hd__tap_1 TAP_10595 (  );
sky130_fd_sc_hd__tap_1 TAP_10596 (  );
sky130_fd_sc_hd__tap_1 TAP_10597 (  );
sky130_fd_sc_hd__tap_1 TAP_10598 (  );
sky130_fd_sc_hd__tap_1 TAP_10599 (  );
sky130_fd_sc_hd__tap_1 TAP_1060 (  );
sky130_fd_sc_hd__tap_1 TAP_10600 (  );
sky130_fd_sc_hd__tap_1 TAP_10601 (  );
sky130_fd_sc_hd__tap_1 TAP_10602 (  );
sky130_fd_sc_hd__tap_1 TAP_10603 (  );
sky130_fd_sc_hd__tap_1 TAP_10604 (  );
sky130_fd_sc_hd__tap_1 TAP_10605 (  );
sky130_fd_sc_hd__tap_1 TAP_10606 (  );
sky130_fd_sc_hd__tap_1 TAP_10607 (  );
sky130_fd_sc_hd__tap_1 TAP_10608 (  );
sky130_fd_sc_hd__tap_1 TAP_10609 (  );
sky130_fd_sc_hd__tap_1 TAP_1061 (  );
sky130_fd_sc_hd__tap_1 TAP_10610 (  );
sky130_fd_sc_hd__tap_1 TAP_10611 (  );
sky130_fd_sc_hd__tap_1 TAP_10612 (  );
sky130_fd_sc_hd__tap_1 TAP_10613 (  );
sky130_fd_sc_hd__tap_1 TAP_10614 (  );
sky130_fd_sc_hd__tap_1 TAP_10615 (  );
sky130_fd_sc_hd__tap_1 TAP_10616 (  );
sky130_fd_sc_hd__tap_1 TAP_10617 (  );
sky130_fd_sc_hd__tap_1 TAP_10618 (  );
sky130_fd_sc_hd__tap_1 TAP_10619 (  );
sky130_fd_sc_hd__tap_1 TAP_1062 (  );
sky130_fd_sc_hd__tap_1 TAP_10620 (  );
sky130_fd_sc_hd__tap_1 TAP_10621 (  );
sky130_fd_sc_hd__tap_1 TAP_10622 (  );
sky130_fd_sc_hd__tap_1 TAP_10623 (  );
sky130_fd_sc_hd__tap_1 TAP_10624 (  );
sky130_fd_sc_hd__tap_1 TAP_10625 (  );
sky130_fd_sc_hd__tap_1 TAP_10626 (  );
sky130_fd_sc_hd__tap_1 TAP_10627 (  );
sky130_fd_sc_hd__tap_1 TAP_10628 (  );
sky130_fd_sc_hd__tap_1 TAP_10629 (  );
sky130_fd_sc_hd__tap_1 TAP_1063 (  );
sky130_fd_sc_hd__tap_1 TAP_10630 (  );
sky130_fd_sc_hd__tap_1 TAP_10631 (  );
sky130_fd_sc_hd__tap_1 TAP_10632 (  );
sky130_fd_sc_hd__tap_1 TAP_10633 (  );
sky130_fd_sc_hd__tap_1 TAP_10634 (  );
sky130_fd_sc_hd__tap_1 TAP_10635 (  );
sky130_fd_sc_hd__tap_1 TAP_10636 (  );
sky130_fd_sc_hd__tap_1 TAP_10637 (  );
sky130_fd_sc_hd__tap_1 TAP_10638 (  );
sky130_fd_sc_hd__tap_1 TAP_10639 (  );
sky130_fd_sc_hd__tap_1 TAP_1064 (  );
sky130_fd_sc_hd__tap_1 TAP_10640 (  );
sky130_fd_sc_hd__tap_1 TAP_10641 (  );
sky130_fd_sc_hd__tap_1 TAP_10642 (  );
sky130_fd_sc_hd__tap_1 TAP_10643 (  );
sky130_fd_sc_hd__tap_1 TAP_10644 (  );
sky130_fd_sc_hd__tap_1 TAP_10645 (  );
sky130_fd_sc_hd__tap_1 TAP_10646 (  );
sky130_fd_sc_hd__tap_1 TAP_10647 (  );
sky130_fd_sc_hd__tap_1 TAP_10648 (  );
sky130_fd_sc_hd__tap_1 TAP_10649 (  );
sky130_fd_sc_hd__tap_1 TAP_1065 (  );
sky130_fd_sc_hd__tap_1 TAP_10650 (  );
sky130_fd_sc_hd__tap_1 TAP_10651 (  );
sky130_fd_sc_hd__tap_1 TAP_10652 (  );
sky130_fd_sc_hd__tap_1 TAP_10653 (  );
sky130_fd_sc_hd__tap_1 TAP_10654 (  );
sky130_fd_sc_hd__tap_1 TAP_10655 (  );
sky130_fd_sc_hd__tap_1 TAP_10656 (  );
sky130_fd_sc_hd__tap_1 TAP_10657 (  );
sky130_fd_sc_hd__tap_1 TAP_10658 (  );
sky130_fd_sc_hd__tap_1 TAP_10659 (  );
sky130_fd_sc_hd__tap_1 TAP_1066 (  );
sky130_fd_sc_hd__tap_1 TAP_10660 (  );
sky130_fd_sc_hd__tap_1 TAP_10661 (  );
sky130_fd_sc_hd__tap_1 TAP_10662 (  );
sky130_fd_sc_hd__tap_1 TAP_10663 (  );
sky130_fd_sc_hd__tap_1 TAP_10664 (  );
sky130_fd_sc_hd__tap_1 TAP_10665 (  );
sky130_fd_sc_hd__tap_1 TAP_10666 (  );
sky130_fd_sc_hd__tap_1 TAP_10667 (  );
sky130_fd_sc_hd__tap_1 TAP_10668 (  );
sky130_fd_sc_hd__tap_1 TAP_10669 (  );
sky130_fd_sc_hd__tap_1 TAP_1067 (  );
sky130_fd_sc_hd__tap_1 TAP_10670 (  );
sky130_fd_sc_hd__tap_1 TAP_10671 (  );
sky130_fd_sc_hd__tap_1 TAP_10672 (  );
sky130_fd_sc_hd__tap_1 TAP_10673 (  );
sky130_fd_sc_hd__tap_1 TAP_10674 (  );
sky130_fd_sc_hd__tap_1 TAP_10675 (  );
sky130_fd_sc_hd__tap_1 TAP_10676 (  );
sky130_fd_sc_hd__tap_1 TAP_10677 (  );
sky130_fd_sc_hd__tap_1 TAP_10678 (  );
sky130_fd_sc_hd__tap_1 TAP_10679 (  );
sky130_fd_sc_hd__tap_1 TAP_1068 (  );
sky130_fd_sc_hd__tap_1 TAP_10680 (  );
sky130_fd_sc_hd__tap_1 TAP_10681 (  );
sky130_fd_sc_hd__tap_1 TAP_10682 (  );
sky130_fd_sc_hd__tap_1 TAP_10683 (  );
sky130_fd_sc_hd__tap_1 TAP_10684 (  );
sky130_fd_sc_hd__tap_1 TAP_10685 (  );
sky130_fd_sc_hd__tap_1 TAP_10686 (  );
sky130_fd_sc_hd__tap_1 TAP_10687 (  );
sky130_fd_sc_hd__tap_1 TAP_10688 (  );
sky130_fd_sc_hd__tap_1 TAP_10689 (  );
sky130_fd_sc_hd__tap_1 TAP_1069 (  );
sky130_fd_sc_hd__tap_1 TAP_10690 (  );
sky130_fd_sc_hd__tap_1 TAP_10691 (  );
sky130_fd_sc_hd__tap_1 TAP_10692 (  );
sky130_fd_sc_hd__tap_1 TAP_10693 (  );
sky130_fd_sc_hd__tap_1 TAP_10694 (  );
sky130_fd_sc_hd__tap_1 TAP_10695 (  );
sky130_fd_sc_hd__tap_1 TAP_10696 (  );
sky130_fd_sc_hd__tap_1 TAP_10697 (  );
sky130_fd_sc_hd__tap_1 TAP_10698 (  );
sky130_fd_sc_hd__tap_1 TAP_10699 (  );
sky130_fd_sc_hd__tap_1 TAP_1070 (  );
sky130_fd_sc_hd__tap_1 TAP_10700 (  );
sky130_fd_sc_hd__tap_1 TAP_10701 (  );
sky130_fd_sc_hd__tap_1 TAP_10702 (  );
sky130_fd_sc_hd__tap_1 TAP_10703 (  );
sky130_fd_sc_hd__tap_1 TAP_10704 (  );
sky130_fd_sc_hd__tap_1 TAP_10705 (  );
sky130_fd_sc_hd__tap_1 TAP_10706 (  );
sky130_fd_sc_hd__tap_1 TAP_10707 (  );
sky130_fd_sc_hd__tap_1 TAP_10708 (  );
sky130_fd_sc_hd__tap_1 TAP_10709 (  );
sky130_fd_sc_hd__tap_1 TAP_1071 (  );
sky130_fd_sc_hd__tap_1 TAP_10710 (  );
sky130_fd_sc_hd__tap_1 TAP_10711 (  );
sky130_fd_sc_hd__tap_1 TAP_10712 (  );
sky130_fd_sc_hd__tap_1 TAP_10713 (  );
sky130_fd_sc_hd__tap_1 TAP_10714 (  );
sky130_fd_sc_hd__tap_1 TAP_10715 (  );
sky130_fd_sc_hd__tap_1 TAP_10716 (  );
sky130_fd_sc_hd__tap_1 TAP_10717 (  );
sky130_fd_sc_hd__tap_1 TAP_10718 (  );
sky130_fd_sc_hd__tap_1 TAP_10719 (  );
sky130_fd_sc_hd__tap_1 TAP_1072 (  );
sky130_fd_sc_hd__tap_1 TAP_10720 (  );
sky130_fd_sc_hd__tap_1 TAP_10721 (  );
sky130_fd_sc_hd__tap_1 TAP_10722 (  );
sky130_fd_sc_hd__tap_1 TAP_10723 (  );
sky130_fd_sc_hd__tap_1 TAP_10724 (  );
sky130_fd_sc_hd__tap_1 TAP_10725 (  );
sky130_fd_sc_hd__tap_1 TAP_10726 (  );
sky130_fd_sc_hd__tap_1 TAP_10727 (  );
sky130_fd_sc_hd__tap_1 TAP_10728 (  );
sky130_fd_sc_hd__tap_1 TAP_10729 (  );
sky130_fd_sc_hd__tap_1 TAP_1073 (  );
sky130_fd_sc_hd__tap_1 TAP_10730 (  );
sky130_fd_sc_hd__tap_1 TAP_10731 (  );
sky130_fd_sc_hd__tap_1 TAP_10732 (  );
sky130_fd_sc_hd__tap_1 TAP_10733 (  );
sky130_fd_sc_hd__tap_1 TAP_10734 (  );
sky130_fd_sc_hd__tap_1 TAP_10735 (  );
sky130_fd_sc_hd__tap_1 TAP_10736 (  );
sky130_fd_sc_hd__tap_1 TAP_10737 (  );
sky130_fd_sc_hd__tap_1 TAP_10738 (  );
sky130_fd_sc_hd__tap_1 TAP_10739 (  );
sky130_fd_sc_hd__tap_1 TAP_1074 (  );
sky130_fd_sc_hd__tap_1 TAP_10740 (  );
sky130_fd_sc_hd__tap_1 TAP_10741 (  );
sky130_fd_sc_hd__tap_1 TAP_10742 (  );
sky130_fd_sc_hd__tap_1 TAP_10743 (  );
sky130_fd_sc_hd__tap_1 TAP_10744 (  );
sky130_fd_sc_hd__tap_1 TAP_10745 (  );
sky130_fd_sc_hd__tap_1 TAP_10746 (  );
sky130_fd_sc_hd__tap_1 TAP_10747 (  );
sky130_fd_sc_hd__tap_1 TAP_10748 (  );
sky130_fd_sc_hd__tap_1 TAP_10749 (  );
sky130_fd_sc_hd__tap_1 TAP_1075 (  );
sky130_fd_sc_hd__tap_1 TAP_10750 (  );
sky130_fd_sc_hd__tap_1 TAP_10751 (  );
sky130_fd_sc_hd__tap_1 TAP_10752 (  );
sky130_fd_sc_hd__tap_1 TAP_10753 (  );
sky130_fd_sc_hd__tap_1 TAP_10754 (  );
sky130_fd_sc_hd__tap_1 TAP_10755 (  );
sky130_fd_sc_hd__tap_1 TAP_10756 (  );
sky130_fd_sc_hd__tap_1 TAP_10757 (  );
sky130_fd_sc_hd__tap_1 TAP_10758 (  );
sky130_fd_sc_hd__tap_1 TAP_10759 (  );
sky130_fd_sc_hd__tap_1 TAP_1076 (  );
sky130_fd_sc_hd__tap_1 TAP_10760 (  );
sky130_fd_sc_hd__tap_1 TAP_10761 (  );
sky130_fd_sc_hd__tap_1 TAP_10762 (  );
sky130_fd_sc_hd__tap_1 TAP_10763 (  );
sky130_fd_sc_hd__tap_1 TAP_10764 (  );
sky130_fd_sc_hd__tap_1 TAP_10765 (  );
sky130_fd_sc_hd__tap_1 TAP_10766 (  );
sky130_fd_sc_hd__tap_1 TAP_10767 (  );
sky130_fd_sc_hd__tap_1 TAP_10768 (  );
sky130_fd_sc_hd__tap_1 TAP_10769 (  );
sky130_fd_sc_hd__tap_1 TAP_1077 (  );
sky130_fd_sc_hd__tap_1 TAP_10770 (  );
sky130_fd_sc_hd__tap_1 TAP_10771 (  );
sky130_fd_sc_hd__tap_1 TAP_10772 (  );
sky130_fd_sc_hd__tap_1 TAP_10773 (  );
sky130_fd_sc_hd__tap_1 TAP_10774 (  );
sky130_fd_sc_hd__tap_1 TAP_10775 (  );
sky130_fd_sc_hd__tap_1 TAP_10776 (  );
sky130_fd_sc_hd__tap_1 TAP_10777 (  );
sky130_fd_sc_hd__tap_1 TAP_10778 (  );
sky130_fd_sc_hd__tap_1 TAP_10779 (  );
sky130_fd_sc_hd__tap_1 TAP_1078 (  );
sky130_fd_sc_hd__tap_1 TAP_10780 (  );
sky130_fd_sc_hd__tap_1 TAP_10781 (  );
sky130_fd_sc_hd__tap_1 TAP_10782 (  );
sky130_fd_sc_hd__tap_1 TAP_10783 (  );
sky130_fd_sc_hd__tap_1 TAP_10784 (  );
sky130_fd_sc_hd__tap_1 TAP_10785 (  );
sky130_fd_sc_hd__tap_1 TAP_10786 (  );
sky130_fd_sc_hd__tap_1 TAP_10787 (  );
sky130_fd_sc_hd__tap_1 TAP_10788 (  );
sky130_fd_sc_hd__tap_1 TAP_10789 (  );
sky130_fd_sc_hd__tap_1 TAP_1079 (  );
sky130_fd_sc_hd__tap_1 TAP_10790 (  );
sky130_fd_sc_hd__tap_1 TAP_10791 (  );
sky130_fd_sc_hd__tap_1 TAP_10792 (  );
sky130_fd_sc_hd__tap_1 TAP_10793 (  );
sky130_fd_sc_hd__tap_1 TAP_10794 (  );
sky130_fd_sc_hd__tap_1 TAP_10795 (  );
sky130_fd_sc_hd__tap_1 TAP_10796 (  );
sky130_fd_sc_hd__tap_1 TAP_10797 (  );
sky130_fd_sc_hd__tap_1 TAP_10798 (  );
sky130_fd_sc_hd__tap_1 TAP_10799 (  );
sky130_fd_sc_hd__tap_1 TAP_1080 (  );
sky130_fd_sc_hd__tap_1 TAP_10800 (  );
sky130_fd_sc_hd__tap_1 TAP_10801 (  );
sky130_fd_sc_hd__tap_1 TAP_10802 (  );
sky130_fd_sc_hd__tap_1 TAP_10803 (  );
sky130_fd_sc_hd__tap_1 TAP_10804 (  );
sky130_fd_sc_hd__tap_1 TAP_10805 (  );
sky130_fd_sc_hd__tap_1 TAP_10806 (  );
sky130_fd_sc_hd__tap_1 TAP_10807 (  );
sky130_fd_sc_hd__tap_1 TAP_10808 (  );
sky130_fd_sc_hd__tap_1 TAP_10809 (  );
sky130_fd_sc_hd__tap_1 TAP_1081 (  );
sky130_fd_sc_hd__tap_1 TAP_10810 (  );
sky130_fd_sc_hd__tap_1 TAP_10811 (  );
sky130_fd_sc_hd__tap_1 TAP_10812 (  );
sky130_fd_sc_hd__tap_1 TAP_10813 (  );
sky130_fd_sc_hd__tap_1 TAP_10814 (  );
sky130_fd_sc_hd__tap_1 TAP_10815 (  );
sky130_fd_sc_hd__tap_1 TAP_10816 (  );
sky130_fd_sc_hd__tap_1 TAP_10817 (  );
sky130_fd_sc_hd__tap_1 TAP_10818 (  );
sky130_fd_sc_hd__tap_1 TAP_10819 (  );
sky130_fd_sc_hd__tap_1 TAP_1082 (  );
sky130_fd_sc_hd__tap_1 TAP_10820 (  );
sky130_fd_sc_hd__tap_1 TAP_10821 (  );
sky130_fd_sc_hd__tap_1 TAP_10822 (  );
sky130_fd_sc_hd__tap_1 TAP_10823 (  );
sky130_fd_sc_hd__tap_1 TAP_10824 (  );
sky130_fd_sc_hd__tap_1 TAP_10825 (  );
sky130_fd_sc_hd__tap_1 TAP_10826 (  );
sky130_fd_sc_hd__tap_1 TAP_10827 (  );
sky130_fd_sc_hd__tap_1 TAP_10828 (  );
sky130_fd_sc_hd__tap_1 TAP_10829 (  );
sky130_fd_sc_hd__tap_1 TAP_1083 (  );
sky130_fd_sc_hd__tap_1 TAP_10830 (  );
sky130_fd_sc_hd__tap_1 TAP_10831 (  );
sky130_fd_sc_hd__tap_1 TAP_10832 (  );
sky130_fd_sc_hd__tap_1 TAP_10833 (  );
sky130_fd_sc_hd__tap_1 TAP_10834 (  );
sky130_fd_sc_hd__tap_1 TAP_10835 (  );
sky130_fd_sc_hd__tap_1 TAP_10836 (  );
sky130_fd_sc_hd__tap_1 TAP_10837 (  );
sky130_fd_sc_hd__tap_1 TAP_10838 (  );
sky130_fd_sc_hd__tap_1 TAP_10839 (  );
sky130_fd_sc_hd__tap_1 TAP_1084 (  );
sky130_fd_sc_hd__tap_1 TAP_10840 (  );
sky130_fd_sc_hd__tap_1 TAP_10841 (  );
sky130_fd_sc_hd__tap_1 TAP_10842 (  );
sky130_fd_sc_hd__tap_1 TAP_10843 (  );
sky130_fd_sc_hd__tap_1 TAP_10844 (  );
sky130_fd_sc_hd__tap_1 TAP_10845 (  );
sky130_fd_sc_hd__tap_1 TAP_10846 (  );
sky130_fd_sc_hd__tap_1 TAP_10847 (  );
sky130_fd_sc_hd__tap_1 TAP_10848 (  );
sky130_fd_sc_hd__tap_1 TAP_10849 (  );
sky130_fd_sc_hd__tap_1 TAP_1085 (  );
sky130_fd_sc_hd__tap_1 TAP_10850 (  );
sky130_fd_sc_hd__tap_1 TAP_10851 (  );
sky130_fd_sc_hd__tap_1 TAP_10852 (  );
sky130_fd_sc_hd__tap_1 TAP_10853 (  );
sky130_fd_sc_hd__tap_1 TAP_10854 (  );
sky130_fd_sc_hd__tap_1 TAP_10855 (  );
sky130_fd_sc_hd__tap_1 TAP_10856 (  );
sky130_fd_sc_hd__tap_1 TAP_10857 (  );
sky130_fd_sc_hd__tap_1 TAP_10858 (  );
sky130_fd_sc_hd__tap_1 TAP_10859 (  );
sky130_fd_sc_hd__tap_1 TAP_1086 (  );
sky130_fd_sc_hd__tap_1 TAP_10860 (  );
sky130_fd_sc_hd__tap_1 TAP_10861 (  );
sky130_fd_sc_hd__tap_1 TAP_10862 (  );
sky130_fd_sc_hd__tap_1 TAP_10863 (  );
sky130_fd_sc_hd__tap_1 TAP_10864 (  );
sky130_fd_sc_hd__tap_1 TAP_10865 (  );
sky130_fd_sc_hd__tap_1 TAP_10866 (  );
sky130_fd_sc_hd__tap_1 TAP_10867 (  );
sky130_fd_sc_hd__tap_1 TAP_10868 (  );
sky130_fd_sc_hd__tap_1 TAP_10869 (  );
sky130_fd_sc_hd__tap_1 TAP_1087 (  );
sky130_fd_sc_hd__tap_1 TAP_10870 (  );
sky130_fd_sc_hd__tap_1 TAP_10871 (  );
sky130_fd_sc_hd__tap_1 TAP_10872 (  );
sky130_fd_sc_hd__tap_1 TAP_10873 (  );
sky130_fd_sc_hd__tap_1 TAP_10874 (  );
sky130_fd_sc_hd__tap_1 TAP_10875 (  );
sky130_fd_sc_hd__tap_1 TAP_10876 (  );
sky130_fd_sc_hd__tap_1 TAP_10877 (  );
sky130_fd_sc_hd__tap_1 TAP_10878 (  );
sky130_fd_sc_hd__tap_1 TAP_10879 (  );
sky130_fd_sc_hd__tap_1 TAP_1088 (  );
sky130_fd_sc_hd__tap_1 TAP_10880 (  );
sky130_fd_sc_hd__tap_1 TAP_10881 (  );
sky130_fd_sc_hd__tap_1 TAP_10882 (  );
sky130_fd_sc_hd__tap_1 TAP_10883 (  );
sky130_fd_sc_hd__tap_1 TAP_10884 (  );
sky130_fd_sc_hd__tap_1 TAP_10885 (  );
sky130_fd_sc_hd__tap_1 TAP_10886 (  );
sky130_fd_sc_hd__tap_1 TAP_10887 (  );
sky130_fd_sc_hd__tap_1 TAP_10888 (  );
sky130_fd_sc_hd__tap_1 TAP_10889 (  );
sky130_fd_sc_hd__tap_1 TAP_1089 (  );
sky130_fd_sc_hd__tap_1 TAP_10890 (  );
sky130_fd_sc_hd__tap_1 TAP_10891 (  );
sky130_fd_sc_hd__tap_1 TAP_10892 (  );
sky130_fd_sc_hd__tap_1 TAP_10893 (  );
sky130_fd_sc_hd__tap_1 TAP_10894 (  );
sky130_fd_sc_hd__tap_1 TAP_10895 (  );
sky130_fd_sc_hd__tap_1 TAP_10896 (  );
sky130_fd_sc_hd__tap_1 TAP_10897 (  );
sky130_fd_sc_hd__tap_1 TAP_10898 (  );
sky130_fd_sc_hd__tap_1 TAP_10899 (  );
sky130_fd_sc_hd__tap_1 TAP_1090 (  );
sky130_fd_sc_hd__tap_1 TAP_10900 (  );
sky130_fd_sc_hd__tap_1 TAP_10901 (  );
sky130_fd_sc_hd__tap_1 TAP_10902 (  );
sky130_fd_sc_hd__tap_1 TAP_10903 (  );
sky130_fd_sc_hd__tap_1 TAP_10904 (  );
sky130_fd_sc_hd__tap_1 TAP_10905 (  );
sky130_fd_sc_hd__tap_1 TAP_10906 (  );
sky130_fd_sc_hd__tap_1 TAP_10907 (  );
sky130_fd_sc_hd__tap_1 TAP_10908 (  );
sky130_fd_sc_hd__tap_1 TAP_10909 (  );
sky130_fd_sc_hd__tap_1 TAP_1091 (  );
sky130_fd_sc_hd__tap_1 TAP_10910 (  );
sky130_fd_sc_hd__tap_1 TAP_10911 (  );
sky130_fd_sc_hd__tap_1 TAP_10912 (  );
sky130_fd_sc_hd__tap_1 TAP_10913 (  );
sky130_fd_sc_hd__tap_1 TAP_10914 (  );
sky130_fd_sc_hd__tap_1 TAP_10915 (  );
sky130_fd_sc_hd__tap_1 TAP_10916 (  );
sky130_fd_sc_hd__tap_1 TAP_10917 (  );
sky130_fd_sc_hd__tap_1 TAP_10918 (  );
sky130_fd_sc_hd__tap_1 TAP_10919 (  );
sky130_fd_sc_hd__tap_1 TAP_1092 (  );
sky130_fd_sc_hd__tap_1 TAP_10920 (  );
sky130_fd_sc_hd__tap_1 TAP_10921 (  );
sky130_fd_sc_hd__tap_1 TAP_10922 (  );
sky130_fd_sc_hd__tap_1 TAP_10923 (  );
sky130_fd_sc_hd__tap_1 TAP_10924 (  );
sky130_fd_sc_hd__tap_1 TAP_10925 (  );
sky130_fd_sc_hd__tap_1 TAP_10926 (  );
sky130_fd_sc_hd__tap_1 TAP_10927 (  );
sky130_fd_sc_hd__tap_1 TAP_10928 (  );
sky130_fd_sc_hd__tap_1 TAP_10929 (  );
sky130_fd_sc_hd__tap_1 TAP_1093 (  );
sky130_fd_sc_hd__tap_1 TAP_10930 (  );
sky130_fd_sc_hd__tap_1 TAP_10931 (  );
sky130_fd_sc_hd__tap_1 TAP_10932 (  );
sky130_fd_sc_hd__tap_1 TAP_10933 (  );
sky130_fd_sc_hd__tap_1 TAP_10934 (  );
sky130_fd_sc_hd__tap_1 TAP_10935 (  );
sky130_fd_sc_hd__tap_1 TAP_10936 (  );
sky130_fd_sc_hd__tap_1 TAP_10937 (  );
sky130_fd_sc_hd__tap_1 TAP_10938 (  );
sky130_fd_sc_hd__tap_1 TAP_10939 (  );
sky130_fd_sc_hd__tap_1 TAP_1094 (  );
sky130_fd_sc_hd__tap_1 TAP_10940 (  );
sky130_fd_sc_hd__tap_1 TAP_10941 (  );
sky130_fd_sc_hd__tap_1 TAP_10942 (  );
sky130_fd_sc_hd__tap_1 TAP_10943 (  );
sky130_fd_sc_hd__tap_1 TAP_10944 (  );
sky130_fd_sc_hd__tap_1 TAP_10945 (  );
sky130_fd_sc_hd__tap_1 TAP_10946 (  );
sky130_fd_sc_hd__tap_1 TAP_10947 (  );
sky130_fd_sc_hd__tap_1 TAP_10948 (  );
sky130_fd_sc_hd__tap_1 TAP_10949 (  );
sky130_fd_sc_hd__tap_1 TAP_1095 (  );
sky130_fd_sc_hd__tap_1 TAP_10950 (  );
sky130_fd_sc_hd__tap_1 TAP_10951 (  );
sky130_fd_sc_hd__tap_1 TAP_10952 (  );
sky130_fd_sc_hd__tap_1 TAP_10953 (  );
sky130_fd_sc_hd__tap_1 TAP_10954 (  );
sky130_fd_sc_hd__tap_1 TAP_10955 (  );
sky130_fd_sc_hd__tap_1 TAP_10956 (  );
sky130_fd_sc_hd__tap_1 TAP_10957 (  );
sky130_fd_sc_hd__tap_1 TAP_10958 (  );
sky130_fd_sc_hd__tap_1 TAP_10959 (  );
sky130_fd_sc_hd__tap_1 TAP_1096 (  );
sky130_fd_sc_hd__tap_1 TAP_10960 (  );
sky130_fd_sc_hd__tap_1 TAP_10961 (  );
sky130_fd_sc_hd__tap_1 TAP_10962 (  );
sky130_fd_sc_hd__tap_1 TAP_10963 (  );
sky130_fd_sc_hd__tap_1 TAP_10964 (  );
sky130_fd_sc_hd__tap_1 TAP_10965 (  );
sky130_fd_sc_hd__tap_1 TAP_10966 (  );
sky130_fd_sc_hd__tap_1 TAP_10967 (  );
sky130_fd_sc_hd__tap_1 TAP_10968 (  );
sky130_fd_sc_hd__tap_1 TAP_10969 (  );
sky130_fd_sc_hd__tap_1 TAP_1097 (  );
sky130_fd_sc_hd__tap_1 TAP_10970 (  );
sky130_fd_sc_hd__tap_1 TAP_10971 (  );
sky130_fd_sc_hd__tap_1 TAP_10972 (  );
sky130_fd_sc_hd__tap_1 TAP_10973 (  );
sky130_fd_sc_hd__tap_1 TAP_10974 (  );
sky130_fd_sc_hd__tap_1 TAP_10975 (  );
sky130_fd_sc_hd__tap_1 TAP_10976 (  );
sky130_fd_sc_hd__tap_1 TAP_10977 (  );
sky130_fd_sc_hd__tap_1 TAP_10978 (  );
sky130_fd_sc_hd__tap_1 TAP_10979 (  );
sky130_fd_sc_hd__tap_1 TAP_1098 (  );
sky130_fd_sc_hd__tap_1 TAP_10980 (  );
sky130_fd_sc_hd__tap_1 TAP_10981 (  );
sky130_fd_sc_hd__tap_1 TAP_10982 (  );
sky130_fd_sc_hd__tap_1 TAP_10983 (  );
sky130_fd_sc_hd__tap_1 TAP_10984 (  );
sky130_fd_sc_hd__tap_1 TAP_10985 (  );
sky130_fd_sc_hd__tap_1 TAP_10986 (  );
sky130_fd_sc_hd__tap_1 TAP_10987 (  );
sky130_fd_sc_hd__tap_1 TAP_10988 (  );
sky130_fd_sc_hd__tap_1 TAP_10989 (  );
sky130_fd_sc_hd__tap_1 TAP_1099 (  );
sky130_fd_sc_hd__tap_1 TAP_10990 (  );
sky130_fd_sc_hd__tap_1 TAP_10991 (  );
sky130_fd_sc_hd__tap_1 TAP_10992 (  );
sky130_fd_sc_hd__tap_1 TAP_10993 (  );
sky130_fd_sc_hd__tap_1 TAP_10994 (  );
sky130_fd_sc_hd__tap_1 TAP_10995 (  );
sky130_fd_sc_hd__tap_1 TAP_10996 (  );
sky130_fd_sc_hd__tap_1 TAP_10997 (  );
sky130_fd_sc_hd__tap_1 TAP_10998 (  );
sky130_fd_sc_hd__tap_1 TAP_10999 (  );
sky130_fd_sc_hd__tap_1 TAP_1100 (  );
sky130_fd_sc_hd__tap_1 TAP_11000 (  );
sky130_fd_sc_hd__tap_1 TAP_11001 (  );
sky130_fd_sc_hd__tap_1 TAP_11002 (  );
sky130_fd_sc_hd__tap_1 TAP_11003 (  );
sky130_fd_sc_hd__tap_1 TAP_11004 (  );
sky130_fd_sc_hd__tap_1 TAP_11005 (  );
sky130_fd_sc_hd__tap_1 TAP_11006 (  );
sky130_fd_sc_hd__tap_1 TAP_11007 (  );
sky130_fd_sc_hd__tap_1 TAP_11008 (  );
sky130_fd_sc_hd__tap_1 TAP_11009 (  );
sky130_fd_sc_hd__tap_1 TAP_1101 (  );
sky130_fd_sc_hd__tap_1 TAP_11010 (  );
sky130_fd_sc_hd__tap_1 TAP_11011 (  );
sky130_fd_sc_hd__tap_1 TAP_11012 (  );
sky130_fd_sc_hd__tap_1 TAP_11013 (  );
sky130_fd_sc_hd__tap_1 TAP_11014 (  );
sky130_fd_sc_hd__tap_1 TAP_11015 (  );
sky130_fd_sc_hd__tap_1 TAP_11016 (  );
sky130_fd_sc_hd__tap_1 TAP_11017 (  );
sky130_fd_sc_hd__tap_1 TAP_11018 (  );
sky130_fd_sc_hd__tap_1 TAP_11019 (  );
sky130_fd_sc_hd__tap_1 TAP_1102 (  );
sky130_fd_sc_hd__tap_1 TAP_11020 (  );
sky130_fd_sc_hd__tap_1 TAP_11021 (  );
sky130_fd_sc_hd__tap_1 TAP_11022 (  );
sky130_fd_sc_hd__tap_1 TAP_11023 (  );
sky130_fd_sc_hd__tap_1 TAP_11024 (  );
sky130_fd_sc_hd__tap_1 TAP_11025 (  );
sky130_fd_sc_hd__tap_1 TAP_11026 (  );
sky130_fd_sc_hd__tap_1 TAP_11027 (  );
sky130_fd_sc_hd__tap_1 TAP_11028 (  );
sky130_fd_sc_hd__tap_1 TAP_11029 (  );
sky130_fd_sc_hd__tap_1 TAP_1103 (  );
sky130_fd_sc_hd__tap_1 TAP_11030 (  );
sky130_fd_sc_hd__tap_1 TAP_11031 (  );
sky130_fd_sc_hd__tap_1 TAP_11032 (  );
sky130_fd_sc_hd__tap_1 TAP_11033 (  );
sky130_fd_sc_hd__tap_1 TAP_11034 (  );
sky130_fd_sc_hd__tap_1 TAP_11035 (  );
sky130_fd_sc_hd__tap_1 TAP_11036 (  );
sky130_fd_sc_hd__tap_1 TAP_11037 (  );
sky130_fd_sc_hd__tap_1 TAP_11038 (  );
sky130_fd_sc_hd__tap_1 TAP_11039 (  );
sky130_fd_sc_hd__tap_1 TAP_1104 (  );
sky130_fd_sc_hd__tap_1 TAP_11040 (  );
sky130_fd_sc_hd__tap_1 TAP_11041 (  );
sky130_fd_sc_hd__tap_1 TAP_11042 (  );
sky130_fd_sc_hd__tap_1 TAP_11043 (  );
sky130_fd_sc_hd__tap_1 TAP_11044 (  );
sky130_fd_sc_hd__tap_1 TAP_11045 (  );
sky130_fd_sc_hd__tap_1 TAP_11046 (  );
sky130_fd_sc_hd__tap_1 TAP_11047 (  );
sky130_fd_sc_hd__tap_1 TAP_11048 (  );
sky130_fd_sc_hd__tap_1 TAP_11049 (  );
sky130_fd_sc_hd__tap_1 TAP_1105 (  );
sky130_fd_sc_hd__tap_1 TAP_11050 (  );
sky130_fd_sc_hd__tap_1 TAP_11051 (  );
sky130_fd_sc_hd__tap_1 TAP_11052 (  );
sky130_fd_sc_hd__tap_1 TAP_11053 (  );
sky130_fd_sc_hd__tap_1 TAP_11054 (  );
sky130_fd_sc_hd__tap_1 TAP_11055 (  );
sky130_fd_sc_hd__tap_1 TAP_11056 (  );
sky130_fd_sc_hd__tap_1 TAP_11057 (  );
sky130_fd_sc_hd__tap_1 TAP_11058 (  );
sky130_fd_sc_hd__tap_1 TAP_11059 (  );
sky130_fd_sc_hd__tap_1 TAP_1106 (  );
sky130_fd_sc_hd__tap_1 TAP_11060 (  );
sky130_fd_sc_hd__tap_1 TAP_11061 (  );
sky130_fd_sc_hd__tap_1 TAP_11062 (  );
sky130_fd_sc_hd__tap_1 TAP_11063 (  );
sky130_fd_sc_hd__tap_1 TAP_11064 (  );
sky130_fd_sc_hd__tap_1 TAP_11065 (  );
sky130_fd_sc_hd__tap_1 TAP_11066 (  );
sky130_fd_sc_hd__tap_1 TAP_11067 (  );
sky130_fd_sc_hd__tap_1 TAP_11068 (  );
sky130_fd_sc_hd__tap_1 TAP_11069 (  );
sky130_fd_sc_hd__tap_1 TAP_1107 (  );
sky130_fd_sc_hd__tap_1 TAP_11070 (  );
sky130_fd_sc_hd__tap_1 TAP_11071 (  );
sky130_fd_sc_hd__tap_1 TAP_11072 (  );
sky130_fd_sc_hd__tap_1 TAP_11073 (  );
sky130_fd_sc_hd__tap_1 TAP_11074 (  );
sky130_fd_sc_hd__tap_1 TAP_11075 (  );
sky130_fd_sc_hd__tap_1 TAP_11076 (  );
sky130_fd_sc_hd__tap_1 TAP_11077 (  );
sky130_fd_sc_hd__tap_1 TAP_11078 (  );
sky130_fd_sc_hd__tap_1 TAP_11079 (  );
sky130_fd_sc_hd__tap_1 TAP_1108 (  );
sky130_fd_sc_hd__tap_1 TAP_11080 (  );
sky130_fd_sc_hd__tap_1 TAP_11081 (  );
sky130_fd_sc_hd__tap_1 TAP_11082 (  );
sky130_fd_sc_hd__tap_1 TAP_11083 (  );
sky130_fd_sc_hd__tap_1 TAP_11084 (  );
sky130_fd_sc_hd__tap_1 TAP_11085 (  );
sky130_fd_sc_hd__tap_1 TAP_11086 (  );
sky130_fd_sc_hd__tap_1 TAP_11087 (  );
sky130_fd_sc_hd__tap_1 TAP_11088 (  );
sky130_fd_sc_hd__tap_1 TAP_11089 (  );
sky130_fd_sc_hd__tap_1 TAP_1109 (  );
sky130_fd_sc_hd__tap_1 TAP_11090 (  );
sky130_fd_sc_hd__tap_1 TAP_11091 (  );
sky130_fd_sc_hd__tap_1 TAP_11092 (  );
sky130_fd_sc_hd__tap_1 TAP_11093 (  );
sky130_fd_sc_hd__tap_1 TAP_11094 (  );
sky130_fd_sc_hd__tap_1 TAP_11095 (  );
sky130_fd_sc_hd__tap_1 TAP_11096 (  );
sky130_fd_sc_hd__tap_1 TAP_11097 (  );
sky130_fd_sc_hd__tap_1 TAP_11098 (  );
sky130_fd_sc_hd__tap_1 TAP_11099 (  );
sky130_fd_sc_hd__tap_1 TAP_1110 (  );
sky130_fd_sc_hd__tap_1 TAP_11100 (  );
sky130_fd_sc_hd__tap_1 TAP_11101 (  );
sky130_fd_sc_hd__tap_1 TAP_11102 (  );
sky130_fd_sc_hd__tap_1 TAP_11103 (  );
sky130_fd_sc_hd__tap_1 TAP_11104 (  );
sky130_fd_sc_hd__tap_1 TAP_11105 (  );
sky130_fd_sc_hd__tap_1 TAP_11106 (  );
sky130_fd_sc_hd__tap_1 TAP_11107 (  );
sky130_fd_sc_hd__tap_1 TAP_11108 (  );
sky130_fd_sc_hd__tap_1 TAP_11109 (  );
sky130_fd_sc_hd__tap_1 TAP_1111 (  );
sky130_fd_sc_hd__tap_1 TAP_11110 (  );
sky130_fd_sc_hd__tap_1 TAP_11111 (  );
sky130_fd_sc_hd__tap_1 TAP_11112 (  );
sky130_fd_sc_hd__tap_1 TAP_11113 (  );
sky130_fd_sc_hd__tap_1 TAP_11114 (  );
sky130_fd_sc_hd__tap_1 TAP_11115 (  );
sky130_fd_sc_hd__tap_1 TAP_11116 (  );
sky130_fd_sc_hd__tap_1 TAP_11117 (  );
sky130_fd_sc_hd__tap_1 TAP_11118 (  );
sky130_fd_sc_hd__tap_1 TAP_11119 (  );
sky130_fd_sc_hd__tap_1 TAP_1112 (  );
sky130_fd_sc_hd__tap_1 TAP_11120 (  );
sky130_fd_sc_hd__tap_1 TAP_11121 (  );
sky130_fd_sc_hd__tap_1 TAP_11122 (  );
sky130_fd_sc_hd__tap_1 TAP_11123 (  );
sky130_fd_sc_hd__tap_1 TAP_11124 (  );
sky130_fd_sc_hd__tap_1 TAP_11125 (  );
sky130_fd_sc_hd__tap_1 TAP_11126 (  );
sky130_fd_sc_hd__tap_1 TAP_11127 (  );
sky130_fd_sc_hd__tap_1 TAP_11128 (  );
sky130_fd_sc_hd__tap_1 TAP_11129 (  );
sky130_fd_sc_hd__tap_1 TAP_1113 (  );
sky130_fd_sc_hd__tap_1 TAP_11130 (  );
sky130_fd_sc_hd__tap_1 TAP_11131 (  );
sky130_fd_sc_hd__tap_1 TAP_11132 (  );
sky130_fd_sc_hd__tap_1 TAP_11133 (  );
sky130_fd_sc_hd__tap_1 TAP_11134 (  );
sky130_fd_sc_hd__tap_1 TAP_11135 (  );
sky130_fd_sc_hd__tap_1 TAP_11136 (  );
sky130_fd_sc_hd__tap_1 TAP_11137 (  );
sky130_fd_sc_hd__tap_1 TAP_11138 (  );
sky130_fd_sc_hd__tap_1 TAP_11139 (  );
sky130_fd_sc_hd__tap_1 TAP_1114 (  );
sky130_fd_sc_hd__tap_1 TAP_11140 (  );
sky130_fd_sc_hd__tap_1 TAP_11141 (  );
sky130_fd_sc_hd__tap_1 TAP_11142 (  );
sky130_fd_sc_hd__tap_1 TAP_11143 (  );
sky130_fd_sc_hd__tap_1 TAP_11144 (  );
sky130_fd_sc_hd__tap_1 TAP_11145 (  );
sky130_fd_sc_hd__tap_1 TAP_11146 (  );
sky130_fd_sc_hd__tap_1 TAP_11147 (  );
sky130_fd_sc_hd__tap_1 TAP_11148 (  );
sky130_fd_sc_hd__tap_1 TAP_11149 (  );
sky130_fd_sc_hd__tap_1 TAP_1115 (  );
sky130_fd_sc_hd__tap_1 TAP_11150 (  );
sky130_fd_sc_hd__tap_1 TAP_11151 (  );
sky130_fd_sc_hd__tap_1 TAP_11152 (  );
sky130_fd_sc_hd__tap_1 TAP_11153 (  );
sky130_fd_sc_hd__tap_1 TAP_11154 (  );
sky130_fd_sc_hd__tap_1 TAP_11155 (  );
sky130_fd_sc_hd__tap_1 TAP_11156 (  );
sky130_fd_sc_hd__tap_1 TAP_11157 (  );
sky130_fd_sc_hd__tap_1 TAP_11158 (  );
sky130_fd_sc_hd__tap_1 TAP_11159 (  );
sky130_fd_sc_hd__tap_1 TAP_1116 (  );
sky130_fd_sc_hd__tap_1 TAP_11160 (  );
sky130_fd_sc_hd__tap_1 TAP_11161 (  );
sky130_fd_sc_hd__tap_1 TAP_11162 (  );
sky130_fd_sc_hd__tap_1 TAP_11163 (  );
sky130_fd_sc_hd__tap_1 TAP_11164 (  );
sky130_fd_sc_hd__tap_1 TAP_11165 (  );
sky130_fd_sc_hd__tap_1 TAP_11166 (  );
sky130_fd_sc_hd__tap_1 TAP_11167 (  );
sky130_fd_sc_hd__tap_1 TAP_11168 (  );
sky130_fd_sc_hd__tap_1 TAP_11169 (  );
sky130_fd_sc_hd__tap_1 TAP_1117 (  );
sky130_fd_sc_hd__tap_1 TAP_11170 (  );
sky130_fd_sc_hd__tap_1 TAP_11171 (  );
sky130_fd_sc_hd__tap_1 TAP_11172 (  );
sky130_fd_sc_hd__tap_1 TAP_11173 (  );
sky130_fd_sc_hd__tap_1 TAP_11174 (  );
sky130_fd_sc_hd__tap_1 TAP_11175 (  );
sky130_fd_sc_hd__tap_1 TAP_11176 (  );
sky130_fd_sc_hd__tap_1 TAP_11177 (  );
sky130_fd_sc_hd__tap_1 TAP_11178 (  );
sky130_fd_sc_hd__tap_1 TAP_11179 (  );
sky130_fd_sc_hd__tap_1 TAP_1118 (  );
sky130_fd_sc_hd__tap_1 TAP_11180 (  );
sky130_fd_sc_hd__tap_1 TAP_11181 (  );
sky130_fd_sc_hd__tap_1 TAP_11182 (  );
sky130_fd_sc_hd__tap_1 TAP_11183 (  );
sky130_fd_sc_hd__tap_1 TAP_11184 (  );
sky130_fd_sc_hd__tap_1 TAP_11185 (  );
sky130_fd_sc_hd__tap_1 TAP_11186 (  );
sky130_fd_sc_hd__tap_1 TAP_11187 (  );
sky130_fd_sc_hd__tap_1 TAP_11188 (  );
sky130_fd_sc_hd__tap_1 TAP_11189 (  );
sky130_fd_sc_hd__tap_1 TAP_1119 (  );
sky130_fd_sc_hd__tap_1 TAP_11190 (  );
sky130_fd_sc_hd__tap_1 TAP_11191 (  );
sky130_fd_sc_hd__tap_1 TAP_11192 (  );
sky130_fd_sc_hd__tap_1 TAP_11193 (  );
sky130_fd_sc_hd__tap_1 TAP_11194 (  );
sky130_fd_sc_hd__tap_1 TAP_11195 (  );
sky130_fd_sc_hd__tap_1 TAP_11196 (  );
sky130_fd_sc_hd__tap_1 TAP_11197 (  );
sky130_fd_sc_hd__tap_1 TAP_11198 (  );
sky130_fd_sc_hd__tap_1 TAP_11199 (  );
sky130_fd_sc_hd__tap_1 TAP_1120 (  );
sky130_fd_sc_hd__tap_1 TAP_11200 (  );
sky130_fd_sc_hd__tap_1 TAP_11201 (  );
sky130_fd_sc_hd__tap_1 TAP_11202 (  );
sky130_fd_sc_hd__tap_1 TAP_11203 (  );
sky130_fd_sc_hd__tap_1 TAP_11204 (  );
sky130_fd_sc_hd__tap_1 TAP_11205 (  );
sky130_fd_sc_hd__tap_1 TAP_11206 (  );
sky130_fd_sc_hd__tap_1 TAP_11207 (  );
sky130_fd_sc_hd__tap_1 TAP_11208 (  );
sky130_fd_sc_hd__tap_1 TAP_11209 (  );
sky130_fd_sc_hd__tap_1 TAP_1121 (  );
sky130_fd_sc_hd__tap_1 TAP_11210 (  );
sky130_fd_sc_hd__tap_1 TAP_11211 (  );
sky130_fd_sc_hd__tap_1 TAP_11212 (  );
sky130_fd_sc_hd__tap_1 TAP_11213 (  );
sky130_fd_sc_hd__tap_1 TAP_11214 (  );
sky130_fd_sc_hd__tap_1 TAP_11215 (  );
sky130_fd_sc_hd__tap_1 TAP_11216 (  );
sky130_fd_sc_hd__tap_1 TAP_11217 (  );
sky130_fd_sc_hd__tap_1 TAP_11218 (  );
sky130_fd_sc_hd__tap_1 TAP_11219 (  );
sky130_fd_sc_hd__tap_1 TAP_1122 (  );
sky130_fd_sc_hd__tap_1 TAP_11220 (  );
sky130_fd_sc_hd__tap_1 TAP_11221 (  );
sky130_fd_sc_hd__tap_1 TAP_11222 (  );
sky130_fd_sc_hd__tap_1 TAP_11223 (  );
sky130_fd_sc_hd__tap_1 TAP_11224 (  );
sky130_fd_sc_hd__tap_1 TAP_11225 (  );
sky130_fd_sc_hd__tap_1 TAP_11226 (  );
sky130_fd_sc_hd__tap_1 TAP_11227 (  );
sky130_fd_sc_hd__tap_1 TAP_11228 (  );
sky130_fd_sc_hd__tap_1 TAP_11229 (  );
sky130_fd_sc_hd__tap_1 TAP_1123 (  );
sky130_fd_sc_hd__tap_1 TAP_11230 (  );
sky130_fd_sc_hd__tap_1 TAP_11231 (  );
sky130_fd_sc_hd__tap_1 TAP_11232 (  );
sky130_fd_sc_hd__tap_1 TAP_11233 (  );
sky130_fd_sc_hd__tap_1 TAP_11234 (  );
sky130_fd_sc_hd__tap_1 TAP_11235 (  );
sky130_fd_sc_hd__tap_1 TAP_11236 (  );
sky130_fd_sc_hd__tap_1 TAP_11237 (  );
sky130_fd_sc_hd__tap_1 TAP_11238 (  );
sky130_fd_sc_hd__tap_1 TAP_11239 (  );
sky130_fd_sc_hd__tap_1 TAP_1124 (  );
sky130_fd_sc_hd__tap_1 TAP_11240 (  );
sky130_fd_sc_hd__tap_1 TAP_11241 (  );
sky130_fd_sc_hd__tap_1 TAP_11242 (  );
sky130_fd_sc_hd__tap_1 TAP_11243 (  );
sky130_fd_sc_hd__tap_1 TAP_11244 (  );
sky130_fd_sc_hd__tap_1 TAP_11245 (  );
sky130_fd_sc_hd__tap_1 TAP_11246 (  );
sky130_fd_sc_hd__tap_1 TAP_11247 (  );
sky130_fd_sc_hd__tap_1 TAP_11248 (  );
sky130_fd_sc_hd__tap_1 TAP_11249 (  );
sky130_fd_sc_hd__tap_1 TAP_1125 (  );
sky130_fd_sc_hd__tap_1 TAP_11250 (  );
sky130_fd_sc_hd__tap_1 TAP_11251 (  );
sky130_fd_sc_hd__tap_1 TAP_11252 (  );
sky130_fd_sc_hd__tap_1 TAP_11253 (  );
sky130_fd_sc_hd__tap_1 TAP_11254 (  );
sky130_fd_sc_hd__tap_1 TAP_11255 (  );
sky130_fd_sc_hd__tap_1 TAP_11256 (  );
sky130_fd_sc_hd__tap_1 TAP_11257 (  );
sky130_fd_sc_hd__tap_1 TAP_11258 (  );
sky130_fd_sc_hd__tap_1 TAP_11259 (  );
sky130_fd_sc_hd__tap_1 TAP_1126 (  );
sky130_fd_sc_hd__tap_1 TAP_11260 (  );
sky130_fd_sc_hd__tap_1 TAP_11261 (  );
sky130_fd_sc_hd__tap_1 TAP_11262 (  );
sky130_fd_sc_hd__tap_1 TAP_11263 (  );
sky130_fd_sc_hd__tap_1 TAP_11264 (  );
sky130_fd_sc_hd__tap_1 TAP_11265 (  );
sky130_fd_sc_hd__tap_1 TAP_11266 (  );
sky130_fd_sc_hd__tap_1 TAP_11267 (  );
sky130_fd_sc_hd__tap_1 TAP_11268 (  );
sky130_fd_sc_hd__tap_1 TAP_11269 (  );
sky130_fd_sc_hd__tap_1 TAP_1127 (  );
sky130_fd_sc_hd__tap_1 TAP_11270 (  );
sky130_fd_sc_hd__tap_1 TAP_11271 (  );
sky130_fd_sc_hd__tap_1 TAP_11272 (  );
sky130_fd_sc_hd__tap_1 TAP_11273 (  );
sky130_fd_sc_hd__tap_1 TAP_11274 (  );
sky130_fd_sc_hd__tap_1 TAP_11275 (  );
sky130_fd_sc_hd__tap_1 TAP_11276 (  );
sky130_fd_sc_hd__tap_1 TAP_11277 (  );
sky130_fd_sc_hd__tap_1 TAP_11278 (  );
sky130_fd_sc_hd__tap_1 TAP_11279 (  );
sky130_fd_sc_hd__tap_1 TAP_1128 (  );
sky130_fd_sc_hd__tap_1 TAP_11280 (  );
sky130_fd_sc_hd__tap_1 TAP_11281 (  );
sky130_fd_sc_hd__tap_1 TAP_11282 (  );
sky130_fd_sc_hd__tap_1 TAP_11283 (  );
sky130_fd_sc_hd__tap_1 TAP_11284 (  );
sky130_fd_sc_hd__tap_1 TAP_11285 (  );
sky130_fd_sc_hd__tap_1 TAP_11286 (  );
sky130_fd_sc_hd__tap_1 TAP_11287 (  );
sky130_fd_sc_hd__tap_1 TAP_11288 (  );
sky130_fd_sc_hd__tap_1 TAP_11289 (  );
sky130_fd_sc_hd__tap_1 TAP_1129 (  );
sky130_fd_sc_hd__tap_1 TAP_11290 (  );
sky130_fd_sc_hd__tap_1 TAP_11291 (  );
sky130_fd_sc_hd__tap_1 TAP_11292 (  );
sky130_fd_sc_hd__tap_1 TAP_11293 (  );
sky130_fd_sc_hd__tap_1 TAP_11294 (  );
sky130_fd_sc_hd__tap_1 TAP_11295 (  );
sky130_fd_sc_hd__tap_1 TAP_11296 (  );
sky130_fd_sc_hd__tap_1 TAP_11297 (  );
sky130_fd_sc_hd__tap_1 TAP_11298 (  );
sky130_fd_sc_hd__tap_1 TAP_11299 (  );
sky130_fd_sc_hd__tap_1 TAP_1130 (  );
sky130_fd_sc_hd__tap_1 TAP_11300 (  );
sky130_fd_sc_hd__tap_1 TAP_11301 (  );
sky130_fd_sc_hd__tap_1 TAP_11302 (  );
sky130_fd_sc_hd__tap_1 TAP_11303 (  );
sky130_fd_sc_hd__tap_1 TAP_11304 (  );
sky130_fd_sc_hd__tap_1 TAP_11305 (  );
sky130_fd_sc_hd__tap_1 TAP_11306 (  );
sky130_fd_sc_hd__tap_1 TAP_11307 (  );
sky130_fd_sc_hd__tap_1 TAP_11308 (  );
sky130_fd_sc_hd__tap_1 TAP_11309 (  );
sky130_fd_sc_hd__tap_1 TAP_1131 (  );
sky130_fd_sc_hd__tap_1 TAP_11310 (  );
sky130_fd_sc_hd__tap_1 TAP_11311 (  );
sky130_fd_sc_hd__tap_1 TAP_11312 (  );
sky130_fd_sc_hd__tap_1 TAP_11313 (  );
sky130_fd_sc_hd__tap_1 TAP_11314 (  );
sky130_fd_sc_hd__tap_1 TAP_11315 (  );
sky130_fd_sc_hd__tap_1 TAP_11316 (  );
sky130_fd_sc_hd__tap_1 TAP_11317 (  );
sky130_fd_sc_hd__tap_1 TAP_11318 (  );
sky130_fd_sc_hd__tap_1 TAP_11319 (  );
sky130_fd_sc_hd__tap_1 TAP_1132 (  );
sky130_fd_sc_hd__tap_1 TAP_11320 (  );
sky130_fd_sc_hd__tap_1 TAP_11321 (  );
sky130_fd_sc_hd__tap_1 TAP_11322 (  );
sky130_fd_sc_hd__tap_1 TAP_11323 (  );
sky130_fd_sc_hd__tap_1 TAP_11324 (  );
sky130_fd_sc_hd__tap_1 TAP_11325 (  );
sky130_fd_sc_hd__tap_1 TAP_11326 (  );
sky130_fd_sc_hd__tap_1 TAP_11327 (  );
sky130_fd_sc_hd__tap_1 TAP_11328 (  );
sky130_fd_sc_hd__tap_1 TAP_11329 (  );
sky130_fd_sc_hd__tap_1 TAP_1133 (  );
sky130_fd_sc_hd__tap_1 TAP_11330 (  );
sky130_fd_sc_hd__tap_1 TAP_11331 (  );
sky130_fd_sc_hd__tap_1 TAP_11332 (  );
sky130_fd_sc_hd__tap_1 TAP_11333 (  );
sky130_fd_sc_hd__tap_1 TAP_11334 (  );
sky130_fd_sc_hd__tap_1 TAP_11335 (  );
sky130_fd_sc_hd__tap_1 TAP_11336 (  );
sky130_fd_sc_hd__tap_1 TAP_11337 (  );
sky130_fd_sc_hd__tap_1 TAP_11338 (  );
sky130_fd_sc_hd__tap_1 TAP_11339 (  );
sky130_fd_sc_hd__tap_1 TAP_1134 (  );
sky130_fd_sc_hd__tap_1 TAP_11340 (  );
sky130_fd_sc_hd__tap_1 TAP_11341 (  );
sky130_fd_sc_hd__tap_1 TAP_11342 (  );
sky130_fd_sc_hd__tap_1 TAP_11343 (  );
sky130_fd_sc_hd__tap_1 TAP_11344 (  );
sky130_fd_sc_hd__tap_1 TAP_11345 (  );
sky130_fd_sc_hd__tap_1 TAP_11346 (  );
sky130_fd_sc_hd__tap_1 TAP_11347 (  );
sky130_fd_sc_hd__tap_1 TAP_11348 (  );
sky130_fd_sc_hd__tap_1 TAP_11349 (  );
sky130_fd_sc_hd__tap_1 TAP_1135 (  );
sky130_fd_sc_hd__tap_1 TAP_11350 (  );
sky130_fd_sc_hd__tap_1 TAP_11351 (  );
sky130_fd_sc_hd__tap_1 TAP_11352 (  );
sky130_fd_sc_hd__tap_1 TAP_11353 (  );
sky130_fd_sc_hd__tap_1 TAP_11354 (  );
sky130_fd_sc_hd__tap_1 TAP_11355 (  );
sky130_fd_sc_hd__tap_1 TAP_11356 (  );
sky130_fd_sc_hd__tap_1 TAP_11357 (  );
sky130_fd_sc_hd__tap_1 TAP_11358 (  );
sky130_fd_sc_hd__tap_1 TAP_11359 (  );
sky130_fd_sc_hd__tap_1 TAP_1136 (  );
sky130_fd_sc_hd__tap_1 TAP_11360 (  );
sky130_fd_sc_hd__tap_1 TAP_11361 (  );
sky130_fd_sc_hd__tap_1 TAP_11362 (  );
sky130_fd_sc_hd__tap_1 TAP_11363 (  );
sky130_fd_sc_hd__tap_1 TAP_11364 (  );
sky130_fd_sc_hd__tap_1 TAP_11365 (  );
sky130_fd_sc_hd__tap_1 TAP_11366 (  );
sky130_fd_sc_hd__tap_1 TAP_11367 (  );
sky130_fd_sc_hd__tap_1 TAP_11368 (  );
sky130_fd_sc_hd__tap_1 TAP_11369 (  );
sky130_fd_sc_hd__tap_1 TAP_1137 (  );
sky130_fd_sc_hd__tap_1 TAP_11370 (  );
sky130_fd_sc_hd__tap_1 TAP_11371 (  );
sky130_fd_sc_hd__tap_1 TAP_11372 (  );
sky130_fd_sc_hd__tap_1 TAP_11373 (  );
sky130_fd_sc_hd__tap_1 TAP_11374 (  );
sky130_fd_sc_hd__tap_1 TAP_11375 (  );
sky130_fd_sc_hd__tap_1 TAP_11376 (  );
sky130_fd_sc_hd__tap_1 TAP_11377 (  );
sky130_fd_sc_hd__tap_1 TAP_11378 (  );
sky130_fd_sc_hd__tap_1 TAP_11379 (  );
sky130_fd_sc_hd__tap_1 TAP_1138 (  );
sky130_fd_sc_hd__tap_1 TAP_11380 (  );
sky130_fd_sc_hd__tap_1 TAP_11381 (  );
sky130_fd_sc_hd__tap_1 TAP_11382 (  );
sky130_fd_sc_hd__tap_1 TAP_11383 (  );
sky130_fd_sc_hd__tap_1 TAP_11384 (  );
sky130_fd_sc_hd__tap_1 TAP_11385 (  );
sky130_fd_sc_hd__tap_1 TAP_11386 (  );
sky130_fd_sc_hd__tap_1 TAP_11387 (  );
sky130_fd_sc_hd__tap_1 TAP_11388 (  );
sky130_fd_sc_hd__tap_1 TAP_11389 (  );
sky130_fd_sc_hd__tap_1 TAP_1139 (  );
sky130_fd_sc_hd__tap_1 TAP_11390 (  );
sky130_fd_sc_hd__tap_1 TAP_11391 (  );
sky130_fd_sc_hd__tap_1 TAP_11392 (  );
sky130_fd_sc_hd__tap_1 TAP_11393 (  );
sky130_fd_sc_hd__tap_1 TAP_11394 (  );
sky130_fd_sc_hd__tap_1 TAP_11395 (  );
sky130_fd_sc_hd__tap_1 TAP_11396 (  );
sky130_fd_sc_hd__tap_1 TAP_11397 (  );
sky130_fd_sc_hd__tap_1 TAP_11398 (  );
sky130_fd_sc_hd__tap_1 TAP_11399 (  );
sky130_fd_sc_hd__tap_1 TAP_1140 (  );
sky130_fd_sc_hd__tap_1 TAP_11400 (  );
sky130_fd_sc_hd__tap_1 TAP_11401 (  );
sky130_fd_sc_hd__tap_1 TAP_11402 (  );
sky130_fd_sc_hd__tap_1 TAP_11403 (  );
sky130_fd_sc_hd__tap_1 TAP_11404 (  );
sky130_fd_sc_hd__tap_1 TAP_11405 (  );
sky130_fd_sc_hd__tap_1 TAP_11406 (  );
sky130_fd_sc_hd__tap_1 TAP_11407 (  );
sky130_fd_sc_hd__tap_1 TAP_11408 (  );
sky130_fd_sc_hd__tap_1 TAP_11409 (  );
sky130_fd_sc_hd__tap_1 TAP_1141 (  );
sky130_fd_sc_hd__tap_1 TAP_11410 (  );
sky130_fd_sc_hd__tap_1 TAP_11411 (  );
sky130_fd_sc_hd__tap_1 TAP_11412 (  );
sky130_fd_sc_hd__tap_1 TAP_11413 (  );
sky130_fd_sc_hd__tap_1 TAP_11414 (  );
sky130_fd_sc_hd__tap_1 TAP_11415 (  );
sky130_fd_sc_hd__tap_1 TAP_11416 (  );
sky130_fd_sc_hd__tap_1 TAP_11417 (  );
sky130_fd_sc_hd__tap_1 TAP_11418 (  );
sky130_fd_sc_hd__tap_1 TAP_11419 (  );
sky130_fd_sc_hd__tap_1 TAP_1142 (  );
sky130_fd_sc_hd__tap_1 TAP_11420 (  );
sky130_fd_sc_hd__tap_1 TAP_11421 (  );
sky130_fd_sc_hd__tap_1 TAP_11422 (  );
sky130_fd_sc_hd__tap_1 TAP_11423 (  );
sky130_fd_sc_hd__tap_1 TAP_11424 (  );
sky130_fd_sc_hd__tap_1 TAP_11425 (  );
sky130_fd_sc_hd__tap_1 TAP_11426 (  );
sky130_fd_sc_hd__tap_1 TAP_11427 (  );
sky130_fd_sc_hd__tap_1 TAP_11428 (  );
sky130_fd_sc_hd__tap_1 TAP_11429 (  );
sky130_fd_sc_hd__tap_1 TAP_1143 (  );
sky130_fd_sc_hd__tap_1 TAP_11430 (  );
sky130_fd_sc_hd__tap_1 TAP_11431 (  );
sky130_fd_sc_hd__tap_1 TAP_11432 (  );
sky130_fd_sc_hd__tap_1 TAP_11433 (  );
sky130_fd_sc_hd__tap_1 TAP_11434 (  );
sky130_fd_sc_hd__tap_1 TAP_11435 (  );
sky130_fd_sc_hd__tap_1 TAP_11436 (  );
sky130_fd_sc_hd__tap_1 TAP_11437 (  );
sky130_fd_sc_hd__tap_1 TAP_11438 (  );
sky130_fd_sc_hd__tap_1 TAP_11439 (  );
sky130_fd_sc_hd__tap_1 TAP_1144 (  );
sky130_fd_sc_hd__tap_1 TAP_11440 (  );
sky130_fd_sc_hd__tap_1 TAP_11441 (  );
sky130_fd_sc_hd__tap_1 TAP_11442 (  );
sky130_fd_sc_hd__tap_1 TAP_11443 (  );
sky130_fd_sc_hd__tap_1 TAP_11444 (  );
sky130_fd_sc_hd__tap_1 TAP_11445 (  );
sky130_fd_sc_hd__tap_1 TAP_11446 (  );
sky130_fd_sc_hd__tap_1 TAP_11447 (  );
sky130_fd_sc_hd__tap_1 TAP_11448 (  );
sky130_fd_sc_hd__tap_1 TAP_11449 (  );
sky130_fd_sc_hd__tap_1 TAP_1145 (  );
sky130_fd_sc_hd__tap_1 TAP_11450 (  );
sky130_fd_sc_hd__tap_1 TAP_11451 (  );
sky130_fd_sc_hd__tap_1 TAP_11452 (  );
sky130_fd_sc_hd__tap_1 TAP_11453 (  );
sky130_fd_sc_hd__tap_1 TAP_11454 (  );
sky130_fd_sc_hd__tap_1 TAP_11455 (  );
sky130_fd_sc_hd__tap_1 TAP_11456 (  );
sky130_fd_sc_hd__tap_1 TAP_11457 (  );
sky130_fd_sc_hd__tap_1 TAP_11458 (  );
sky130_fd_sc_hd__tap_1 TAP_11459 (  );
sky130_fd_sc_hd__tap_1 TAP_1146 (  );
sky130_fd_sc_hd__tap_1 TAP_11460 (  );
sky130_fd_sc_hd__tap_1 TAP_11461 (  );
sky130_fd_sc_hd__tap_1 TAP_11462 (  );
sky130_fd_sc_hd__tap_1 TAP_11463 (  );
sky130_fd_sc_hd__tap_1 TAP_11464 (  );
sky130_fd_sc_hd__tap_1 TAP_11465 (  );
sky130_fd_sc_hd__tap_1 TAP_11466 (  );
sky130_fd_sc_hd__tap_1 TAP_11467 (  );
sky130_fd_sc_hd__tap_1 TAP_11468 (  );
sky130_fd_sc_hd__tap_1 TAP_11469 (  );
sky130_fd_sc_hd__tap_1 TAP_1147 (  );
sky130_fd_sc_hd__tap_1 TAP_11470 (  );
sky130_fd_sc_hd__tap_1 TAP_11471 (  );
sky130_fd_sc_hd__tap_1 TAP_11472 (  );
sky130_fd_sc_hd__tap_1 TAP_11473 (  );
sky130_fd_sc_hd__tap_1 TAP_11474 (  );
sky130_fd_sc_hd__tap_1 TAP_11475 (  );
sky130_fd_sc_hd__tap_1 TAP_11476 (  );
sky130_fd_sc_hd__tap_1 TAP_11477 (  );
sky130_fd_sc_hd__tap_1 TAP_11478 (  );
sky130_fd_sc_hd__tap_1 TAP_11479 (  );
sky130_fd_sc_hd__tap_1 TAP_1148 (  );
sky130_fd_sc_hd__tap_1 TAP_11480 (  );
sky130_fd_sc_hd__tap_1 TAP_11481 (  );
sky130_fd_sc_hd__tap_1 TAP_11482 (  );
sky130_fd_sc_hd__tap_1 TAP_11483 (  );
sky130_fd_sc_hd__tap_1 TAP_11484 (  );
sky130_fd_sc_hd__tap_1 TAP_11485 (  );
sky130_fd_sc_hd__tap_1 TAP_11486 (  );
sky130_fd_sc_hd__tap_1 TAP_11487 (  );
sky130_fd_sc_hd__tap_1 TAP_11488 (  );
sky130_fd_sc_hd__tap_1 TAP_11489 (  );
sky130_fd_sc_hd__tap_1 TAP_1149 (  );
sky130_fd_sc_hd__tap_1 TAP_11490 (  );
sky130_fd_sc_hd__tap_1 TAP_11491 (  );
sky130_fd_sc_hd__tap_1 TAP_11492 (  );
sky130_fd_sc_hd__tap_1 TAP_11493 (  );
sky130_fd_sc_hd__tap_1 TAP_11494 (  );
sky130_fd_sc_hd__tap_1 TAP_11495 (  );
sky130_fd_sc_hd__tap_1 TAP_11496 (  );
sky130_fd_sc_hd__tap_1 TAP_11497 (  );
sky130_fd_sc_hd__tap_1 TAP_11498 (  );
sky130_fd_sc_hd__tap_1 TAP_11499 (  );
sky130_fd_sc_hd__tap_1 TAP_1150 (  );
sky130_fd_sc_hd__tap_1 TAP_11500 (  );
sky130_fd_sc_hd__tap_1 TAP_11501 (  );
sky130_fd_sc_hd__tap_1 TAP_11502 (  );
sky130_fd_sc_hd__tap_1 TAP_11503 (  );
sky130_fd_sc_hd__tap_1 TAP_11504 (  );
sky130_fd_sc_hd__tap_1 TAP_11505 (  );
sky130_fd_sc_hd__tap_1 TAP_11506 (  );
sky130_fd_sc_hd__tap_1 TAP_11507 (  );
sky130_fd_sc_hd__tap_1 TAP_11508 (  );
sky130_fd_sc_hd__tap_1 TAP_11509 (  );
sky130_fd_sc_hd__tap_1 TAP_1151 (  );
sky130_fd_sc_hd__tap_1 TAP_11510 (  );
sky130_fd_sc_hd__tap_1 TAP_11511 (  );
sky130_fd_sc_hd__tap_1 TAP_11512 (  );
sky130_fd_sc_hd__tap_1 TAP_11513 (  );
sky130_fd_sc_hd__tap_1 TAP_11514 (  );
sky130_fd_sc_hd__tap_1 TAP_11515 (  );
sky130_fd_sc_hd__tap_1 TAP_11516 (  );
sky130_fd_sc_hd__tap_1 TAP_11517 (  );
sky130_fd_sc_hd__tap_1 TAP_11518 (  );
sky130_fd_sc_hd__tap_1 TAP_11519 (  );
sky130_fd_sc_hd__tap_1 TAP_1152 (  );
sky130_fd_sc_hd__tap_1 TAP_11520 (  );
sky130_fd_sc_hd__tap_1 TAP_11521 (  );
sky130_fd_sc_hd__tap_1 TAP_11522 (  );
sky130_fd_sc_hd__tap_1 TAP_11523 (  );
sky130_fd_sc_hd__tap_1 TAP_11524 (  );
sky130_fd_sc_hd__tap_1 TAP_11525 (  );
sky130_fd_sc_hd__tap_1 TAP_11526 (  );
sky130_fd_sc_hd__tap_1 TAP_11527 (  );
sky130_fd_sc_hd__tap_1 TAP_11528 (  );
sky130_fd_sc_hd__tap_1 TAP_11529 (  );
sky130_fd_sc_hd__tap_1 TAP_1153 (  );
sky130_fd_sc_hd__tap_1 TAP_11530 (  );
sky130_fd_sc_hd__tap_1 TAP_11531 (  );
sky130_fd_sc_hd__tap_1 TAP_11532 (  );
sky130_fd_sc_hd__tap_1 TAP_11533 (  );
sky130_fd_sc_hd__tap_1 TAP_11534 (  );
sky130_fd_sc_hd__tap_1 TAP_11535 (  );
sky130_fd_sc_hd__tap_1 TAP_11536 (  );
sky130_fd_sc_hd__tap_1 TAP_11537 (  );
sky130_fd_sc_hd__tap_1 TAP_11538 (  );
sky130_fd_sc_hd__tap_1 TAP_11539 (  );
sky130_fd_sc_hd__tap_1 TAP_1154 (  );
sky130_fd_sc_hd__tap_1 TAP_11540 (  );
sky130_fd_sc_hd__tap_1 TAP_11541 (  );
sky130_fd_sc_hd__tap_1 TAP_11542 (  );
sky130_fd_sc_hd__tap_1 TAP_11543 (  );
sky130_fd_sc_hd__tap_1 TAP_11544 (  );
sky130_fd_sc_hd__tap_1 TAP_11545 (  );
sky130_fd_sc_hd__tap_1 TAP_11546 (  );
sky130_fd_sc_hd__tap_1 TAP_11547 (  );
sky130_fd_sc_hd__tap_1 TAP_11548 (  );
sky130_fd_sc_hd__tap_1 TAP_11549 (  );
sky130_fd_sc_hd__tap_1 TAP_1155 (  );
sky130_fd_sc_hd__tap_1 TAP_11550 (  );
sky130_fd_sc_hd__tap_1 TAP_11551 (  );
sky130_fd_sc_hd__tap_1 TAP_11552 (  );
sky130_fd_sc_hd__tap_1 TAP_11553 (  );
sky130_fd_sc_hd__tap_1 TAP_11554 (  );
sky130_fd_sc_hd__tap_1 TAP_11555 (  );
sky130_fd_sc_hd__tap_1 TAP_11556 (  );
sky130_fd_sc_hd__tap_1 TAP_11557 (  );
sky130_fd_sc_hd__tap_1 TAP_11558 (  );
sky130_fd_sc_hd__tap_1 TAP_11559 (  );
sky130_fd_sc_hd__tap_1 TAP_1156 (  );
sky130_fd_sc_hd__tap_1 TAP_11560 (  );
sky130_fd_sc_hd__tap_1 TAP_11561 (  );
sky130_fd_sc_hd__tap_1 TAP_11562 (  );
sky130_fd_sc_hd__tap_1 TAP_11563 (  );
sky130_fd_sc_hd__tap_1 TAP_11564 (  );
sky130_fd_sc_hd__tap_1 TAP_11565 (  );
sky130_fd_sc_hd__tap_1 TAP_11566 (  );
sky130_fd_sc_hd__tap_1 TAP_11567 (  );
sky130_fd_sc_hd__tap_1 TAP_11568 (  );
sky130_fd_sc_hd__tap_1 TAP_11569 (  );
sky130_fd_sc_hd__tap_1 TAP_1157 (  );
sky130_fd_sc_hd__tap_1 TAP_11570 (  );
sky130_fd_sc_hd__tap_1 TAP_11571 (  );
sky130_fd_sc_hd__tap_1 TAP_11572 (  );
sky130_fd_sc_hd__tap_1 TAP_11573 (  );
sky130_fd_sc_hd__tap_1 TAP_11574 (  );
sky130_fd_sc_hd__tap_1 TAP_11575 (  );
sky130_fd_sc_hd__tap_1 TAP_11576 (  );
sky130_fd_sc_hd__tap_1 TAP_11577 (  );
sky130_fd_sc_hd__tap_1 TAP_11578 (  );
sky130_fd_sc_hd__tap_1 TAP_11579 (  );
sky130_fd_sc_hd__tap_1 TAP_1158 (  );
sky130_fd_sc_hd__tap_1 TAP_11580 (  );
sky130_fd_sc_hd__tap_1 TAP_11581 (  );
sky130_fd_sc_hd__tap_1 TAP_11582 (  );
sky130_fd_sc_hd__tap_1 TAP_11583 (  );
sky130_fd_sc_hd__tap_1 TAP_11584 (  );
sky130_fd_sc_hd__tap_1 TAP_11585 (  );
sky130_fd_sc_hd__tap_1 TAP_11586 (  );
sky130_fd_sc_hd__tap_1 TAP_11587 (  );
sky130_fd_sc_hd__tap_1 TAP_11588 (  );
sky130_fd_sc_hd__tap_1 TAP_11589 (  );
sky130_fd_sc_hd__tap_1 TAP_1159 (  );
sky130_fd_sc_hd__tap_1 TAP_11590 (  );
sky130_fd_sc_hd__tap_1 TAP_11591 (  );
sky130_fd_sc_hd__tap_1 TAP_11592 (  );
sky130_fd_sc_hd__tap_1 TAP_11593 (  );
sky130_fd_sc_hd__tap_1 TAP_11594 (  );
sky130_fd_sc_hd__tap_1 TAP_11595 (  );
sky130_fd_sc_hd__tap_1 TAP_11596 (  );
sky130_fd_sc_hd__tap_1 TAP_11597 (  );
sky130_fd_sc_hd__tap_1 TAP_11598 (  );
sky130_fd_sc_hd__tap_1 TAP_11599 (  );
sky130_fd_sc_hd__tap_1 TAP_1160 (  );
sky130_fd_sc_hd__tap_1 TAP_11600 (  );
sky130_fd_sc_hd__tap_1 TAP_11601 (  );
sky130_fd_sc_hd__tap_1 TAP_11602 (  );
sky130_fd_sc_hd__tap_1 TAP_11603 (  );
sky130_fd_sc_hd__tap_1 TAP_11604 (  );
sky130_fd_sc_hd__tap_1 TAP_11605 (  );
sky130_fd_sc_hd__tap_1 TAP_11606 (  );
sky130_fd_sc_hd__tap_1 TAP_11607 (  );
sky130_fd_sc_hd__tap_1 TAP_11608 (  );
sky130_fd_sc_hd__tap_1 TAP_11609 (  );
sky130_fd_sc_hd__tap_1 TAP_1161 (  );
sky130_fd_sc_hd__tap_1 TAP_11610 (  );
sky130_fd_sc_hd__tap_1 TAP_11611 (  );
sky130_fd_sc_hd__tap_1 TAP_11612 (  );
sky130_fd_sc_hd__tap_1 TAP_11613 (  );
sky130_fd_sc_hd__tap_1 TAP_11614 (  );
sky130_fd_sc_hd__tap_1 TAP_11615 (  );
sky130_fd_sc_hd__tap_1 TAP_11616 (  );
sky130_fd_sc_hd__tap_1 TAP_11617 (  );
sky130_fd_sc_hd__tap_1 TAP_11618 (  );
sky130_fd_sc_hd__tap_1 TAP_11619 (  );
sky130_fd_sc_hd__tap_1 TAP_1162 (  );
sky130_fd_sc_hd__tap_1 TAP_11620 (  );
sky130_fd_sc_hd__tap_1 TAP_11621 (  );
sky130_fd_sc_hd__tap_1 TAP_11622 (  );
sky130_fd_sc_hd__tap_1 TAP_11623 (  );
sky130_fd_sc_hd__tap_1 TAP_11624 (  );
sky130_fd_sc_hd__tap_1 TAP_11625 (  );
sky130_fd_sc_hd__tap_1 TAP_11626 (  );
sky130_fd_sc_hd__tap_1 TAP_11627 (  );
sky130_fd_sc_hd__tap_1 TAP_11628 (  );
sky130_fd_sc_hd__tap_1 TAP_11629 (  );
sky130_fd_sc_hd__tap_1 TAP_1163 (  );
sky130_fd_sc_hd__tap_1 TAP_11630 (  );
sky130_fd_sc_hd__tap_1 TAP_11631 (  );
sky130_fd_sc_hd__tap_1 TAP_11632 (  );
sky130_fd_sc_hd__tap_1 TAP_11633 (  );
sky130_fd_sc_hd__tap_1 TAP_11634 (  );
sky130_fd_sc_hd__tap_1 TAP_11635 (  );
sky130_fd_sc_hd__tap_1 TAP_11636 (  );
sky130_fd_sc_hd__tap_1 TAP_11637 (  );
sky130_fd_sc_hd__tap_1 TAP_11638 (  );
sky130_fd_sc_hd__tap_1 TAP_11639 (  );
sky130_fd_sc_hd__tap_1 TAP_1164 (  );
sky130_fd_sc_hd__tap_1 TAP_11640 (  );
sky130_fd_sc_hd__tap_1 TAP_11641 (  );
sky130_fd_sc_hd__tap_1 TAP_11642 (  );
sky130_fd_sc_hd__tap_1 TAP_11643 (  );
sky130_fd_sc_hd__tap_1 TAP_11644 (  );
sky130_fd_sc_hd__tap_1 TAP_11645 (  );
sky130_fd_sc_hd__tap_1 TAP_11646 (  );
sky130_fd_sc_hd__tap_1 TAP_11647 (  );
sky130_fd_sc_hd__tap_1 TAP_11648 (  );
sky130_fd_sc_hd__tap_1 TAP_11649 (  );
sky130_fd_sc_hd__tap_1 TAP_1165 (  );
sky130_fd_sc_hd__tap_1 TAP_11650 (  );
sky130_fd_sc_hd__tap_1 TAP_11651 (  );
sky130_fd_sc_hd__tap_1 TAP_11652 (  );
sky130_fd_sc_hd__tap_1 TAP_11653 (  );
sky130_fd_sc_hd__tap_1 TAP_11654 (  );
sky130_fd_sc_hd__tap_1 TAP_11655 (  );
sky130_fd_sc_hd__tap_1 TAP_11656 (  );
sky130_fd_sc_hd__tap_1 TAP_11657 (  );
sky130_fd_sc_hd__tap_1 TAP_11658 (  );
sky130_fd_sc_hd__tap_1 TAP_11659 (  );
sky130_fd_sc_hd__tap_1 TAP_1166 (  );
sky130_fd_sc_hd__tap_1 TAP_11660 (  );
sky130_fd_sc_hd__tap_1 TAP_11661 (  );
sky130_fd_sc_hd__tap_1 TAP_11662 (  );
sky130_fd_sc_hd__tap_1 TAP_11663 (  );
sky130_fd_sc_hd__tap_1 TAP_11664 (  );
sky130_fd_sc_hd__tap_1 TAP_11665 (  );
sky130_fd_sc_hd__tap_1 TAP_11666 (  );
sky130_fd_sc_hd__tap_1 TAP_11667 (  );
sky130_fd_sc_hd__tap_1 TAP_11668 (  );
sky130_fd_sc_hd__tap_1 TAP_11669 (  );
sky130_fd_sc_hd__tap_1 TAP_1167 (  );
sky130_fd_sc_hd__tap_1 TAP_11670 (  );
sky130_fd_sc_hd__tap_1 TAP_11671 (  );
sky130_fd_sc_hd__tap_1 TAP_11672 (  );
sky130_fd_sc_hd__tap_1 TAP_11673 (  );
sky130_fd_sc_hd__tap_1 TAP_11674 (  );
sky130_fd_sc_hd__tap_1 TAP_11675 (  );
sky130_fd_sc_hd__tap_1 TAP_11676 (  );
sky130_fd_sc_hd__tap_1 TAP_11677 (  );
sky130_fd_sc_hd__tap_1 TAP_11678 (  );
sky130_fd_sc_hd__tap_1 TAP_11679 (  );
sky130_fd_sc_hd__tap_1 TAP_1168 (  );
sky130_fd_sc_hd__tap_1 TAP_11680 (  );
sky130_fd_sc_hd__tap_1 TAP_11681 (  );
sky130_fd_sc_hd__tap_1 TAP_11682 (  );
sky130_fd_sc_hd__tap_1 TAP_11683 (  );
sky130_fd_sc_hd__tap_1 TAP_11684 (  );
sky130_fd_sc_hd__tap_1 TAP_11685 (  );
sky130_fd_sc_hd__tap_1 TAP_11686 (  );
sky130_fd_sc_hd__tap_1 TAP_11687 (  );
sky130_fd_sc_hd__tap_1 TAP_11688 (  );
sky130_fd_sc_hd__tap_1 TAP_11689 (  );
sky130_fd_sc_hd__tap_1 TAP_1169 (  );
sky130_fd_sc_hd__tap_1 TAP_11690 (  );
sky130_fd_sc_hd__tap_1 TAP_11691 (  );
sky130_fd_sc_hd__tap_1 TAP_11692 (  );
sky130_fd_sc_hd__tap_1 TAP_11693 (  );
sky130_fd_sc_hd__tap_1 TAP_11694 (  );
sky130_fd_sc_hd__tap_1 TAP_11695 (  );
sky130_fd_sc_hd__tap_1 TAP_11696 (  );
sky130_fd_sc_hd__tap_1 TAP_11697 (  );
sky130_fd_sc_hd__tap_1 TAP_11698 (  );
sky130_fd_sc_hd__tap_1 TAP_11699 (  );
sky130_fd_sc_hd__tap_1 TAP_1170 (  );
sky130_fd_sc_hd__tap_1 TAP_11700 (  );
sky130_fd_sc_hd__tap_1 TAP_11701 (  );
sky130_fd_sc_hd__tap_1 TAP_11702 (  );
sky130_fd_sc_hd__tap_1 TAP_11703 (  );
sky130_fd_sc_hd__tap_1 TAP_11704 (  );
sky130_fd_sc_hd__tap_1 TAP_11705 (  );
sky130_fd_sc_hd__tap_1 TAP_11706 (  );
sky130_fd_sc_hd__tap_1 TAP_11707 (  );
sky130_fd_sc_hd__tap_1 TAP_11708 (  );
sky130_fd_sc_hd__tap_1 TAP_11709 (  );
sky130_fd_sc_hd__tap_1 TAP_1171 (  );
sky130_fd_sc_hd__tap_1 TAP_11710 (  );
sky130_fd_sc_hd__tap_1 TAP_11711 (  );
sky130_fd_sc_hd__tap_1 TAP_11712 (  );
sky130_fd_sc_hd__tap_1 TAP_11713 (  );
sky130_fd_sc_hd__tap_1 TAP_11714 (  );
sky130_fd_sc_hd__tap_1 TAP_11715 (  );
sky130_fd_sc_hd__tap_1 TAP_11716 (  );
sky130_fd_sc_hd__tap_1 TAP_11717 (  );
sky130_fd_sc_hd__tap_1 TAP_11718 (  );
sky130_fd_sc_hd__tap_1 TAP_11719 (  );
sky130_fd_sc_hd__tap_1 TAP_1172 (  );
sky130_fd_sc_hd__tap_1 TAP_11720 (  );
sky130_fd_sc_hd__tap_1 TAP_11721 (  );
sky130_fd_sc_hd__tap_1 TAP_11722 (  );
sky130_fd_sc_hd__tap_1 TAP_11723 (  );
sky130_fd_sc_hd__tap_1 TAP_11724 (  );
sky130_fd_sc_hd__tap_1 TAP_11725 (  );
sky130_fd_sc_hd__tap_1 TAP_11726 (  );
sky130_fd_sc_hd__tap_1 TAP_11727 (  );
sky130_fd_sc_hd__tap_1 TAP_11728 (  );
sky130_fd_sc_hd__tap_1 TAP_11729 (  );
sky130_fd_sc_hd__tap_1 TAP_1173 (  );
sky130_fd_sc_hd__tap_1 TAP_11730 (  );
sky130_fd_sc_hd__tap_1 TAP_11731 (  );
sky130_fd_sc_hd__tap_1 TAP_11732 (  );
sky130_fd_sc_hd__tap_1 TAP_11733 (  );
sky130_fd_sc_hd__tap_1 TAP_11734 (  );
sky130_fd_sc_hd__tap_1 TAP_11735 (  );
sky130_fd_sc_hd__tap_1 TAP_11736 (  );
sky130_fd_sc_hd__tap_1 TAP_11737 (  );
sky130_fd_sc_hd__tap_1 TAP_11738 (  );
sky130_fd_sc_hd__tap_1 TAP_11739 (  );
sky130_fd_sc_hd__tap_1 TAP_1174 (  );
sky130_fd_sc_hd__tap_1 TAP_11740 (  );
sky130_fd_sc_hd__tap_1 TAP_11741 (  );
sky130_fd_sc_hd__tap_1 TAP_11742 (  );
sky130_fd_sc_hd__tap_1 TAP_11743 (  );
sky130_fd_sc_hd__tap_1 TAP_11744 (  );
sky130_fd_sc_hd__tap_1 TAP_11745 (  );
sky130_fd_sc_hd__tap_1 TAP_11746 (  );
sky130_fd_sc_hd__tap_1 TAP_11747 (  );
sky130_fd_sc_hd__tap_1 TAP_11748 (  );
sky130_fd_sc_hd__tap_1 TAP_11749 (  );
sky130_fd_sc_hd__tap_1 TAP_1175 (  );
sky130_fd_sc_hd__tap_1 TAP_11750 (  );
sky130_fd_sc_hd__tap_1 TAP_11751 (  );
sky130_fd_sc_hd__tap_1 TAP_11752 (  );
sky130_fd_sc_hd__tap_1 TAP_11753 (  );
sky130_fd_sc_hd__tap_1 TAP_11754 (  );
sky130_fd_sc_hd__tap_1 TAP_11755 (  );
sky130_fd_sc_hd__tap_1 TAP_11756 (  );
sky130_fd_sc_hd__tap_1 TAP_11757 (  );
sky130_fd_sc_hd__tap_1 TAP_11758 (  );
sky130_fd_sc_hd__tap_1 TAP_11759 (  );
sky130_fd_sc_hd__tap_1 TAP_1176 (  );
sky130_fd_sc_hd__tap_1 TAP_11760 (  );
sky130_fd_sc_hd__tap_1 TAP_11761 (  );
sky130_fd_sc_hd__tap_1 TAP_11762 (  );
sky130_fd_sc_hd__tap_1 TAP_11763 (  );
sky130_fd_sc_hd__tap_1 TAP_11764 (  );
sky130_fd_sc_hd__tap_1 TAP_11765 (  );
sky130_fd_sc_hd__tap_1 TAP_11766 (  );
sky130_fd_sc_hd__tap_1 TAP_11767 (  );
sky130_fd_sc_hd__tap_1 TAP_11768 (  );
sky130_fd_sc_hd__tap_1 TAP_11769 (  );
sky130_fd_sc_hd__tap_1 TAP_1177 (  );
sky130_fd_sc_hd__tap_1 TAP_11770 (  );
sky130_fd_sc_hd__tap_1 TAP_11771 (  );
sky130_fd_sc_hd__tap_1 TAP_11772 (  );
sky130_fd_sc_hd__tap_1 TAP_11773 (  );
sky130_fd_sc_hd__tap_1 TAP_11774 (  );
sky130_fd_sc_hd__tap_1 TAP_11775 (  );
sky130_fd_sc_hd__tap_1 TAP_11776 (  );
sky130_fd_sc_hd__tap_1 TAP_11777 (  );
sky130_fd_sc_hd__tap_1 TAP_11778 (  );
sky130_fd_sc_hd__tap_1 TAP_11779 (  );
sky130_fd_sc_hd__tap_1 TAP_1178 (  );
sky130_fd_sc_hd__tap_1 TAP_11780 (  );
sky130_fd_sc_hd__tap_1 TAP_11781 (  );
sky130_fd_sc_hd__tap_1 TAP_11782 (  );
sky130_fd_sc_hd__tap_1 TAP_11783 (  );
sky130_fd_sc_hd__tap_1 TAP_11784 (  );
sky130_fd_sc_hd__tap_1 TAP_11785 (  );
sky130_fd_sc_hd__tap_1 TAP_11786 (  );
sky130_fd_sc_hd__tap_1 TAP_11787 (  );
sky130_fd_sc_hd__tap_1 TAP_11788 (  );
sky130_fd_sc_hd__tap_1 TAP_11789 (  );
sky130_fd_sc_hd__tap_1 TAP_1179 (  );
sky130_fd_sc_hd__tap_1 TAP_11790 (  );
sky130_fd_sc_hd__tap_1 TAP_11791 (  );
sky130_fd_sc_hd__tap_1 TAP_11792 (  );
sky130_fd_sc_hd__tap_1 TAP_11793 (  );
sky130_fd_sc_hd__tap_1 TAP_11794 (  );
sky130_fd_sc_hd__tap_1 TAP_11795 (  );
sky130_fd_sc_hd__tap_1 TAP_11796 (  );
sky130_fd_sc_hd__tap_1 TAP_11797 (  );
sky130_fd_sc_hd__tap_1 TAP_11798 (  );
sky130_fd_sc_hd__tap_1 TAP_11799 (  );
sky130_fd_sc_hd__tap_1 TAP_1180 (  );
sky130_fd_sc_hd__tap_1 TAP_11800 (  );
sky130_fd_sc_hd__tap_1 TAP_11801 (  );
sky130_fd_sc_hd__tap_1 TAP_11802 (  );
sky130_fd_sc_hd__tap_1 TAP_11803 (  );
sky130_fd_sc_hd__tap_1 TAP_11804 (  );
sky130_fd_sc_hd__tap_1 TAP_11805 (  );
sky130_fd_sc_hd__tap_1 TAP_11806 (  );
sky130_fd_sc_hd__tap_1 TAP_11807 (  );
sky130_fd_sc_hd__tap_1 TAP_11808 (  );
sky130_fd_sc_hd__tap_1 TAP_11809 (  );
sky130_fd_sc_hd__tap_1 TAP_1181 (  );
sky130_fd_sc_hd__tap_1 TAP_11810 (  );
sky130_fd_sc_hd__tap_1 TAP_11811 (  );
sky130_fd_sc_hd__tap_1 TAP_11812 (  );
sky130_fd_sc_hd__tap_1 TAP_11813 (  );
sky130_fd_sc_hd__tap_1 TAP_11814 (  );
sky130_fd_sc_hd__tap_1 TAP_11815 (  );
sky130_fd_sc_hd__tap_1 TAP_11816 (  );
sky130_fd_sc_hd__tap_1 TAP_11817 (  );
sky130_fd_sc_hd__tap_1 TAP_11818 (  );
sky130_fd_sc_hd__tap_1 TAP_11819 (  );
sky130_fd_sc_hd__tap_1 TAP_1182 (  );
sky130_fd_sc_hd__tap_1 TAP_11820 (  );
sky130_fd_sc_hd__tap_1 TAP_11821 (  );
sky130_fd_sc_hd__tap_1 TAP_11822 (  );
sky130_fd_sc_hd__tap_1 TAP_11823 (  );
sky130_fd_sc_hd__tap_1 TAP_11824 (  );
sky130_fd_sc_hd__tap_1 TAP_11825 (  );
sky130_fd_sc_hd__tap_1 TAP_11826 (  );
sky130_fd_sc_hd__tap_1 TAP_11827 (  );
sky130_fd_sc_hd__tap_1 TAP_11828 (  );
sky130_fd_sc_hd__tap_1 TAP_11829 (  );
sky130_fd_sc_hd__tap_1 TAP_1183 (  );
sky130_fd_sc_hd__tap_1 TAP_11830 (  );
sky130_fd_sc_hd__tap_1 TAP_11831 (  );
sky130_fd_sc_hd__tap_1 TAP_11832 (  );
sky130_fd_sc_hd__tap_1 TAP_11833 (  );
sky130_fd_sc_hd__tap_1 TAP_11834 (  );
sky130_fd_sc_hd__tap_1 TAP_11835 (  );
sky130_fd_sc_hd__tap_1 TAP_11836 (  );
sky130_fd_sc_hd__tap_1 TAP_11837 (  );
sky130_fd_sc_hd__tap_1 TAP_11838 (  );
sky130_fd_sc_hd__tap_1 TAP_11839 (  );
sky130_fd_sc_hd__tap_1 TAP_1184 (  );
sky130_fd_sc_hd__tap_1 TAP_11840 (  );
sky130_fd_sc_hd__tap_1 TAP_11841 (  );
sky130_fd_sc_hd__tap_1 TAP_11842 (  );
sky130_fd_sc_hd__tap_1 TAP_11843 (  );
sky130_fd_sc_hd__tap_1 TAP_11844 (  );
sky130_fd_sc_hd__tap_1 TAP_11845 (  );
sky130_fd_sc_hd__tap_1 TAP_11846 (  );
sky130_fd_sc_hd__tap_1 TAP_11847 (  );
sky130_fd_sc_hd__tap_1 TAP_11848 (  );
sky130_fd_sc_hd__tap_1 TAP_11849 (  );
sky130_fd_sc_hd__tap_1 TAP_1185 (  );
sky130_fd_sc_hd__tap_1 TAP_11850 (  );
sky130_fd_sc_hd__tap_1 TAP_11851 (  );
sky130_fd_sc_hd__tap_1 TAP_11852 (  );
sky130_fd_sc_hd__tap_1 TAP_11853 (  );
sky130_fd_sc_hd__tap_1 TAP_11854 (  );
sky130_fd_sc_hd__tap_1 TAP_11855 (  );
sky130_fd_sc_hd__tap_1 TAP_11856 (  );
sky130_fd_sc_hd__tap_1 TAP_11857 (  );
sky130_fd_sc_hd__tap_1 TAP_11858 (  );
sky130_fd_sc_hd__tap_1 TAP_11859 (  );
sky130_fd_sc_hd__tap_1 TAP_1186 (  );
sky130_fd_sc_hd__tap_1 TAP_11860 (  );
sky130_fd_sc_hd__tap_1 TAP_11861 (  );
sky130_fd_sc_hd__tap_1 TAP_11862 (  );
sky130_fd_sc_hd__tap_1 TAP_11863 (  );
sky130_fd_sc_hd__tap_1 TAP_11864 (  );
sky130_fd_sc_hd__tap_1 TAP_11865 (  );
sky130_fd_sc_hd__tap_1 TAP_11866 (  );
sky130_fd_sc_hd__tap_1 TAP_11867 (  );
sky130_fd_sc_hd__tap_1 TAP_11868 (  );
sky130_fd_sc_hd__tap_1 TAP_11869 (  );
sky130_fd_sc_hd__tap_1 TAP_1187 (  );
sky130_fd_sc_hd__tap_1 TAP_11870 (  );
sky130_fd_sc_hd__tap_1 TAP_11871 (  );
sky130_fd_sc_hd__tap_1 TAP_11872 (  );
sky130_fd_sc_hd__tap_1 TAP_11873 (  );
sky130_fd_sc_hd__tap_1 TAP_11874 (  );
sky130_fd_sc_hd__tap_1 TAP_11875 (  );
sky130_fd_sc_hd__tap_1 TAP_11876 (  );
sky130_fd_sc_hd__tap_1 TAP_11877 (  );
sky130_fd_sc_hd__tap_1 TAP_11878 (  );
sky130_fd_sc_hd__tap_1 TAP_11879 (  );
sky130_fd_sc_hd__tap_1 TAP_1188 (  );
sky130_fd_sc_hd__tap_1 TAP_11880 (  );
sky130_fd_sc_hd__tap_1 TAP_11881 (  );
sky130_fd_sc_hd__tap_1 TAP_11882 (  );
sky130_fd_sc_hd__tap_1 TAP_11883 (  );
sky130_fd_sc_hd__tap_1 TAP_11884 (  );
sky130_fd_sc_hd__tap_1 TAP_11885 (  );
sky130_fd_sc_hd__tap_1 TAP_11886 (  );
sky130_fd_sc_hd__tap_1 TAP_11887 (  );
sky130_fd_sc_hd__tap_1 TAP_11888 (  );
sky130_fd_sc_hd__tap_1 TAP_11889 (  );
sky130_fd_sc_hd__tap_1 TAP_1189 (  );
sky130_fd_sc_hd__tap_1 TAP_11890 (  );
sky130_fd_sc_hd__tap_1 TAP_11891 (  );
sky130_fd_sc_hd__tap_1 TAP_11892 (  );
sky130_fd_sc_hd__tap_1 TAP_11893 (  );
sky130_fd_sc_hd__tap_1 TAP_11894 (  );
sky130_fd_sc_hd__tap_1 TAP_11895 (  );
sky130_fd_sc_hd__tap_1 TAP_11896 (  );
sky130_fd_sc_hd__tap_1 TAP_11897 (  );
sky130_fd_sc_hd__tap_1 TAP_11898 (  );
sky130_fd_sc_hd__tap_1 TAP_11899 (  );
sky130_fd_sc_hd__tap_1 TAP_1190 (  );
sky130_fd_sc_hd__tap_1 TAP_11900 (  );
sky130_fd_sc_hd__tap_1 TAP_11901 (  );
sky130_fd_sc_hd__tap_1 TAP_11902 (  );
sky130_fd_sc_hd__tap_1 TAP_11903 (  );
sky130_fd_sc_hd__tap_1 TAP_11904 (  );
sky130_fd_sc_hd__tap_1 TAP_11905 (  );
sky130_fd_sc_hd__tap_1 TAP_11906 (  );
sky130_fd_sc_hd__tap_1 TAP_11907 (  );
sky130_fd_sc_hd__tap_1 TAP_11908 (  );
sky130_fd_sc_hd__tap_1 TAP_11909 (  );
sky130_fd_sc_hd__tap_1 TAP_1191 (  );
sky130_fd_sc_hd__tap_1 TAP_11910 (  );
sky130_fd_sc_hd__tap_1 TAP_11911 (  );
sky130_fd_sc_hd__tap_1 TAP_11912 (  );
sky130_fd_sc_hd__tap_1 TAP_11913 (  );
sky130_fd_sc_hd__tap_1 TAP_11914 (  );
sky130_fd_sc_hd__tap_1 TAP_11915 (  );
sky130_fd_sc_hd__tap_1 TAP_11916 (  );
sky130_fd_sc_hd__tap_1 TAP_11917 (  );
sky130_fd_sc_hd__tap_1 TAP_11918 (  );
sky130_fd_sc_hd__tap_1 TAP_11919 (  );
sky130_fd_sc_hd__tap_1 TAP_1192 (  );
sky130_fd_sc_hd__tap_1 TAP_11920 (  );
sky130_fd_sc_hd__tap_1 TAP_11921 (  );
sky130_fd_sc_hd__tap_1 TAP_11922 (  );
sky130_fd_sc_hd__tap_1 TAP_11923 (  );
sky130_fd_sc_hd__tap_1 TAP_11924 (  );
sky130_fd_sc_hd__tap_1 TAP_11925 (  );
sky130_fd_sc_hd__tap_1 TAP_11926 (  );
sky130_fd_sc_hd__tap_1 TAP_11927 (  );
sky130_fd_sc_hd__tap_1 TAP_11928 (  );
sky130_fd_sc_hd__tap_1 TAP_11929 (  );
sky130_fd_sc_hd__tap_1 TAP_1193 (  );
sky130_fd_sc_hd__tap_1 TAP_11930 (  );
sky130_fd_sc_hd__tap_1 TAP_11931 (  );
sky130_fd_sc_hd__tap_1 TAP_11932 (  );
sky130_fd_sc_hd__tap_1 TAP_11933 (  );
sky130_fd_sc_hd__tap_1 TAP_11934 (  );
sky130_fd_sc_hd__tap_1 TAP_11935 (  );
sky130_fd_sc_hd__tap_1 TAP_11936 (  );
sky130_fd_sc_hd__tap_1 TAP_11937 (  );
sky130_fd_sc_hd__tap_1 TAP_11938 (  );
sky130_fd_sc_hd__tap_1 TAP_11939 (  );
sky130_fd_sc_hd__tap_1 TAP_1194 (  );
sky130_fd_sc_hd__tap_1 TAP_11940 (  );
sky130_fd_sc_hd__tap_1 TAP_11941 (  );
sky130_fd_sc_hd__tap_1 TAP_11942 (  );
sky130_fd_sc_hd__tap_1 TAP_11943 (  );
sky130_fd_sc_hd__tap_1 TAP_11944 (  );
sky130_fd_sc_hd__tap_1 TAP_11945 (  );
sky130_fd_sc_hd__tap_1 TAP_11946 (  );
sky130_fd_sc_hd__tap_1 TAP_11947 (  );
sky130_fd_sc_hd__tap_1 TAP_11948 (  );
sky130_fd_sc_hd__tap_1 TAP_11949 (  );
sky130_fd_sc_hd__tap_1 TAP_1195 (  );
sky130_fd_sc_hd__tap_1 TAP_11950 (  );
sky130_fd_sc_hd__tap_1 TAP_11951 (  );
sky130_fd_sc_hd__tap_1 TAP_11952 (  );
sky130_fd_sc_hd__tap_1 TAP_11953 (  );
sky130_fd_sc_hd__tap_1 TAP_11954 (  );
sky130_fd_sc_hd__tap_1 TAP_11955 (  );
sky130_fd_sc_hd__tap_1 TAP_11956 (  );
sky130_fd_sc_hd__tap_1 TAP_11957 (  );
sky130_fd_sc_hd__tap_1 TAP_11958 (  );
sky130_fd_sc_hd__tap_1 TAP_11959 (  );
sky130_fd_sc_hd__tap_1 TAP_1196 (  );
sky130_fd_sc_hd__tap_1 TAP_11960 (  );
sky130_fd_sc_hd__tap_1 TAP_11961 (  );
sky130_fd_sc_hd__tap_1 TAP_11962 (  );
sky130_fd_sc_hd__tap_1 TAP_11963 (  );
sky130_fd_sc_hd__tap_1 TAP_11964 (  );
sky130_fd_sc_hd__tap_1 TAP_11965 (  );
sky130_fd_sc_hd__tap_1 TAP_11966 (  );
sky130_fd_sc_hd__tap_1 TAP_11967 (  );
sky130_fd_sc_hd__tap_1 TAP_11968 (  );
sky130_fd_sc_hd__tap_1 TAP_11969 (  );
sky130_fd_sc_hd__tap_1 TAP_1197 (  );
sky130_fd_sc_hd__tap_1 TAP_11970 (  );
sky130_fd_sc_hd__tap_1 TAP_11971 (  );
sky130_fd_sc_hd__tap_1 TAP_11972 (  );
sky130_fd_sc_hd__tap_1 TAP_11973 (  );
sky130_fd_sc_hd__tap_1 TAP_11974 (  );
sky130_fd_sc_hd__tap_1 TAP_11975 (  );
sky130_fd_sc_hd__tap_1 TAP_11976 (  );
sky130_fd_sc_hd__tap_1 TAP_11977 (  );
sky130_fd_sc_hd__tap_1 TAP_11978 (  );
sky130_fd_sc_hd__tap_1 TAP_11979 (  );
sky130_fd_sc_hd__tap_1 TAP_1198 (  );
sky130_fd_sc_hd__tap_1 TAP_11980 (  );
sky130_fd_sc_hd__tap_1 TAP_11981 (  );
sky130_fd_sc_hd__tap_1 TAP_11982 (  );
sky130_fd_sc_hd__tap_1 TAP_11983 (  );
sky130_fd_sc_hd__tap_1 TAP_11984 (  );
sky130_fd_sc_hd__tap_1 TAP_11985 (  );
sky130_fd_sc_hd__tap_1 TAP_11986 (  );
sky130_fd_sc_hd__tap_1 TAP_11987 (  );
sky130_fd_sc_hd__tap_1 TAP_11988 (  );
sky130_fd_sc_hd__tap_1 TAP_11989 (  );
sky130_fd_sc_hd__tap_1 TAP_1199 (  );
sky130_fd_sc_hd__tap_1 TAP_11990 (  );
sky130_fd_sc_hd__tap_1 TAP_11991 (  );
sky130_fd_sc_hd__tap_1 TAP_11992 (  );
sky130_fd_sc_hd__tap_1 TAP_11993 (  );
sky130_fd_sc_hd__tap_1 TAP_11994 (  );
sky130_fd_sc_hd__tap_1 TAP_11995 (  );
sky130_fd_sc_hd__tap_1 TAP_11996 (  );
sky130_fd_sc_hd__tap_1 TAP_11997 (  );
sky130_fd_sc_hd__tap_1 TAP_11998 (  );
sky130_fd_sc_hd__tap_1 TAP_11999 (  );
sky130_fd_sc_hd__tap_1 TAP_1200 (  );
sky130_fd_sc_hd__tap_1 TAP_12000 (  );
sky130_fd_sc_hd__tap_1 TAP_12001 (  );
sky130_fd_sc_hd__tap_1 TAP_12002 (  );
sky130_fd_sc_hd__tap_1 TAP_12003 (  );
sky130_fd_sc_hd__tap_1 TAP_12004 (  );
sky130_fd_sc_hd__tap_1 TAP_12005 (  );
sky130_fd_sc_hd__tap_1 TAP_12006 (  );
sky130_fd_sc_hd__tap_1 TAP_12007 (  );
sky130_fd_sc_hd__tap_1 TAP_12008 (  );
sky130_fd_sc_hd__tap_1 TAP_12009 (  );
sky130_fd_sc_hd__tap_1 TAP_1201 (  );
sky130_fd_sc_hd__tap_1 TAP_12010 (  );
sky130_fd_sc_hd__tap_1 TAP_12011 (  );
sky130_fd_sc_hd__tap_1 TAP_12012 (  );
sky130_fd_sc_hd__tap_1 TAP_12013 (  );
sky130_fd_sc_hd__tap_1 TAP_12014 (  );
sky130_fd_sc_hd__tap_1 TAP_12015 (  );
sky130_fd_sc_hd__tap_1 TAP_12016 (  );
sky130_fd_sc_hd__tap_1 TAP_12017 (  );
sky130_fd_sc_hd__tap_1 TAP_12018 (  );
sky130_fd_sc_hd__tap_1 TAP_12019 (  );
sky130_fd_sc_hd__tap_1 TAP_1202 (  );
sky130_fd_sc_hd__tap_1 TAP_12020 (  );
sky130_fd_sc_hd__tap_1 TAP_12021 (  );
sky130_fd_sc_hd__tap_1 TAP_12022 (  );
sky130_fd_sc_hd__tap_1 TAP_12023 (  );
sky130_fd_sc_hd__tap_1 TAP_12024 (  );
sky130_fd_sc_hd__tap_1 TAP_12025 (  );
sky130_fd_sc_hd__tap_1 TAP_12026 (  );
sky130_fd_sc_hd__tap_1 TAP_12027 (  );
sky130_fd_sc_hd__tap_1 TAP_12028 (  );
sky130_fd_sc_hd__tap_1 TAP_12029 (  );
sky130_fd_sc_hd__tap_1 TAP_1203 (  );
sky130_fd_sc_hd__tap_1 TAP_12030 (  );
sky130_fd_sc_hd__tap_1 TAP_12031 (  );
sky130_fd_sc_hd__tap_1 TAP_12032 (  );
sky130_fd_sc_hd__tap_1 TAP_12033 (  );
sky130_fd_sc_hd__tap_1 TAP_12034 (  );
sky130_fd_sc_hd__tap_1 TAP_12035 (  );
sky130_fd_sc_hd__tap_1 TAP_12036 (  );
sky130_fd_sc_hd__tap_1 TAP_12037 (  );
sky130_fd_sc_hd__tap_1 TAP_12038 (  );
sky130_fd_sc_hd__tap_1 TAP_12039 (  );
sky130_fd_sc_hd__tap_1 TAP_1204 (  );
sky130_fd_sc_hd__tap_1 TAP_12040 (  );
sky130_fd_sc_hd__tap_1 TAP_12041 (  );
sky130_fd_sc_hd__tap_1 TAP_12042 (  );
sky130_fd_sc_hd__tap_1 TAP_12043 (  );
sky130_fd_sc_hd__tap_1 TAP_12044 (  );
sky130_fd_sc_hd__tap_1 TAP_12045 (  );
sky130_fd_sc_hd__tap_1 TAP_12046 (  );
sky130_fd_sc_hd__tap_1 TAP_12047 (  );
sky130_fd_sc_hd__tap_1 TAP_12048 (  );
sky130_fd_sc_hd__tap_1 TAP_12049 (  );
sky130_fd_sc_hd__tap_1 TAP_1205 (  );
sky130_fd_sc_hd__tap_1 TAP_12050 (  );
sky130_fd_sc_hd__tap_1 TAP_12051 (  );
sky130_fd_sc_hd__tap_1 TAP_12052 (  );
sky130_fd_sc_hd__tap_1 TAP_12053 (  );
sky130_fd_sc_hd__tap_1 TAP_12054 (  );
sky130_fd_sc_hd__tap_1 TAP_12055 (  );
sky130_fd_sc_hd__tap_1 TAP_12056 (  );
sky130_fd_sc_hd__tap_1 TAP_12057 (  );
sky130_fd_sc_hd__tap_1 TAP_12058 (  );
sky130_fd_sc_hd__tap_1 TAP_12059 (  );
sky130_fd_sc_hd__tap_1 TAP_1206 (  );
sky130_fd_sc_hd__tap_1 TAP_12060 (  );
sky130_fd_sc_hd__tap_1 TAP_12061 (  );
sky130_fd_sc_hd__tap_1 TAP_12062 (  );
sky130_fd_sc_hd__tap_1 TAP_12063 (  );
sky130_fd_sc_hd__tap_1 TAP_12064 (  );
sky130_fd_sc_hd__tap_1 TAP_12065 (  );
sky130_fd_sc_hd__tap_1 TAP_12066 (  );
sky130_fd_sc_hd__tap_1 TAP_12067 (  );
sky130_fd_sc_hd__tap_1 TAP_12068 (  );
sky130_fd_sc_hd__tap_1 TAP_12069 (  );
sky130_fd_sc_hd__tap_1 TAP_1207 (  );
sky130_fd_sc_hd__tap_1 TAP_12070 (  );
sky130_fd_sc_hd__tap_1 TAP_12071 (  );
sky130_fd_sc_hd__tap_1 TAP_12072 (  );
sky130_fd_sc_hd__tap_1 TAP_12073 (  );
sky130_fd_sc_hd__tap_1 TAP_12074 (  );
sky130_fd_sc_hd__tap_1 TAP_12075 (  );
sky130_fd_sc_hd__tap_1 TAP_12076 (  );
sky130_fd_sc_hd__tap_1 TAP_12077 (  );
sky130_fd_sc_hd__tap_1 TAP_12078 (  );
sky130_fd_sc_hd__tap_1 TAP_12079 (  );
sky130_fd_sc_hd__tap_1 TAP_1208 (  );
sky130_fd_sc_hd__tap_1 TAP_12080 (  );
sky130_fd_sc_hd__tap_1 TAP_12081 (  );
sky130_fd_sc_hd__tap_1 TAP_12082 (  );
sky130_fd_sc_hd__tap_1 TAP_12083 (  );
sky130_fd_sc_hd__tap_1 TAP_12084 (  );
sky130_fd_sc_hd__tap_1 TAP_12085 (  );
sky130_fd_sc_hd__tap_1 TAP_12086 (  );
sky130_fd_sc_hd__tap_1 TAP_12087 (  );
sky130_fd_sc_hd__tap_1 TAP_12088 (  );
sky130_fd_sc_hd__tap_1 TAP_12089 (  );
sky130_fd_sc_hd__tap_1 TAP_1209 (  );
sky130_fd_sc_hd__tap_1 TAP_12090 (  );
sky130_fd_sc_hd__tap_1 TAP_12091 (  );
sky130_fd_sc_hd__tap_1 TAP_12092 (  );
sky130_fd_sc_hd__tap_1 TAP_12093 (  );
sky130_fd_sc_hd__tap_1 TAP_12094 (  );
sky130_fd_sc_hd__tap_1 TAP_12095 (  );
sky130_fd_sc_hd__tap_1 TAP_12096 (  );
sky130_fd_sc_hd__tap_1 TAP_12097 (  );
sky130_fd_sc_hd__tap_1 TAP_12098 (  );
sky130_fd_sc_hd__tap_1 TAP_12099 (  );
sky130_fd_sc_hd__tap_1 TAP_1210 (  );
sky130_fd_sc_hd__tap_1 TAP_12100 (  );
sky130_fd_sc_hd__tap_1 TAP_12101 (  );
sky130_fd_sc_hd__tap_1 TAP_12102 (  );
sky130_fd_sc_hd__tap_1 TAP_12103 (  );
sky130_fd_sc_hd__tap_1 TAP_12104 (  );
sky130_fd_sc_hd__tap_1 TAP_12105 (  );
sky130_fd_sc_hd__tap_1 TAP_12106 (  );
sky130_fd_sc_hd__tap_1 TAP_12107 (  );
sky130_fd_sc_hd__tap_1 TAP_12108 (  );
sky130_fd_sc_hd__tap_1 TAP_12109 (  );
sky130_fd_sc_hd__tap_1 TAP_1211 (  );
sky130_fd_sc_hd__tap_1 TAP_12110 (  );
sky130_fd_sc_hd__tap_1 TAP_12111 (  );
sky130_fd_sc_hd__tap_1 TAP_12112 (  );
sky130_fd_sc_hd__tap_1 TAP_12113 (  );
sky130_fd_sc_hd__tap_1 TAP_12114 (  );
sky130_fd_sc_hd__tap_1 TAP_12115 (  );
sky130_fd_sc_hd__tap_1 TAP_12116 (  );
sky130_fd_sc_hd__tap_1 TAP_12117 (  );
sky130_fd_sc_hd__tap_1 TAP_12118 (  );
sky130_fd_sc_hd__tap_1 TAP_12119 (  );
sky130_fd_sc_hd__tap_1 TAP_1212 (  );
sky130_fd_sc_hd__tap_1 TAP_12120 (  );
sky130_fd_sc_hd__tap_1 TAP_12121 (  );
sky130_fd_sc_hd__tap_1 TAP_12122 (  );
sky130_fd_sc_hd__tap_1 TAP_12123 (  );
sky130_fd_sc_hd__tap_1 TAP_12124 (  );
sky130_fd_sc_hd__tap_1 TAP_12125 (  );
sky130_fd_sc_hd__tap_1 TAP_12126 (  );
sky130_fd_sc_hd__tap_1 TAP_12127 (  );
sky130_fd_sc_hd__tap_1 TAP_12128 (  );
sky130_fd_sc_hd__tap_1 TAP_12129 (  );
sky130_fd_sc_hd__tap_1 TAP_1213 (  );
sky130_fd_sc_hd__tap_1 TAP_12130 (  );
sky130_fd_sc_hd__tap_1 TAP_12131 (  );
sky130_fd_sc_hd__tap_1 TAP_12132 (  );
sky130_fd_sc_hd__tap_1 TAP_12133 (  );
sky130_fd_sc_hd__tap_1 TAP_12134 (  );
sky130_fd_sc_hd__tap_1 TAP_12135 (  );
sky130_fd_sc_hd__tap_1 TAP_12136 (  );
sky130_fd_sc_hd__tap_1 TAP_12137 (  );
sky130_fd_sc_hd__tap_1 TAP_12138 (  );
sky130_fd_sc_hd__tap_1 TAP_12139 (  );
sky130_fd_sc_hd__tap_1 TAP_1214 (  );
sky130_fd_sc_hd__tap_1 TAP_12140 (  );
sky130_fd_sc_hd__tap_1 TAP_12141 (  );
sky130_fd_sc_hd__tap_1 TAP_12142 (  );
sky130_fd_sc_hd__tap_1 TAP_12143 (  );
sky130_fd_sc_hd__tap_1 TAP_12144 (  );
sky130_fd_sc_hd__tap_1 TAP_12145 (  );
sky130_fd_sc_hd__tap_1 TAP_12146 (  );
sky130_fd_sc_hd__tap_1 TAP_12147 (  );
sky130_fd_sc_hd__tap_1 TAP_12148 (  );
sky130_fd_sc_hd__tap_1 TAP_12149 (  );
sky130_fd_sc_hd__tap_1 TAP_1215 (  );
sky130_fd_sc_hd__tap_1 TAP_12150 (  );
sky130_fd_sc_hd__tap_1 TAP_12151 (  );
sky130_fd_sc_hd__tap_1 TAP_12152 (  );
sky130_fd_sc_hd__tap_1 TAP_12153 (  );
sky130_fd_sc_hd__tap_1 TAP_12154 (  );
sky130_fd_sc_hd__tap_1 TAP_12155 (  );
sky130_fd_sc_hd__tap_1 TAP_12156 (  );
sky130_fd_sc_hd__tap_1 TAP_12157 (  );
sky130_fd_sc_hd__tap_1 TAP_12158 (  );
sky130_fd_sc_hd__tap_1 TAP_12159 (  );
sky130_fd_sc_hd__tap_1 TAP_1216 (  );
sky130_fd_sc_hd__tap_1 TAP_12160 (  );
sky130_fd_sc_hd__tap_1 TAP_12161 (  );
sky130_fd_sc_hd__tap_1 TAP_12162 (  );
sky130_fd_sc_hd__tap_1 TAP_12163 (  );
sky130_fd_sc_hd__tap_1 TAP_12164 (  );
sky130_fd_sc_hd__tap_1 TAP_12165 (  );
sky130_fd_sc_hd__tap_1 TAP_12166 (  );
sky130_fd_sc_hd__tap_1 TAP_12167 (  );
sky130_fd_sc_hd__tap_1 TAP_12168 (  );
sky130_fd_sc_hd__tap_1 TAP_12169 (  );
sky130_fd_sc_hd__tap_1 TAP_1217 (  );
sky130_fd_sc_hd__tap_1 TAP_12170 (  );
sky130_fd_sc_hd__tap_1 TAP_12171 (  );
sky130_fd_sc_hd__tap_1 TAP_12172 (  );
sky130_fd_sc_hd__tap_1 TAP_12173 (  );
sky130_fd_sc_hd__tap_1 TAP_12174 (  );
sky130_fd_sc_hd__tap_1 TAP_12175 (  );
sky130_fd_sc_hd__tap_1 TAP_12176 (  );
sky130_fd_sc_hd__tap_1 TAP_12177 (  );
sky130_fd_sc_hd__tap_1 TAP_12178 (  );
sky130_fd_sc_hd__tap_1 TAP_12179 (  );
sky130_fd_sc_hd__tap_1 TAP_1218 (  );
sky130_fd_sc_hd__tap_1 TAP_12180 (  );
sky130_fd_sc_hd__tap_1 TAP_12181 (  );
sky130_fd_sc_hd__tap_1 TAP_12182 (  );
sky130_fd_sc_hd__tap_1 TAP_12183 (  );
sky130_fd_sc_hd__tap_1 TAP_12184 (  );
sky130_fd_sc_hd__tap_1 TAP_12185 (  );
sky130_fd_sc_hd__tap_1 TAP_12186 (  );
sky130_fd_sc_hd__tap_1 TAP_12187 (  );
sky130_fd_sc_hd__tap_1 TAP_12188 (  );
sky130_fd_sc_hd__tap_1 TAP_12189 (  );
sky130_fd_sc_hd__tap_1 TAP_1219 (  );
sky130_fd_sc_hd__tap_1 TAP_12190 (  );
sky130_fd_sc_hd__tap_1 TAP_12191 (  );
sky130_fd_sc_hd__tap_1 TAP_12192 (  );
sky130_fd_sc_hd__tap_1 TAP_12193 (  );
sky130_fd_sc_hd__tap_1 TAP_12194 (  );
sky130_fd_sc_hd__tap_1 TAP_12195 (  );
sky130_fd_sc_hd__tap_1 TAP_12196 (  );
sky130_fd_sc_hd__tap_1 TAP_12197 (  );
sky130_fd_sc_hd__tap_1 TAP_12198 (  );
sky130_fd_sc_hd__tap_1 TAP_12199 (  );
sky130_fd_sc_hd__tap_1 TAP_1220 (  );
sky130_fd_sc_hd__tap_1 TAP_12200 (  );
sky130_fd_sc_hd__tap_1 TAP_12201 (  );
sky130_fd_sc_hd__tap_1 TAP_12202 (  );
sky130_fd_sc_hd__tap_1 TAP_12203 (  );
sky130_fd_sc_hd__tap_1 TAP_12204 (  );
sky130_fd_sc_hd__tap_1 TAP_12205 (  );
sky130_fd_sc_hd__tap_1 TAP_12206 (  );
sky130_fd_sc_hd__tap_1 TAP_12207 (  );
sky130_fd_sc_hd__tap_1 TAP_12208 (  );
sky130_fd_sc_hd__tap_1 TAP_12209 (  );
sky130_fd_sc_hd__tap_1 TAP_1221 (  );
sky130_fd_sc_hd__tap_1 TAP_12210 (  );
sky130_fd_sc_hd__tap_1 TAP_12211 (  );
sky130_fd_sc_hd__tap_1 TAP_12212 (  );
sky130_fd_sc_hd__tap_1 TAP_12213 (  );
sky130_fd_sc_hd__tap_1 TAP_12214 (  );
sky130_fd_sc_hd__tap_1 TAP_12215 (  );
sky130_fd_sc_hd__tap_1 TAP_12216 (  );
sky130_fd_sc_hd__tap_1 TAP_12217 (  );
sky130_fd_sc_hd__tap_1 TAP_12218 (  );
sky130_fd_sc_hd__tap_1 TAP_12219 (  );
sky130_fd_sc_hd__tap_1 TAP_1222 (  );
sky130_fd_sc_hd__tap_1 TAP_12220 (  );
sky130_fd_sc_hd__tap_1 TAP_12221 (  );
sky130_fd_sc_hd__tap_1 TAP_12222 (  );
sky130_fd_sc_hd__tap_1 TAP_12223 (  );
sky130_fd_sc_hd__tap_1 TAP_12224 (  );
sky130_fd_sc_hd__tap_1 TAP_12225 (  );
sky130_fd_sc_hd__tap_1 TAP_12226 (  );
sky130_fd_sc_hd__tap_1 TAP_12227 (  );
sky130_fd_sc_hd__tap_1 TAP_12228 (  );
sky130_fd_sc_hd__tap_1 TAP_12229 (  );
sky130_fd_sc_hd__tap_1 TAP_1223 (  );
sky130_fd_sc_hd__tap_1 TAP_12230 (  );
sky130_fd_sc_hd__tap_1 TAP_12231 (  );
sky130_fd_sc_hd__tap_1 TAP_12232 (  );
sky130_fd_sc_hd__tap_1 TAP_12233 (  );
sky130_fd_sc_hd__tap_1 TAP_12234 (  );
sky130_fd_sc_hd__tap_1 TAP_12235 (  );
sky130_fd_sc_hd__tap_1 TAP_12236 (  );
sky130_fd_sc_hd__tap_1 TAP_12237 (  );
sky130_fd_sc_hd__tap_1 TAP_12238 (  );
sky130_fd_sc_hd__tap_1 TAP_12239 (  );
sky130_fd_sc_hd__tap_1 TAP_1224 (  );
sky130_fd_sc_hd__tap_1 TAP_12240 (  );
sky130_fd_sc_hd__tap_1 TAP_12241 (  );
sky130_fd_sc_hd__tap_1 TAP_12242 (  );
sky130_fd_sc_hd__tap_1 TAP_12243 (  );
sky130_fd_sc_hd__tap_1 TAP_12244 (  );
sky130_fd_sc_hd__tap_1 TAP_12245 (  );
sky130_fd_sc_hd__tap_1 TAP_12246 (  );
sky130_fd_sc_hd__tap_1 TAP_12247 (  );
sky130_fd_sc_hd__tap_1 TAP_12248 (  );
sky130_fd_sc_hd__tap_1 TAP_12249 (  );
sky130_fd_sc_hd__tap_1 TAP_1225 (  );
sky130_fd_sc_hd__tap_1 TAP_12250 (  );
sky130_fd_sc_hd__tap_1 TAP_12251 (  );
sky130_fd_sc_hd__tap_1 TAP_12252 (  );
sky130_fd_sc_hd__tap_1 TAP_12253 (  );
sky130_fd_sc_hd__tap_1 TAP_12254 (  );
sky130_fd_sc_hd__tap_1 TAP_12255 (  );
sky130_fd_sc_hd__tap_1 TAP_12256 (  );
sky130_fd_sc_hd__tap_1 TAP_12257 (  );
sky130_fd_sc_hd__tap_1 TAP_12258 (  );
sky130_fd_sc_hd__tap_1 TAP_12259 (  );
sky130_fd_sc_hd__tap_1 TAP_1226 (  );
sky130_fd_sc_hd__tap_1 TAP_12260 (  );
sky130_fd_sc_hd__tap_1 TAP_12261 (  );
sky130_fd_sc_hd__tap_1 TAP_12262 (  );
sky130_fd_sc_hd__tap_1 TAP_12263 (  );
sky130_fd_sc_hd__tap_1 TAP_12264 (  );
sky130_fd_sc_hd__tap_1 TAP_12265 (  );
sky130_fd_sc_hd__tap_1 TAP_12266 (  );
sky130_fd_sc_hd__tap_1 TAP_12267 (  );
sky130_fd_sc_hd__tap_1 TAP_12268 (  );
sky130_fd_sc_hd__tap_1 TAP_12269 (  );
sky130_fd_sc_hd__tap_1 TAP_1227 (  );
sky130_fd_sc_hd__tap_1 TAP_12270 (  );
sky130_fd_sc_hd__tap_1 TAP_12271 (  );
sky130_fd_sc_hd__tap_1 TAP_12272 (  );
sky130_fd_sc_hd__tap_1 TAP_12273 (  );
sky130_fd_sc_hd__tap_1 TAP_12274 (  );
sky130_fd_sc_hd__tap_1 TAP_12275 (  );
sky130_fd_sc_hd__tap_1 TAP_12276 (  );
sky130_fd_sc_hd__tap_1 TAP_12277 (  );
sky130_fd_sc_hd__tap_1 TAP_12278 (  );
sky130_fd_sc_hd__tap_1 TAP_12279 (  );
sky130_fd_sc_hd__tap_1 TAP_1228 (  );
sky130_fd_sc_hd__tap_1 TAP_12280 (  );
sky130_fd_sc_hd__tap_1 TAP_12281 (  );
sky130_fd_sc_hd__tap_1 TAP_12282 (  );
sky130_fd_sc_hd__tap_1 TAP_12283 (  );
sky130_fd_sc_hd__tap_1 TAP_12284 (  );
sky130_fd_sc_hd__tap_1 TAP_12285 (  );
sky130_fd_sc_hd__tap_1 TAP_12286 (  );
sky130_fd_sc_hd__tap_1 TAP_12287 (  );
sky130_fd_sc_hd__tap_1 TAP_12288 (  );
sky130_fd_sc_hd__tap_1 TAP_12289 (  );
sky130_fd_sc_hd__tap_1 TAP_1229 (  );
sky130_fd_sc_hd__tap_1 TAP_12290 (  );
sky130_fd_sc_hd__tap_1 TAP_12291 (  );
sky130_fd_sc_hd__tap_1 TAP_12292 (  );
sky130_fd_sc_hd__tap_1 TAP_12293 (  );
sky130_fd_sc_hd__tap_1 TAP_12294 (  );
sky130_fd_sc_hd__tap_1 TAP_12295 (  );
sky130_fd_sc_hd__tap_1 TAP_12296 (  );
sky130_fd_sc_hd__tap_1 TAP_12297 (  );
sky130_fd_sc_hd__tap_1 TAP_12298 (  );
sky130_fd_sc_hd__tap_1 TAP_12299 (  );
sky130_fd_sc_hd__tap_1 TAP_1230 (  );
sky130_fd_sc_hd__tap_1 TAP_12300 (  );
sky130_fd_sc_hd__tap_1 TAP_12301 (  );
sky130_fd_sc_hd__tap_1 TAP_12302 (  );
sky130_fd_sc_hd__tap_1 TAP_12303 (  );
sky130_fd_sc_hd__tap_1 TAP_12304 (  );
sky130_fd_sc_hd__tap_1 TAP_12305 (  );
sky130_fd_sc_hd__tap_1 TAP_12306 (  );
sky130_fd_sc_hd__tap_1 TAP_12307 (  );
sky130_fd_sc_hd__tap_1 TAP_12308 (  );
sky130_fd_sc_hd__tap_1 TAP_12309 (  );
sky130_fd_sc_hd__tap_1 TAP_1231 (  );
sky130_fd_sc_hd__tap_1 TAP_12310 (  );
sky130_fd_sc_hd__tap_1 TAP_12311 (  );
sky130_fd_sc_hd__tap_1 TAP_12312 (  );
sky130_fd_sc_hd__tap_1 TAP_12313 (  );
sky130_fd_sc_hd__tap_1 TAP_12314 (  );
sky130_fd_sc_hd__tap_1 TAP_12315 (  );
sky130_fd_sc_hd__tap_1 TAP_12316 (  );
sky130_fd_sc_hd__tap_1 TAP_12317 (  );
sky130_fd_sc_hd__tap_1 TAP_12318 (  );
sky130_fd_sc_hd__tap_1 TAP_12319 (  );
sky130_fd_sc_hd__tap_1 TAP_1232 (  );
sky130_fd_sc_hd__tap_1 TAP_12320 (  );
sky130_fd_sc_hd__tap_1 TAP_12321 (  );
sky130_fd_sc_hd__tap_1 TAP_12322 (  );
sky130_fd_sc_hd__tap_1 TAP_12323 (  );
sky130_fd_sc_hd__tap_1 TAP_12324 (  );
sky130_fd_sc_hd__tap_1 TAP_12325 (  );
sky130_fd_sc_hd__tap_1 TAP_12326 (  );
sky130_fd_sc_hd__tap_1 TAP_12327 (  );
sky130_fd_sc_hd__tap_1 TAP_12328 (  );
sky130_fd_sc_hd__tap_1 TAP_12329 (  );
sky130_fd_sc_hd__tap_1 TAP_1233 (  );
sky130_fd_sc_hd__tap_1 TAP_12330 (  );
sky130_fd_sc_hd__tap_1 TAP_12331 (  );
sky130_fd_sc_hd__tap_1 TAP_12332 (  );
sky130_fd_sc_hd__tap_1 TAP_12333 (  );
sky130_fd_sc_hd__tap_1 TAP_12334 (  );
sky130_fd_sc_hd__tap_1 TAP_12335 (  );
sky130_fd_sc_hd__tap_1 TAP_12336 (  );
sky130_fd_sc_hd__tap_1 TAP_12337 (  );
sky130_fd_sc_hd__tap_1 TAP_12338 (  );
sky130_fd_sc_hd__tap_1 TAP_12339 (  );
sky130_fd_sc_hd__tap_1 TAP_1234 (  );
sky130_fd_sc_hd__tap_1 TAP_12340 (  );
sky130_fd_sc_hd__tap_1 TAP_12341 (  );
sky130_fd_sc_hd__tap_1 TAP_12342 (  );
sky130_fd_sc_hd__tap_1 TAP_12343 (  );
sky130_fd_sc_hd__tap_1 TAP_12344 (  );
sky130_fd_sc_hd__tap_1 TAP_12345 (  );
sky130_fd_sc_hd__tap_1 TAP_12346 (  );
sky130_fd_sc_hd__tap_1 TAP_12347 (  );
sky130_fd_sc_hd__tap_1 TAP_12348 (  );
sky130_fd_sc_hd__tap_1 TAP_12349 (  );
sky130_fd_sc_hd__tap_1 TAP_1235 (  );
sky130_fd_sc_hd__tap_1 TAP_12350 (  );
sky130_fd_sc_hd__tap_1 TAP_12351 (  );
sky130_fd_sc_hd__tap_1 TAP_12352 (  );
sky130_fd_sc_hd__tap_1 TAP_12353 (  );
sky130_fd_sc_hd__tap_1 TAP_12354 (  );
sky130_fd_sc_hd__tap_1 TAP_12355 (  );
sky130_fd_sc_hd__tap_1 TAP_12356 (  );
sky130_fd_sc_hd__tap_1 TAP_12357 (  );
sky130_fd_sc_hd__tap_1 TAP_12358 (  );
sky130_fd_sc_hd__tap_1 TAP_12359 (  );
sky130_fd_sc_hd__tap_1 TAP_1236 (  );
sky130_fd_sc_hd__tap_1 TAP_12360 (  );
sky130_fd_sc_hd__tap_1 TAP_12361 (  );
sky130_fd_sc_hd__tap_1 TAP_12362 (  );
sky130_fd_sc_hd__tap_1 TAP_12363 (  );
sky130_fd_sc_hd__tap_1 TAP_12364 (  );
sky130_fd_sc_hd__tap_1 TAP_12365 (  );
sky130_fd_sc_hd__tap_1 TAP_12366 (  );
sky130_fd_sc_hd__tap_1 TAP_12367 (  );
sky130_fd_sc_hd__tap_1 TAP_12368 (  );
sky130_fd_sc_hd__tap_1 TAP_12369 (  );
sky130_fd_sc_hd__tap_1 TAP_1237 (  );
sky130_fd_sc_hd__tap_1 TAP_12370 (  );
sky130_fd_sc_hd__tap_1 TAP_12371 (  );
sky130_fd_sc_hd__tap_1 TAP_12372 (  );
sky130_fd_sc_hd__tap_1 TAP_12373 (  );
sky130_fd_sc_hd__tap_1 TAP_12374 (  );
sky130_fd_sc_hd__tap_1 TAP_12375 (  );
sky130_fd_sc_hd__tap_1 TAP_12376 (  );
sky130_fd_sc_hd__tap_1 TAP_12377 (  );
sky130_fd_sc_hd__tap_1 TAP_12378 (  );
sky130_fd_sc_hd__tap_1 TAP_12379 (  );
sky130_fd_sc_hd__tap_1 TAP_1238 (  );
sky130_fd_sc_hd__tap_1 TAP_12380 (  );
sky130_fd_sc_hd__tap_1 TAP_12381 (  );
sky130_fd_sc_hd__tap_1 TAP_12382 (  );
sky130_fd_sc_hd__tap_1 TAP_12383 (  );
sky130_fd_sc_hd__tap_1 TAP_12384 (  );
sky130_fd_sc_hd__tap_1 TAP_12385 (  );
sky130_fd_sc_hd__tap_1 TAP_12386 (  );
sky130_fd_sc_hd__tap_1 TAP_12387 (  );
sky130_fd_sc_hd__tap_1 TAP_12388 (  );
sky130_fd_sc_hd__tap_1 TAP_12389 (  );
sky130_fd_sc_hd__tap_1 TAP_1239 (  );
sky130_fd_sc_hd__tap_1 TAP_12390 (  );
sky130_fd_sc_hd__tap_1 TAP_12391 (  );
sky130_fd_sc_hd__tap_1 TAP_12392 (  );
sky130_fd_sc_hd__tap_1 TAP_12393 (  );
sky130_fd_sc_hd__tap_1 TAP_12394 (  );
sky130_fd_sc_hd__tap_1 TAP_12395 (  );
sky130_fd_sc_hd__tap_1 TAP_12396 (  );
sky130_fd_sc_hd__tap_1 TAP_12397 (  );
sky130_fd_sc_hd__tap_1 TAP_12398 (  );
sky130_fd_sc_hd__tap_1 TAP_12399 (  );
sky130_fd_sc_hd__tap_1 TAP_1240 (  );
sky130_fd_sc_hd__tap_1 TAP_12400 (  );
sky130_fd_sc_hd__tap_1 TAP_12401 (  );
sky130_fd_sc_hd__tap_1 TAP_12402 (  );
sky130_fd_sc_hd__tap_1 TAP_12403 (  );
sky130_fd_sc_hd__tap_1 TAP_12404 (  );
sky130_fd_sc_hd__tap_1 TAP_12405 (  );
sky130_fd_sc_hd__tap_1 TAP_12406 (  );
sky130_fd_sc_hd__tap_1 TAP_12407 (  );
sky130_fd_sc_hd__tap_1 TAP_12408 (  );
sky130_fd_sc_hd__tap_1 TAP_12409 (  );
sky130_fd_sc_hd__tap_1 TAP_1241 (  );
sky130_fd_sc_hd__tap_1 TAP_12410 (  );
sky130_fd_sc_hd__tap_1 TAP_12411 (  );
sky130_fd_sc_hd__tap_1 TAP_12412 (  );
sky130_fd_sc_hd__tap_1 TAP_12413 (  );
sky130_fd_sc_hd__tap_1 TAP_12414 (  );
sky130_fd_sc_hd__tap_1 TAP_12415 (  );
sky130_fd_sc_hd__tap_1 TAP_12416 (  );
sky130_fd_sc_hd__tap_1 TAP_12417 (  );
sky130_fd_sc_hd__tap_1 TAP_12418 (  );
sky130_fd_sc_hd__tap_1 TAP_12419 (  );
sky130_fd_sc_hd__tap_1 TAP_1242 (  );
sky130_fd_sc_hd__tap_1 TAP_12420 (  );
sky130_fd_sc_hd__tap_1 TAP_12421 (  );
sky130_fd_sc_hd__tap_1 TAP_12422 (  );
sky130_fd_sc_hd__tap_1 TAP_12423 (  );
sky130_fd_sc_hd__tap_1 TAP_12424 (  );
sky130_fd_sc_hd__tap_1 TAP_12425 (  );
sky130_fd_sc_hd__tap_1 TAP_12426 (  );
sky130_fd_sc_hd__tap_1 TAP_12427 (  );
sky130_fd_sc_hd__tap_1 TAP_12428 (  );
sky130_fd_sc_hd__tap_1 TAP_12429 (  );
sky130_fd_sc_hd__tap_1 TAP_1243 (  );
sky130_fd_sc_hd__tap_1 TAP_12430 (  );
sky130_fd_sc_hd__tap_1 TAP_12431 (  );
sky130_fd_sc_hd__tap_1 TAP_12432 (  );
sky130_fd_sc_hd__tap_1 TAP_12433 (  );
sky130_fd_sc_hd__tap_1 TAP_12434 (  );
sky130_fd_sc_hd__tap_1 TAP_12435 (  );
sky130_fd_sc_hd__tap_1 TAP_12436 (  );
sky130_fd_sc_hd__tap_1 TAP_12437 (  );
sky130_fd_sc_hd__tap_1 TAP_12438 (  );
sky130_fd_sc_hd__tap_1 TAP_12439 (  );
sky130_fd_sc_hd__tap_1 TAP_1244 (  );
sky130_fd_sc_hd__tap_1 TAP_12440 (  );
sky130_fd_sc_hd__tap_1 TAP_12441 (  );
sky130_fd_sc_hd__tap_1 TAP_12442 (  );
sky130_fd_sc_hd__tap_1 TAP_12443 (  );
sky130_fd_sc_hd__tap_1 TAP_12444 (  );
sky130_fd_sc_hd__tap_1 TAP_12445 (  );
sky130_fd_sc_hd__tap_1 TAP_12446 (  );
sky130_fd_sc_hd__tap_1 TAP_12447 (  );
sky130_fd_sc_hd__tap_1 TAP_12448 (  );
sky130_fd_sc_hd__tap_1 TAP_12449 (  );
sky130_fd_sc_hd__tap_1 TAP_1245 (  );
sky130_fd_sc_hd__tap_1 TAP_12450 (  );
sky130_fd_sc_hd__tap_1 TAP_12451 (  );
sky130_fd_sc_hd__tap_1 TAP_12452 (  );
sky130_fd_sc_hd__tap_1 TAP_12453 (  );
sky130_fd_sc_hd__tap_1 TAP_12454 (  );
sky130_fd_sc_hd__tap_1 TAP_12455 (  );
sky130_fd_sc_hd__tap_1 TAP_12456 (  );
sky130_fd_sc_hd__tap_1 TAP_12457 (  );
sky130_fd_sc_hd__tap_1 TAP_12458 (  );
sky130_fd_sc_hd__tap_1 TAP_12459 (  );
sky130_fd_sc_hd__tap_1 TAP_1246 (  );
sky130_fd_sc_hd__tap_1 TAP_12460 (  );
sky130_fd_sc_hd__tap_1 TAP_12461 (  );
sky130_fd_sc_hd__tap_1 TAP_12462 (  );
sky130_fd_sc_hd__tap_1 TAP_12463 (  );
sky130_fd_sc_hd__tap_1 TAP_12464 (  );
sky130_fd_sc_hd__tap_1 TAP_12465 (  );
sky130_fd_sc_hd__tap_1 TAP_12466 (  );
sky130_fd_sc_hd__tap_1 TAP_12467 (  );
sky130_fd_sc_hd__tap_1 TAP_12468 (  );
sky130_fd_sc_hd__tap_1 TAP_12469 (  );
sky130_fd_sc_hd__tap_1 TAP_1247 (  );
sky130_fd_sc_hd__tap_1 TAP_12470 (  );
sky130_fd_sc_hd__tap_1 TAP_12471 (  );
sky130_fd_sc_hd__tap_1 TAP_12472 (  );
sky130_fd_sc_hd__tap_1 TAP_12473 (  );
sky130_fd_sc_hd__tap_1 TAP_12474 (  );
sky130_fd_sc_hd__tap_1 TAP_12475 (  );
sky130_fd_sc_hd__tap_1 TAP_12476 (  );
sky130_fd_sc_hd__tap_1 TAP_12477 (  );
sky130_fd_sc_hd__tap_1 TAP_12478 (  );
sky130_fd_sc_hd__tap_1 TAP_12479 (  );
sky130_fd_sc_hd__tap_1 TAP_1248 (  );
sky130_fd_sc_hd__tap_1 TAP_12480 (  );
sky130_fd_sc_hd__tap_1 TAP_12481 (  );
sky130_fd_sc_hd__tap_1 TAP_12482 (  );
sky130_fd_sc_hd__tap_1 TAP_12483 (  );
sky130_fd_sc_hd__tap_1 TAP_12484 (  );
sky130_fd_sc_hd__tap_1 TAP_12485 (  );
sky130_fd_sc_hd__tap_1 TAP_12486 (  );
sky130_fd_sc_hd__tap_1 TAP_12487 (  );
sky130_fd_sc_hd__tap_1 TAP_12488 (  );
sky130_fd_sc_hd__tap_1 TAP_12489 (  );
sky130_fd_sc_hd__tap_1 TAP_1249 (  );
sky130_fd_sc_hd__tap_1 TAP_12490 (  );
sky130_fd_sc_hd__tap_1 TAP_12491 (  );
sky130_fd_sc_hd__tap_1 TAP_12492 (  );
sky130_fd_sc_hd__tap_1 TAP_12493 (  );
sky130_fd_sc_hd__tap_1 TAP_12494 (  );
sky130_fd_sc_hd__tap_1 TAP_12495 (  );
sky130_fd_sc_hd__tap_1 TAP_12496 (  );
sky130_fd_sc_hd__tap_1 TAP_12497 (  );
sky130_fd_sc_hd__tap_1 TAP_12498 (  );
sky130_fd_sc_hd__tap_1 TAP_12499 (  );
sky130_fd_sc_hd__tap_1 TAP_1250 (  );
sky130_fd_sc_hd__tap_1 TAP_12500 (  );
sky130_fd_sc_hd__tap_1 TAP_12501 (  );
sky130_fd_sc_hd__tap_1 TAP_12502 (  );
sky130_fd_sc_hd__tap_1 TAP_12503 (  );
sky130_fd_sc_hd__tap_1 TAP_12504 (  );
sky130_fd_sc_hd__tap_1 TAP_12505 (  );
sky130_fd_sc_hd__tap_1 TAP_12506 (  );
sky130_fd_sc_hd__tap_1 TAP_12507 (  );
sky130_fd_sc_hd__tap_1 TAP_12508 (  );
sky130_fd_sc_hd__tap_1 TAP_12509 (  );
sky130_fd_sc_hd__tap_1 TAP_1251 (  );
sky130_fd_sc_hd__tap_1 TAP_12510 (  );
sky130_fd_sc_hd__tap_1 TAP_12511 (  );
sky130_fd_sc_hd__tap_1 TAP_12512 (  );
sky130_fd_sc_hd__tap_1 TAP_12513 (  );
sky130_fd_sc_hd__tap_1 TAP_12514 (  );
sky130_fd_sc_hd__tap_1 TAP_12515 (  );
sky130_fd_sc_hd__tap_1 TAP_12516 (  );
sky130_fd_sc_hd__tap_1 TAP_12517 (  );
sky130_fd_sc_hd__tap_1 TAP_12518 (  );
sky130_fd_sc_hd__tap_1 TAP_12519 (  );
sky130_fd_sc_hd__tap_1 TAP_1252 (  );
sky130_fd_sc_hd__tap_1 TAP_12520 (  );
sky130_fd_sc_hd__tap_1 TAP_12521 (  );
sky130_fd_sc_hd__tap_1 TAP_12522 (  );
sky130_fd_sc_hd__tap_1 TAP_12523 (  );
sky130_fd_sc_hd__tap_1 TAP_12524 (  );
sky130_fd_sc_hd__tap_1 TAP_12525 (  );
sky130_fd_sc_hd__tap_1 TAP_12526 (  );
sky130_fd_sc_hd__tap_1 TAP_12527 (  );
sky130_fd_sc_hd__tap_1 TAP_12528 (  );
sky130_fd_sc_hd__tap_1 TAP_12529 (  );
sky130_fd_sc_hd__tap_1 TAP_1253 (  );
sky130_fd_sc_hd__tap_1 TAP_12530 (  );
sky130_fd_sc_hd__tap_1 TAP_12531 (  );
sky130_fd_sc_hd__tap_1 TAP_12532 (  );
sky130_fd_sc_hd__tap_1 TAP_12533 (  );
sky130_fd_sc_hd__tap_1 TAP_12534 (  );
sky130_fd_sc_hd__tap_1 TAP_12535 (  );
sky130_fd_sc_hd__tap_1 TAP_12536 (  );
sky130_fd_sc_hd__tap_1 TAP_12537 (  );
sky130_fd_sc_hd__tap_1 TAP_12538 (  );
sky130_fd_sc_hd__tap_1 TAP_12539 (  );
sky130_fd_sc_hd__tap_1 TAP_1254 (  );
sky130_fd_sc_hd__tap_1 TAP_12540 (  );
sky130_fd_sc_hd__tap_1 TAP_12541 (  );
sky130_fd_sc_hd__tap_1 TAP_12542 (  );
sky130_fd_sc_hd__tap_1 TAP_12543 (  );
sky130_fd_sc_hd__tap_1 TAP_12544 (  );
sky130_fd_sc_hd__tap_1 TAP_12545 (  );
sky130_fd_sc_hd__tap_1 TAP_12546 (  );
sky130_fd_sc_hd__tap_1 TAP_12547 (  );
sky130_fd_sc_hd__tap_1 TAP_12548 (  );
sky130_fd_sc_hd__tap_1 TAP_12549 (  );
sky130_fd_sc_hd__tap_1 TAP_1255 (  );
sky130_fd_sc_hd__tap_1 TAP_12550 (  );
sky130_fd_sc_hd__tap_1 TAP_12551 (  );
sky130_fd_sc_hd__tap_1 TAP_12552 (  );
sky130_fd_sc_hd__tap_1 TAP_12553 (  );
sky130_fd_sc_hd__tap_1 TAP_12554 (  );
sky130_fd_sc_hd__tap_1 TAP_12555 (  );
sky130_fd_sc_hd__tap_1 TAP_12556 (  );
sky130_fd_sc_hd__tap_1 TAP_12557 (  );
sky130_fd_sc_hd__tap_1 TAP_12558 (  );
sky130_fd_sc_hd__tap_1 TAP_12559 (  );
sky130_fd_sc_hd__tap_1 TAP_1256 (  );
sky130_fd_sc_hd__tap_1 TAP_12560 (  );
sky130_fd_sc_hd__tap_1 TAP_12561 (  );
sky130_fd_sc_hd__tap_1 TAP_12562 (  );
sky130_fd_sc_hd__tap_1 TAP_12563 (  );
sky130_fd_sc_hd__tap_1 TAP_12564 (  );
sky130_fd_sc_hd__tap_1 TAP_12565 (  );
sky130_fd_sc_hd__tap_1 TAP_12566 (  );
sky130_fd_sc_hd__tap_1 TAP_12567 (  );
sky130_fd_sc_hd__tap_1 TAP_12568 (  );
sky130_fd_sc_hd__tap_1 TAP_12569 (  );
sky130_fd_sc_hd__tap_1 TAP_1257 (  );
sky130_fd_sc_hd__tap_1 TAP_12570 (  );
sky130_fd_sc_hd__tap_1 TAP_12571 (  );
sky130_fd_sc_hd__tap_1 TAP_12572 (  );
sky130_fd_sc_hd__tap_1 TAP_12573 (  );
sky130_fd_sc_hd__tap_1 TAP_12574 (  );
sky130_fd_sc_hd__tap_1 TAP_12575 (  );
sky130_fd_sc_hd__tap_1 TAP_12576 (  );
sky130_fd_sc_hd__tap_1 TAP_12577 (  );
sky130_fd_sc_hd__tap_1 TAP_12578 (  );
sky130_fd_sc_hd__tap_1 TAP_12579 (  );
sky130_fd_sc_hd__tap_1 TAP_1258 (  );
sky130_fd_sc_hd__tap_1 TAP_12580 (  );
sky130_fd_sc_hd__tap_1 TAP_12581 (  );
sky130_fd_sc_hd__tap_1 TAP_12582 (  );
sky130_fd_sc_hd__tap_1 TAP_12583 (  );
sky130_fd_sc_hd__tap_1 TAP_12584 (  );
sky130_fd_sc_hd__tap_1 TAP_12585 (  );
sky130_fd_sc_hd__tap_1 TAP_12586 (  );
sky130_fd_sc_hd__tap_1 TAP_12587 (  );
sky130_fd_sc_hd__tap_1 TAP_12588 (  );
sky130_fd_sc_hd__tap_1 TAP_12589 (  );
sky130_fd_sc_hd__tap_1 TAP_1259 (  );
sky130_fd_sc_hd__tap_1 TAP_12590 (  );
sky130_fd_sc_hd__tap_1 TAP_12591 (  );
sky130_fd_sc_hd__tap_1 TAP_12592 (  );
sky130_fd_sc_hd__tap_1 TAP_12593 (  );
sky130_fd_sc_hd__tap_1 TAP_12594 (  );
sky130_fd_sc_hd__tap_1 TAP_12595 (  );
sky130_fd_sc_hd__tap_1 TAP_12596 (  );
sky130_fd_sc_hd__tap_1 TAP_12597 (  );
sky130_fd_sc_hd__tap_1 TAP_12598 (  );
sky130_fd_sc_hd__tap_1 TAP_12599 (  );
sky130_fd_sc_hd__tap_1 TAP_1260 (  );
sky130_fd_sc_hd__tap_1 TAP_12600 (  );
sky130_fd_sc_hd__tap_1 TAP_12601 (  );
sky130_fd_sc_hd__tap_1 TAP_12602 (  );
sky130_fd_sc_hd__tap_1 TAP_12603 (  );
sky130_fd_sc_hd__tap_1 TAP_12604 (  );
sky130_fd_sc_hd__tap_1 TAP_12605 (  );
sky130_fd_sc_hd__tap_1 TAP_12606 (  );
sky130_fd_sc_hd__tap_1 TAP_12607 (  );
sky130_fd_sc_hd__tap_1 TAP_12608 (  );
sky130_fd_sc_hd__tap_1 TAP_12609 (  );
sky130_fd_sc_hd__tap_1 TAP_1261 (  );
sky130_fd_sc_hd__tap_1 TAP_12610 (  );
sky130_fd_sc_hd__tap_1 TAP_12611 (  );
sky130_fd_sc_hd__tap_1 TAP_12612 (  );
sky130_fd_sc_hd__tap_1 TAP_12613 (  );
sky130_fd_sc_hd__tap_1 TAP_12614 (  );
sky130_fd_sc_hd__tap_1 TAP_12615 (  );
sky130_fd_sc_hd__tap_1 TAP_12616 (  );
sky130_fd_sc_hd__tap_1 TAP_12617 (  );
sky130_fd_sc_hd__tap_1 TAP_12618 (  );
sky130_fd_sc_hd__tap_1 TAP_12619 (  );
sky130_fd_sc_hd__tap_1 TAP_1262 (  );
sky130_fd_sc_hd__tap_1 TAP_12620 (  );
sky130_fd_sc_hd__tap_1 TAP_12621 (  );
sky130_fd_sc_hd__tap_1 TAP_12622 (  );
sky130_fd_sc_hd__tap_1 TAP_12623 (  );
sky130_fd_sc_hd__tap_1 TAP_12624 (  );
sky130_fd_sc_hd__tap_1 TAP_12625 (  );
sky130_fd_sc_hd__tap_1 TAP_12626 (  );
sky130_fd_sc_hd__tap_1 TAP_12627 (  );
sky130_fd_sc_hd__tap_1 TAP_12628 (  );
sky130_fd_sc_hd__tap_1 TAP_12629 (  );
sky130_fd_sc_hd__tap_1 TAP_1263 (  );
sky130_fd_sc_hd__tap_1 TAP_12630 (  );
sky130_fd_sc_hd__tap_1 TAP_12631 (  );
sky130_fd_sc_hd__tap_1 TAP_12632 (  );
sky130_fd_sc_hd__tap_1 TAP_12633 (  );
sky130_fd_sc_hd__tap_1 TAP_12634 (  );
sky130_fd_sc_hd__tap_1 TAP_12635 (  );
sky130_fd_sc_hd__tap_1 TAP_12636 (  );
sky130_fd_sc_hd__tap_1 TAP_12637 (  );
sky130_fd_sc_hd__tap_1 TAP_12638 (  );
sky130_fd_sc_hd__tap_1 TAP_12639 (  );
sky130_fd_sc_hd__tap_1 TAP_1264 (  );
sky130_fd_sc_hd__tap_1 TAP_12640 (  );
sky130_fd_sc_hd__tap_1 TAP_12641 (  );
sky130_fd_sc_hd__tap_1 TAP_12642 (  );
sky130_fd_sc_hd__tap_1 TAP_12643 (  );
sky130_fd_sc_hd__tap_1 TAP_12644 (  );
sky130_fd_sc_hd__tap_1 TAP_12645 (  );
sky130_fd_sc_hd__tap_1 TAP_12646 (  );
sky130_fd_sc_hd__tap_1 TAP_12647 (  );
sky130_fd_sc_hd__tap_1 TAP_12648 (  );
sky130_fd_sc_hd__tap_1 TAP_12649 (  );
sky130_fd_sc_hd__tap_1 TAP_1265 (  );
sky130_fd_sc_hd__tap_1 TAP_12650 (  );
sky130_fd_sc_hd__tap_1 TAP_12651 (  );
sky130_fd_sc_hd__tap_1 TAP_12652 (  );
sky130_fd_sc_hd__tap_1 TAP_12653 (  );
sky130_fd_sc_hd__tap_1 TAP_12654 (  );
sky130_fd_sc_hd__tap_1 TAP_12655 (  );
sky130_fd_sc_hd__tap_1 TAP_12656 (  );
sky130_fd_sc_hd__tap_1 TAP_12657 (  );
sky130_fd_sc_hd__tap_1 TAP_12658 (  );
sky130_fd_sc_hd__tap_1 TAP_12659 (  );
sky130_fd_sc_hd__tap_1 TAP_1266 (  );
sky130_fd_sc_hd__tap_1 TAP_12660 (  );
sky130_fd_sc_hd__tap_1 TAP_12661 (  );
sky130_fd_sc_hd__tap_1 TAP_12662 (  );
sky130_fd_sc_hd__tap_1 TAP_12663 (  );
sky130_fd_sc_hd__tap_1 TAP_12664 (  );
sky130_fd_sc_hd__tap_1 TAP_12665 (  );
sky130_fd_sc_hd__tap_1 TAP_12666 (  );
sky130_fd_sc_hd__tap_1 TAP_12667 (  );
sky130_fd_sc_hd__tap_1 TAP_12668 (  );
sky130_fd_sc_hd__tap_1 TAP_12669 (  );
sky130_fd_sc_hd__tap_1 TAP_1267 (  );
sky130_fd_sc_hd__tap_1 TAP_12670 (  );
sky130_fd_sc_hd__tap_1 TAP_12671 (  );
sky130_fd_sc_hd__tap_1 TAP_12672 (  );
sky130_fd_sc_hd__tap_1 TAP_12673 (  );
sky130_fd_sc_hd__tap_1 TAP_12674 (  );
sky130_fd_sc_hd__tap_1 TAP_12675 (  );
sky130_fd_sc_hd__tap_1 TAP_12676 (  );
sky130_fd_sc_hd__tap_1 TAP_12677 (  );
sky130_fd_sc_hd__tap_1 TAP_12678 (  );
sky130_fd_sc_hd__tap_1 TAP_12679 (  );
sky130_fd_sc_hd__tap_1 TAP_1268 (  );
sky130_fd_sc_hd__tap_1 TAP_12680 (  );
sky130_fd_sc_hd__tap_1 TAP_12681 (  );
sky130_fd_sc_hd__tap_1 TAP_12682 (  );
sky130_fd_sc_hd__tap_1 TAP_12683 (  );
sky130_fd_sc_hd__tap_1 TAP_12684 (  );
sky130_fd_sc_hd__tap_1 TAP_12685 (  );
sky130_fd_sc_hd__tap_1 TAP_12686 (  );
sky130_fd_sc_hd__tap_1 TAP_12687 (  );
sky130_fd_sc_hd__tap_1 TAP_12688 (  );
sky130_fd_sc_hd__tap_1 TAP_12689 (  );
sky130_fd_sc_hd__tap_1 TAP_1269 (  );
sky130_fd_sc_hd__tap_1 TAP_12690 (  );
sky130_fd_sc_hd__tap_1 TAP_12691 (  );
sky130_fd_sc_hd__tap_1 TAP_12692 (  );
sky130_fd_sc_hd__tap_1 TAP_12693 (  );
sky130_fd_sc_hd__tap_1 TAP_12694 (  );
sky130_fd_sc_hd__tap_1 TAP_12695 (  );
sky130_fd_sc_hd__tap_1 TAP_12696 (  );
sky130_fd_sc_hd__tap_1 TAP_12697 (  );
sky130_fd_sc_hd__tap_1 TAP_12698 (  );
sky130_fd_sc_hd__tap_1 TAP_12699 (  );
sky130_fd_sc_hd__tap_1 TAP_1270 (  );
sky130_fd_sc_hd__tap_1 TAP_12700 (  );
sky130_fd_sc_hd__tap_1 TAP_12701 (  );
sky130_fd_sc_hd__tap_1 TAP_12702 (  );
sky130_fd_sc_hd__tap_1 TAP_12703 (  );
sky130_fd_sc_hd__tap_1 TAP_12704 (  );
sky130_fd_sc_hd__tap_1 TAP_12705 (  );
sky130_fd_sc_hd__tap_1 TAP_12706 (  );
sky130_fd_sc_hd__tap_1 TAP_12707 (  );
sky130_fd_sc_hd__tap_1 TAP_12708 (  );
sky130_fd_sc_hd__tap_1 TAP_12709 (  );
sky130_fd_sc_hd__tap_1 TAP_1271 (  );
sky130_fd_sc_hd__tap_1 TAP_12710 (  );
sky130_fd_sc_hd__tap_1 TAP_12711 (  );
sky130_fd_sc_hd__tap_1 TAP_12712 (  );
sky130_fd_sc_hd__tap_1 TAP_12713 (  );
sky130_fd_sc_hd__tap_1 TAP_12714 (  );
sky130_fd_sc_hd__tap_1 TAP_12715 (  );
sky130_fd_sc_hd__tap_1 TAP_12716 (  );
sky130_fd_sc_hd__tap_1 TAP_12717 (  );
sky130_fd_sc_hd__tap_1 TAP_12718 (  );
sky130_fd_sc_hd__tap_1 TAP_12719 (  );
sky130_fd_sc_hd__tap_1 TAP_1272 (  );
sky130_fd_sc_hd__tap_1 TAP_12720 (  );
sky130_fd_sc_hd__tap_1 TAP_12721 (  );
sky130_fd_sc_hd__tap_1 TAP_12722 (  );
sky130_fd_sc_hd__tap_1 TAP_12723 (  );
sky130_fd_sc_hd__tap_1 TAP_12724 (  );
sky130_fd_sc_hd__tap_1 TAP_12725 (  );
sky130_fd_sc_hd__tap_1 TAP_12726 (  );
sky130_fd_sc_hd__tap_1 TAP_12727 (  );
sky130_fd_sc_hd__tap_1 TAP_12728 (  );
sky130_fd_sc_hd__tap_1 TAP_12729 (  );
sky130_fd_sc_hd__tap_1 TAP_1273 (  );
sky130_fd_sc_hd__tap_1 TAP_12730 (  );
sky130_fd_sc_hd__tap_1 TAP_12731 (  );
sky130_fd_sc_hd__tap_1 TAP_12732 (  );
sky130_fd_sc_hd__tap_1 TAP_12733 (  );
sky130_fd_sc_hd__tap_1 TAP_12734 (  );
sky130_fd_sc_hd__tap_1 TAP_12735 (  );
sky130_fd_sc_hd__tap_1 TAP_12736 (  );
sky130_fd_sc_hd__tap_1 TAP_12737 (  );
sky130_fd_sc_hd__tap_1 TAP_12738 (  );
sky130_fd_sc_hd__tap_1 TAP_12739 (  );
sky130_fd_sc_hd__tap_1 TAP_1274 (  );
sky130_fd_sc_hd__tap_1 TAP_12740 (  );
sky130_fd_sc_hd__tap_1 TAP_12741 (  );
sky130_fd_sc_hd__tap_1 TAP_12742 (  );
sky130_fd_sc_hd__tap_1 TAP_12743 (  );
sky130_fd_sc_hd__tap_1 TAP_12744 (  );
sky130_fd_sc_hd__tap_1 TAP_12745 (  );
sky130_fd_sc_hd__tap_1 TAP_12746 (  );
sky130_fd_sc_hd__tap_1 TAP_12747 (  );
sky130_fd_sc_hd__tap_1 TAP_12748 (  );
sky130_fd_sc_hd__tap_1 TAP_12749 (  );
sky130_fd_sc_hd__tap_1 TAP_1275 (  );
sky130_fd_sc_hd__tap_1 TAP_12750 (  );
sky130_fd_sc_hd__tap_1 TAP_12751 (  );
sky130_fd_sc_hd__tap_1 TAP_12752 (  );
sky130_fd_sc_hd__tap_1 TAP_12753 (  );
sky130_fd_sc_hd__tap_1 TAP_12754 (  );
sky130_fd_sc_hd__tap_1 TAP_12755 (  );
sky130_fd_sc_hd__tap_1 TAP_12756 (  );
sky130_fd_sc_hd__tap_1 TAP_12757 (  );
sky130_fd_sc_hd__tap_1 TAP_12758 (  );
sky130_fd_sc_hd__tap_1 TAP_12759 (  );
sky130_fd_sc_hd__tap_1 TAP_1276 (  );
sky130_fd_sc_hd__tap_1 TAP_12760 (  );
sky130_fd_sc_hd__tap_1 TAP_12761 (  );
sky130_fd_sc_hd__tap_1 TAP_12762 (  );
sky130_fd_sc_hd__tap_1 TAP_12763 (  );
sky130_fd_sc_hd__tap_1 TAP_12764 (  );
sky130_fd_sc_hd__tap_1 TAP_12765 (  );
sky130_fd_sc_hd__tap_1 TAP_12766 (  );
sky130_fd_sc_hd__tap_1 TAP_12767 (  );
sky130_fd_sc_hd__tap_1 TAP_12768 (  );
sky130_fd_sc_hd__tap_1 TAP_12769 (  );
sky130_fd_sc_hd__tap_1 TAP_1277 (  );
sky130_fd_sc_hd__tap_1 TAP_12770 (  );
sky130_fd_sc_hd__tap_1 TAP_12771 (  );
sky130_fd_sc_hd__tap_1 TAP_12772 (  );
sky130_fd_sc_hd__tap_1 TAP_12773 (  );
sky130_fd_sc_hd__tap_1 TAP_12774 (  );
sky130_fd_sc_hd__tap_1 TAP_12775 (  );
sky130_fd_sc_hd__tap_1 TAP_12776 (  );
sky130_fd_sc_hd__tap_1 TAP_12777 (  );
sky130_fd_sc_hd__tap_1 TAP_12778 (  );
sky130_fd_sc_hd__tap_1 TAP_12779 (  );
sky130_fd_sc_hd__tap_1 TAP_1278 (  );
sky130_fd_sc_hd__tap_1 TAP_12780 (  );
sky130_fd_sc_hd__tap_1 TAP_12781 (  );
sky130_fd_sc_hd__tap_1 TAP_12782 (  );
sky130_fd_sc_hd__tap_1 TAP_12783 (  );
sky130_fd_sc_hd__tap_1 TAP_12784 (  );
sky130_fd_sc_hd__tap_1 TAP_12785 (  );
sky130_fd_sc_hd__tap_1 TAP_12786 (  );
sky130_fd_sc_hd__tap_1 TAP_12787 (  );
sky130_fd_sc_hd__tap_1 TAP_12788 (  );
sky130_fd_sc_hd__tap_1 TAP_12789 (  );
sky130_fd_sc_hd__tap_1 TAP_1279 (  );
sky130_fd_sc_hd__tap_1 TAP_12790 (  );
sky130_fd_sc_hd__tap_1 TAP_12791 (  );
sky130_fd_sc_hd__tap_1 TAP_12792 (  );
sky130_fd_sc_hd__tap_1 TAP_12793 (  );
sky130_fd_sc_hd__tap_1 TAP_12794 (  );
sky130_fd_sc_hd__tap_1 TAP_12795 (  );
sky130_fd_sc_hd__tap_1 TAP_12796 (  );
sky130_fd_sc_hd__tap_1 TAP_12797 (  );
sky130_fd_sc_hd__tap_1 TAP_12798 (  );
sky130_fd_sc_hd__tap_1 TAP_12799 (  );
sky130_fd_sc_hd__tap_1 TAP_1280 (  );
sky130_fd_sc_hd__tap_1 TAP_12800 (  );
sky130_fd_sc_hd__tap_1 TAP_12801 (  );
sky130_fd_sc_hd__tap_1 TAP_12802 (  );
sky130_fd_sc_hd__tap_1 TAP_12803 (  );
sky130_fd_sc_hd__tap_1 TAP_12804 (  );
sky130_fd_sc_hd__tap_1 TAP_12805 (  );
sky130_fd_sc_hd__tap_1 TAP_12806 (  );
sky130_fd_sc_hd__tap_1 TAP_12807 (  );
sky130_fd_sc_hd__tap_1 TAP_12808 (  );
sky130_fd_sc_hd__tap_1 TAP_12809 (  );
sky130_fd_sc_hd__tap_1 TAP_1281 (  );
sky130_fd_sc_hd__tap_1 TAP_12810 (  );
sky130_fd_sc_hd__tap_1 TAP_12811 (  );
sky130_fd_sc_hd__tap_1 TAP_12812 (  );
sky130_fd_sc_hd__tap_1 TAP_12813 (  );
sky130_fd_sc_hd__tap_1 TAP_12814 (  );
sky130_fd_sc_hd__tap_1 TAP_12815 (  );
sky130_fd_sc_hd__tap_1 TAP_12816 (  );
sky130_fd_sc_hd__tap_1 TAP_12817 (  );
sky130_fd_sc_hd__tap_1 TAP_12818 (  );
sky130_fd_sc_hd__tap_1 TAP_12819 (  );
sky130_fd_sc_hd__tap_1 TAP_1282 (  );
sky130_fd_sc_hd__tap_1 TAP_12820 (  );
sky130_fd_sc_hd__tap_1 TAP_12821 (  );
sky130_fd_sc_hd__tap_1 TAP_12822 (  );
sky130_fd_sc_hd__tap_1 TAP_12823 (  );
sky130_fd_sc_hd__tap_1 TAP_12824 (  );
sky130_fd_sc_hd__tap_1 TAP_12825 (  );
sky130_fd_sc_hd__tap_1 TAP_12826 (  );
sky130_fd_sc_hd__tap_1 TAP_12827 (  );
sky130_fd_sc_hd__tap_1 TAP_12828 (  );
sky130_fd_sc_hd__tap_1 TAP_12829 (  );
sky130_fd_sc_hd__tap_1 TAP_1283 (  );
sky130_fd_sc_hd__tap_1 TAP_12830 (  );
sky130_fd_sc_hd__tap_1 TAP_12831 (  );
sky130_fd_sc_hd__tap_1 TAP_12832 (  );
sky130_fd_sc_hd__tap_1 TAP_12833 (  );
sky130_fd_sc_hd__tap_1 TAP_12834 (  );
sky130_fd_sc_hd__tap_1 TAP_12835 (  );
sky130_fd_sc_hd__tap_1 TAP_12836 (  );
sky130_fd_sc_hd__tap_1 TAP_12837 (  );
sky130_fd_sc_hd__tap_1 TAP_12838 (  );
sky130_fd_sc_hd__tap_1 TAP_12839 (  );
sky130_fd_sc_hd__tap_1 TAP_1284 (  );
sky130_fd_sc_hd__tap_1 TAP_12840 (  );
sky130_fd_sc_hd__tap_1 TAP_12841 (  );
sky130_fd_sc_hd__tap_1 TAP_12842 (  );
sky130_fd_sc_hd__tap_1 TAP_12843 (  );
sky130_fd_sc_hd__tap_1 TAP_12844 (  );
sky130_fd_sc_hd__tap_1 TAP_12845 (  );
sky130_fd_sc_hd__tap_1 TAP_12846 (  );
sky130_fd_sc_hd__tap_1 TAP_12847 (  );
sky130_fd_sc_hd__tap_1 TAP_12848 (  );
sky130_fd_sc_hd__tap_1 TAP_12849 (  );
sky130_fd_sc_hd__tap_1 TAP_1285 (  );
sky130_fd_sc_hd__tap_1 TAP_12850 (  );
sky130_fd_sc_hd__tap_1 TAP_12851 (  );
sky130_fd_sc_hd__tap_1 TAP_12852 (  );
sky130_fd_sc_hd__tap_1 TAP_12853 (  );
sky130_fd_sc_hd__tap_1 TAP_12854 (  );
sky130_fd_sc_hd__tap_1 TAP_12855 (  );
sky130_fd_sc_hd__tap_1 TAP_12856 (  );
sky130_fd_sc_hd__tap_1 TAP_12857 (  );
sky130_fd_sc_hd__tap_1 TAP_12858 (  );
sky130_fd_sc_hd__tap_1 TAP_12859 (  );
sky130_fd_sc_hd__tap_1 TAP_1286 (  );
sky130_fd_sc_hd__tap_1 TAP_12860 (  );
sky130_fd_sc_hd__tap_1 TAP_12861 (  );
sky130_fd_sc_hd__tap_1 TAP_12862 (  );
sky130_fd_sc_hd__tap_1 TAP_12863 (  );
sky130_fd_sc_hd__tap_1 TAP_12864 (  );
sky130_fd_sc_hd__tap_1 TAP_12865 (  );
sky130_fd_sc_hd__tap_1 TAP_12866 (  );
sky130_fd_sc_hd__tap_1 TAP_12867 (  );
sky130_fd_sc_hd__tap_1 TAP_12868 (  );
sky130_fd_sc_hd__tap_1 TAP_12869 (  );
sky130_fd_sc_hd__tap_1 TAP_1287 (  );
sky130_fd_sc_hd__tap_1 TAP_12870 (  );
sky130_fd_sc_hd__tap_1 TAP_12871 (  );
sky130_fd_sc_hd__tap_1 TAP_12872 (  );
sky130_fd_sc_hd__tap_1 TAP_12873 (  );
sky130_fd_sc_hd__tap_1 TAP_12874 (  );
sky130_fd_sc_hd__tap_1 TAP_12875 (  );
sky130_fd_sc_hd__tap_1 TAP_12876 (  );
sky130_fd_sc_hd__tap_1 TAP_12877 (  );
sky130_fd_sc_hd__tap_1 TAP_12878 (  );
sky130_fd_sc_hd__tap_1 TAP_12879 (  );
sky130_fd_sc_hd__tap_1 TAP_1288 (  );
sky130_fd_sc_hd__tap_1 TAP_12880 (  );
sky130_fd_sc_hd__tap_1 TAP_12881 (  );
sky130_fd_sc_hd__tap_1 TAP_12882 (  );
sky130_fd_sc_hd__tap_1 TAP_12883 (  );
sky130_fd_sc_hd__tap_1 TAP_12884 (  );
sky130_fd_sc_hd__tap_1 TAP_12885 (  );
sky130_fd_sc_hd__tap_1 TAP_12886 (  );
sky130_fd_sc_hd__tap_1 TAP_12887 (  );
sky130_fd_sc_hd__tap_1 TAP_12888 (  );
sky130_fd_sc_hd__tap_1 TAP_12889 (  );
sky130_fd_sc_hd__tap_1 TAP_1289 (  );
sky130_fd_sc_hd__tap_1 TAP_12890 (  );
sky130_fd_sc_hd__tap_1 TAP_12891 (  );
sky130_fd_sc_hd__tap_1 TAP_12892 (  );
sky130_fd_sc_hd__tap_1 TAP_12893 (  );
sky130_fd_sc_hd__tap_1 TAP_12894 (  );
sky130_fd_sc_hd__tap_1 TAP_12895 (  );
sky130_fd_sc_hd__tap_1 TAP_12896 (  );
sky130_fd_sc_hd__tap_1 TAP_12897 (  );
sky130_fd_sc_hd__tap_1 TAP_12898 (  );
sky130_fd_sc_hd__tap_1 TAP_12899 (  );
sky130_fd_sc_hd__tap_1 TAP_1290 (  );
sky130_fd_sc_hd__tap_1 TAP_12900 (  );
sky130_fd_sc_hd__tap_1 TAP_12901 (  );
sky130_fd_sc_hd__tap_1 TAP_12902 (  );
sky130_fd_sc_hd__tap_1 TAP_12903 (  );
sky130_fd_sc_hd__tap_1 TAP_12904 (  );
sky130_fd_sc_hd__tap_1 TAP_12905 (  );
sky130_fd_sc_hd__tap_1 TAP_12906 (  );
sky130_fd_sc_hd__tap_1 TAP_12907 (  );
sky130_fd_sc_hd__tap_1 TAP_12908 (  );
sky130_fd_sc_hd__tap_1 TAP_12909 (  );
sky130_fd_sc_hd__tap_1 TAP_1291 (  );
sky130_fd_sc_hd__tap_1 TAP_12910 (  );
sky130_fd_sc_hd__tap_1 TAP_12911 (  );
sky130_fd_sc_hd__tap_1 TAP_12912 (  );
sky130_fd_sc_hd__tap_1 TAP_12913 (  );
sky130_fd_sc_hd__tap_1 TAP_12914 (  );
sky130_fd_sc_hd__tap_1 TAP_12915 (  );
sky130_fd_sc_hd__tap_1 TAP_12916 (  );
sky130_fd_sc_hd__tap_1 TAP_12917 (  );
sky130_fd_sc_hd__tap_1 TAP_12918 (  );
sky130_fd_sc_hd__tap_1 TAP_12919 (  );
sky130_fd_sc_hd__tap_1 TAP_1292 (  );
sky130_fd_sc_hd__tap_1 TAP_12920 (  );
sky130_fd_sc_hd__tap_1 TAP_12921 (  );
sky130_fd_sc_hd__tap_1 TAP_12922 (  );
sky130_fd_sc_hd__tap_1 TAP_12923 (  );
sky130_fd_sc_hd__tap_1 TAP_12924 (  );
sky130_fd_sc_hd__tap_1 TAP_12925 (  );
sky130_fd_sc_hd__tap_1 TAP_12926 (  );
sky130_fd_sc_hd__tap_1 TAP_12927 (  );
sky130_fd_sc_hd__tap_1 TAP_12928 (  );
sky130_fd_sc_hd__tap_1 TAP_12929 (  );
sky130_fd_sc_hd__tap_1 TAP_1293 (  );
sky130_fd_sc_hd__tap_1 TAP_12930 (  );
sky130_fd_sc_hd__tap_1 TAP_12931 (  );
sky130_fd_sc_hd__tap_1 TAP_12932 (  );
sky130_fd_sc_hd__tap_1 TAP_12933 (  );
sky130_fd_sc_hd__tap_1 TAP_12934 (  );
sky130_fd_sc_hd__tap_1 TAP_12935 (  );
sky130_fd_sc_hd__tap_1 TAP_12936 (  );
sky130_fd_sc_hd__tap_1 TAP_12937 (  );
sky130_fd_sc_hd__tap_1 TAP_12938 (  );
sky130_fd_sc_hd__tap_1 TAP_12939 (  );
sky130_fd_sc_hd__tap_1 TAP_1294 (  );
sky130_fd_sc_hd__tap_1 TAP_12940 (  );
sky130_fd_sc_hd__tap_1 TAP_12941 (  );
sky130_fd_sc_hd__tap_1 TAP_12942 (  );
sky130_fd_sc_hd__tap_1 TAP_12943 (  );
sky130_fd_sc_hd__tap_1 TAP_12944 (  );
sky130_fd_sc_hd__tap_1 TAP_12945 (  );
sky130_fd_sc_hd__tap_1 TAP_12946 (  );
sky130_fd_sc_hd__tap_1 TAP_12947 (  );
sky130_fd_sc_hd__tap_1 TAP_12948 (  );
sky130_fd_sc_hd__tap_1 TAP_12949 (  );
sky130_fd_sc_hd__tap_1 TAP_1295 (  );
sky130_fd_sc_hd__tap_1 TAP_12950 (  );
sky130_fd_sc_hd__tap_1 TAP_12951 (  );
sky130_fd_sc_hd__tap_1 TAP_12952 (  );
sky130_fd_sc_hd__tap_1 TAP_12953 (  );
sky130_fd_sc_hd__tap_1 TAP_12954 (  );
sky130_fd_sc_hd__tap_1 TAP_12955 (  );
sky130_fd_sc_hd__tap_1 TAP_12956 (  );
sky130_fd_sc_hd__tap_1 TAP_12957 (  );
sky130_fd_sc_hd__tap_1 TAP_12958 (  );
sky130_fd_sc_hd__tap_1 TAP_12959 (  );
sky130_fd_sc_hd__tap_1 TAP_1296 (  );
sky130_fd_sc_hd__tap_1 TAP_12960 (  );
sky130_fd_sc_hd__tap_1 TAP_12961 (  );
sky130_fd_sc_hd__tap_1 TAP_12962 (  );
sky130_fd_sc_hd__tap_1 TAP_12963 (  );
sky130_fd_sc_hd__tap_1 TAP_12964 (  );
sky130_fd_sc_hd__tap_1 TAP_12965 (  );
sky130_fd_sc_hd__tap_1 TAP_12966 (  );
sky130_fd_sc_hd__tap_1 TAP_12967 (  );
sky130_fd_sc_hd__tap_1 TAP_12968 (  );
sky130_fd_sc_hd__tap_1 TAP_12969 (  );
sky130_fd_sc_hd__tap_1 TAP_1297 (  );
sky130_fd_sc_hd__tap_1 TAP_12970 (  );
sky130_fd_sc_hd__tap_1 TAP_12971 (  );
sky130_fd_sc_hd__tap_1 TAP_12972 (  );
sky130_fd_sc_hd__tap_1 TAP_12973 (  );
sky130_fd_sc_hd__tap_1 TAP_12974 (  );
sky130_fd_sc_hd__tap_1 TAP_12975 (  );
sky130_fd_sc_hd__tap_1 TAP_12976 (  );
sky130_fd_sc_hd__tap_1 TAP_12977 (  );
sky130_fd_sc_hd__tap_1 TAP_12978 (  );
sky130_fd_sc_hd__tap_1 TAP_12979 (  );
sky130_fd_sc_hd__tap_1 TAP_1298 (  );
sky130_fd_sc_hd__tap_1 TAP_12980 (  );
sky130_fd_sc_hd__tap_1 TAP_12981 (  );
sky130_fd_sc_hd__tap_1 TAP_12982 (  );
sky130_fd_sc_hd__tap_1 TAP_12983 (  );
sky130_fd_sc_hd__tap_1 TAP_12984 (  );
sky130_fd_sc_hd__tap_1 TAP_12985 (  );
sky130_fd_sc_hd__tap_1 TAP_12986 (  );
sky130_fd_sc_hd__tap_1 TAP_12987 (  );
sky130_fd_sc_hd__tap_1 TAP_12988 (  );
sky130_fd_sc_hd__tap_1 TAP_12989 (  );
sky130_fd_sc_hd__tap_1 TAP_1299 (  );
sky130_fd_sc_hd__tap_1 TAP_12990 (  );
sky130_fd_sc_hd__tap_1 TAP_12991 (  );
sky130_fd_sc_hd__tap_1 TAP_12992 (  );
sky130_fd_sc_hd__tap_1 TAP_12993 (  );
sky130_fd_sc_hd__tap_1 TAP_12994 (  );
sky130_fd_sc_hd__tap_1 TAP_12995 (  );
sky130_fd_sc_hd__tap_1 TAP_12996 (  );
sky130_fd_sc_hd__tap_1 TAP_12997 (  );
sky130_fd_sc_hd__tap_1 TAP_12998 (  );
sky130_fd_sc_hd__tap_1 TAP_12999 (  );
sky130_fd_sc_hd__tap_1 TAP_1300 (  );
sky130_fd_sc_hd__tap_1 TAP_13000 (  );
sky130_fd_sc_hd__tap_1 TAP_13001 (  );
sky130_fd_sc_hd__tap_1 TAP_13002 (  );
sky130_fd_sc_hd__tap_1 TAP_13003 (  );
sky130_fd_sc_hd__tap_1 TAP_13004 (  );
sky130_fd_sc_hd__tap_1 TAP_13005 (  );
sky130_fd_sc_hd__tap_1 TAP_13006 (  );
sky130_fd_sc_hd__tap_1 TAP_13007 (  );
sky130_fd_sc_hd__tap_1 TAP_13008 (  );
sky130_fd_sc_hd__tap_1 TAP_13009 (  );
sky130_fd_sc_hd__tap_1 TAP_1301 (  );
sky130_fd_sc_hd__tap_1 TAP_13010 (  );
sky130_fd_sc_hd__tap_1 TAP_13011 (  );
sky130_fd_sc_hd__tap_1 TAP_13012 (  );
sky130_fd_sc_hd__tap_1 TAP_13013 (  );
sky130_fd_sc_hd__tap_1 TAP_13014 (  );
sky130_fd_sc_hd__tap_1 TAP_13015 (  );
sky130_fd_sc_hd__tap_1 TAP_13016 (  );
sky130_fd_sc_hd__tap_1 TAP_13017 (  );
sky130_fd_sc_hd__tap_1 TAP_13018 (  );
sky130_fd_sc_hd__tap_1 TAP_13019 (  );
sky130_fd_sc_hd__tap_1 TAP_1302 (  );
sky130_fd_sc_hd__tap_1 TAP_13020 (  );
sky130_fd_sc_hd__tap_1 TAP_13021 (  );
sky130_fd_sc_hd__tap_1 TAP_13022 (  );
sky130_fd_sc_hd__tap_1 TAP_13023 (  );
sky130_fd_sc_hd__tap_1 TAP_13024 (  );
sky130_fd_sc_hd__tap_1 TAP_13025 (  );
sky130_fd_sc_hd__tap_1 TAP_13026 (  );
sky130_fd_sc_hd__tap_1 TAP_13027 (  );
sky130_fd_sc_hd__tap_1 TAP_13028 (  );
sky130_fd_sc_hd__tap_1 TAP_13029 (  );
sky130_fd_sc_hd__tap_1 TAP_1303 (  );
sky130_fd_sc_hd__tap_1 TAP_13030 (  );
sky130_fd_sc_hd__tap_1 TAP_13031 (  );
sky130_fd_sc_hd__tap_1 TAP_13032 (  );
sky130_fd_sc_hd__tap_1 TAP_13033 (  );
sky130_fd_sc_hd__tap_1 TAP_13034 (  );
sky130_fd_sc_hd__tap_1 TAP_13035 (  );
sky130_fd_sc_hd__tap_1 TAP_13036 (  );
sky130_fd_sc_hd__tap_1 TAP_13037 (  );
sky130_fd_sc_hd__tap_1 TAP_13038 (  );
sky130_fd_sc_hd__tap_1 TAP_13039 (  );
sky130_fd_sc_hd__tap_1 TAP_1304 (  );
sky130_fd_sc_hd__tap_1 TAP_13040 (  );
sky130_fd_sc_hd__tap_1 TAP_13041 (  );
sky130_fd_sc_hd__tap_1 TAP_13042 (  );
sky130_fd_sc_hd__tap_1 TAP_13043 (  );
sky130_fd_sc_hd__tap_1 TAP_13044 (  );
sky130_fd_sc_hd__tap_1 TAP_13045 (  );
sky130_fd_sc_hd__tap_1 TAP_13046 (  );
sky130_fd_sc_hd__tap_1 TAP_13047 (  );
sky130_fd_sc_hd__tap_1 TAP_13048 (  );
sky130_fd_sc_hd__tap_1 TAP_13049 (  );
sky130_fd_sc_hd__tap_1 TAP_1305 (  );
sky130_fd_sc_hd__tap_1 TAP_13050 (  );
sky130_fd_sc_hd__tap_1 TAP_13051 (  );
sky130_fd_sc_hd__tap_1 TAP_13052 (  );
sky130_fd_sc_hd__tap_1 TAP_13053 (  );
sky130_fd_sc_hd__tap_1 TAP_13054 (  );
sky130_fd_sc_hd__tap_1 TAP_13055 (  );
sky130_fd_sc_hd__tap_1 TAP_13056 (  );
sky130_fd_sc_hd__tap_1 TAP_13057 (  );
sky130_fd_sc_hd__tap_1 TAP_13058 (  );
sky130_fd_sc_hd__tap_1 TAP_13059 (  );
sky130_fd_sc_hd__tap_1 TAP_1306 (  );
sky130_fd_sc_hd__tap_1 TAP_13060 (  );
sky130_fd_sc_hd__tap_1 TAP_13061 (  );
sky130_fd_sc_hd__tap_1 TAP_13062 (  );
sky130_fd_sc_hd__tap_1 TAP_13063 (  );
sky130_fd_sc_hd__tap_1 TAP_13064 (  );
sky130_fd_sc_hd__tap_1 TAP_13065 (  );
sky130_fd_sc_hd__tap_1 TAP_13066 (  );
sky130_fd_sc_hd__tap_1 TAP_13067 (  );
sky130_fd_sc_hd__tap_1 TAP_13068 (  );
sky130_fd_sc_hd__tap_1 TAP_13069 (  );
sky130_fd_sc_hd__tap_1 TAP_1307 (  );
sky130_fd_sc_hd__tap_1 TAP_13070 (  );
sky130_fd_sc_hd__tap_1 TAP_13071 (  );
sky130_fd_sc_hd__tap_1 TAP_13072 (  );
sky130_fd_sc_hd__tap_1 TAP_13073 (  );
sky130_fd_sc_hd__tap_1 TAP_13074 (  );
sky130_fd_sc_hd__tap_1 TAP_13075 (  );
sky130_fd_sc_hd__tap_1 TAP_13076 (  );
sky130_fd_sc_hd__tap_1 TAP_13077 (  );
sky130_fd_sc_hd__tap_1 TAP_13078 (  );
sky130_fd_sc_hd__tap_1 TAP_13079 (  );
sky130_fd_sc_hd__tap_1 TAP_1308 (  );
sky130_fd_sc_hd__tap_1 TAP_13080 (  );
sky130_fd_sc_hd__tap_1 TAP_13081 (  );
sky130_fd_sc_hd__tap_1 TAP_13082 (  );
sky130_fd_sc_hd__tap_1 TAP_13083 (  );
sky130_fd_sc_hd__tap_1 TAP_13084 (  );
sky130_fd_sc_hd__tap_1 TAP_13085 (  );
sky130_fd_sc_hd__tap_1 TAP_13086 (  );
sky130_fd_sc_hd__tap_1 TAP_13087 (  );
sky130_fd_sc_hd__tap_1 TAP_13088 (  );
sky130_fd_sc_hd__tap_1 TAP_13089 (  );
sky130_fd_sc_hd__tap_1 TAP_1309 (  );
sky130_fd_sc_hd__tap_1 TAP_13090 (  );
sky130_fd_sc_hd__tap_1 TAP_13091 (  );
sky130_fd_sc_hd__tap_1 TAP_13092 (  );
sky130_fd_sc_hd__tap_1 TAP_13093 (  );
sky130_fd_sc_hd__tap_1 TAP_13094 (  );
sky130_fd_sc_hd__tap_1 TAP_13095 (  );
sky130_fd_sc_hd__tap_1 TAP_13096 (  );
sky130_fd_sc_hd__tap_1 TAP_13097 (  );
sky130_fd_sc_hd__tap_1 TAP_13098 (  );
sky130_fd_sc_hd__tap_1 TAP_13099 (  );
sky130_fd_sc_hd__tap_1 TAP_1310 (  );
sky130_fd_sc_hd__tap_1 TAP_13100 (  );
sky130_fd_sc_hd__tap_1 TAP_13101 (  );
sky130_fd_sc_hd__tap_1 TAP_13102 (  );
sky130_fd_sc_hd__tap_1 TAP_13103 (  );
sky130_fd_sc_hd__tap_1 TAP_13104 (  );
sky130_fd_sc_hd__tap_1 TAP_13105 (  );
sky130_fd_sc_hd__tap_1 TAP_13106 (  );
sky130_fd_sc_hd__tap_1 TAP_13107 (  );
sky130_fd_sc_hd__tap_1 TAP_13108 (  );
sky130_fd_sc_hd__tap_1 TAP_13109 (  );
sky130_fd_sc_hd__tap_1 TAP_1311 (  );
sky130_fd_sc_hd__tap_1 TAP_13110 (  );
sky130_fd_sc_hd__tap_1 TAP_13111 (  );
sky130_fd_sc_hd__tap_1 TAP_13112 (  );
sky130_fd_sc_hd__tap_1 TAP_13113 (  );
sky130_fd_sc_hd__tap_1 TAP_13114 (  );
sky130_fd_sc_hd__tap_1 TAP_13115 (  );
sky130_fd_sc_hd__tap_1 TAP_13116 (  );
sky130_fd_sc_hd__tap_1 TAP_13117 (  );
sky130_fd_sc_hd__tap_1 TAP_13118 (  );
sky130_fd_sc_hd__tap_1 TAP_13119 (  );
sky130_fd_sc_hd__tap_1 TAP_1312 (  );
sky130_fd_sc_hd__tap_1 TAP_13120 (  );
sky130_fd_sc_hd__tap_1 TAP_13121 (  );
sky130_fd_sc_hd__tap_1 TAP_13122 (  );
sky130_fd_sc_hd__tap_1 TAP_13123 (  );
sky130_fd_sc_hd__tap_1 TAP_13124 (  );
sky130_fd_sc_hd__tap_1 TAP_13125 (  );
sky130_fd_sc_hd__tap_1 TAP_13126 (  );
sky130_fd_sc_hd__tap_1 TAP_13127 (  );
sky130_fd_sc_hd__tap_1 TAP_13128 (  );
sky130_fd_sc_hd__tap_1 TAP_13129 (  );
sky130_fd_sc_hd__tap_1 TAP_1313 (  );
sky130_fd_sc_hd__tap_1 TAP_13130 (  );
sky130_fd_sc_hd__tap_1 TAP_13131 (  );
sky130_fd_sc_hd__tap_1 TAP_13132 (  );
sky130_fd_sc_hd__tap_1 TAP_13133 (  );
sky130_fd_sc_hd__tap_1 TAP_13134 (  );
sky130_fd_sc_hd__tap_1 TAP_13135 (  );
sky130_fd_sc_hd__tap_1 TAP_13136 (  );
sky130_fd_sc_hd__tap_1 TAP_13137 (  );
sky130_fd_sc_hd__tap_1 TAP_13138 (  );
sky130_fd_sc_hd__tap_1 TAP_13139 (  );
sky130_fd_sc_hd__tap_1 TAP_1314 (  );
sky130_fd_sc_hd__tap_1 TAP_13140 (  );
sky130_fd_sc_hd__tap_1 TAP_13141 (  );
sky130_fd_sc_hd__tap_1 TAP_13142 (  );
sky130_fd_sc_hd__tap_1 TAP_13143 (  );
sky130_fd_sc_hd__tap_1 TAP_13144 (  );
sky130_fd_sc_hd__tap_1 TAP_13145 (  );
sky130_fd_sc_hd__tap_1 TAP_13146 (  );
sky130_fd_sc_hd__tap_1 TAP_13147 (  );
sky130_fd_sc_hd__tap_1 TAP_13148 (  );
sky130_fd_sc_hd__tap_1 TAP_13149 (  );
sky130_fd_sc_hd__tap_1 TAP_1315 (  );
sky130_fd_sc_hd__tap_1 TAP_13150 (  );
sky130_fd_sc_hd__tap_1 TAP_13151 (  );
sky130_fd_sc_hd__tap_1 TAP_13152 (  );
sky130_fd_sc_hd__tap_1 TAP_13153 (  );
sky130_fd_sc_hd__tap_1 TAP_13154 (  );
sky130_fd_sc_hd__tap_1 TAP_13155 (  );
sky130_fd_sc_hd__tap_1 TAP_13156 (  );
sky130_fd_sc_hd__tap_1 TAP_13157 (  );
sky130_fd_sc_hd__tap_1 TAP_13158 (  );
sky130_fd_sc_hd__tap_1 TAP_13159 (  );
sky130_fd_sc_hd__tap_1 TAP_1316 (  );
sky130_fd_sc_hd__tap_1 TAP_13160 (  );
sky130_fd_sc_hd__tap_1 TAP_13161 (  );
sky130_fd_sc_hd__tap_1 TAP_13162 (  );
sky130_fd_sc_hd__tap_1 TAP_13163 (  );
sky130_fd_sc_hd__tap_1 TAP_13164 (  );
sky130_fd_sc_hd__tap_1 TAP_13165 (  );
sky130_fd_sc_hd__tap_1 TAP_13166 (  );
sky130_fd_sc_hd__tap_1 TAP_13167 (  );
sky130_fd_sc_hd__tap_1 TAP_13168 (  );
sky130_fd_sc_hd__tap_1 TAP_13169 (  );
sky130_fd_sc_hd__tap_1 TAP_1317 (  );
sky130_fd_sc_hd__tap_1 TAP_13170 (  );
sky130_fd_sc_hd__tap_1 TAP_13171 (  );
sky130_fd_sc_hd__tap_1 TAP_13172 (  );
sky130_fd_sc_hd__tap_1 TAP_13173 (  );
sky130_fd_sc_hd__tap_1 TAP_13174 (  );
sky130_fd_sc_hd__tap_1 TAP_13175 (  );
sky130_fd_sc_hd__tap_1 TAP_13176 (  );
sky130_fd_sc_hd__tap_1 TAP_13177 (  );
sky130_fd_sc_hd__tap_1 TAP_13178 (  );
sky130_fd_sc_hd__tap_1 TAP_13179 (  );
sky130_fd_sc_hd__tap_1 TAP_1318 (  );
sky130_fd_sc_hd__tap_1 TAP_13180 (  );
sky130_fd_sc_hd__tap_1 TAP_13181 (  );
sky130_fd_sc_hd__tap_1 TAP_13182 (  );
sky130_fd_sc_hd__tap_1 TAP_13183 (  );
sky130_fd_sc_hd__tap_1 TAP_13184 (  );
sky130_fd_sc_hd__tap_1 TAP_13185 (  );
sky130_fd_sc_hd__tap_1 TAP_13186 (  );
sky130_fd_sc_hd__tap_1 TAP_13187 (  );
sky130_fd_sc_hd__tap_1 TAP_13188 (  );
sky130_fd_sc_hd__tap_1 TAP_13189 (  );
sky130_fd_sc_hd__tap_1 TAP_1319 (  );
sky130_fd_sc_hd__tap_1 TAP_13190 (  );
sky130_fd_sc_hd__tap_1 TAP_13191 (  );
sky130_fd_sc_hd__tap_1 TAP_13192 (  );
sky130_fd_sc_hd__tap_1 TAP_13193 (  );
sky130_fd_sc_hd__tap_1 TAP_13194 (  );
sky130_fd_sc_hd__tap_1 TAP_13195 (  );
sky130_fd_sc_hd__tap_1 TAP_13196 (  );
sky130_fd_sc_hd__tap_1 TAP_13197 (  );
sky130_fd_sc_hd__tap_1 TAP_13198 (  );
sky130_fd_sc_hd__tap_1 TAP_13199 (  );
sky130_fd_sc_hd__tap_1 TAP_1320 (  );
sky130_fd_sc_hd__tap_1 TAP_13200 (  );
sky130_fd_sc_hd__tap_1 TAP_13201 (  );
sky130_fd_sc_hd__tap_1 TAP_13202 (  );
sky130_fd_sc_hd__tap_1 TAP_13203 (  );
sky130_fd_sc_hd__tap_1 TAP_13204 (  );
sky130_fd_sc_hd__tap_1 TAP_13205 (  );
sky130_fd_sc_hd__tap_1 TAP_13206 (  );
sky130_fd_sc_hd__tap_1 TAP_13207 (  );
sky130_fd_sc_hd__tap_1 TAP_13208 (  );
sky130_fd_sc_hd__tap_1 TAP_13209 (  );
sky130_fd_sc_hd__tap_1 TAP_1321 (  );
sky130_fd_sc_hd__tap_1 TAP_13210 (  );
sky130_fd_sc_hd__tap_1 TAP_13211 (  );
sky130_fd_sc_hd__tap_1 TAP_13212 (  );
sky130_fd_sc_hd__tap_1 TAP_13213 (  );
sky130_fd_sc_hd__tap_1 TAP_13214 (  );
sky130_fd_sc_hd__tap_1 TAP_13215 (  );
sky130_fd_sc_hd__tap_1 TAP_13216 (  );
sky130_fd_sc_hd__tap_1 TAP_13217 (  );
sky130_fd_sc_hd__tap_1 TAP_13218 (  );
sky130_fd_sc_hd__tap_1 TAP_13219 (  );
sky130_fd_sc_hd__tap_1 TAP_1322 (  );
sky130_fd_sc_hd__tap_1 TAP_13220 (  );
sky130_fd_sc_hd__tap_1 TAP_13221 (  );
sky130_fd_sc_hd__tap_1 TAP_13222 (  );
sky130_fd_sc_hd__tap_1 TAP_13223 (  );
sky130_fd_sc_hd__tap_1 TAP_13224 (  );
sky130_fd_sc_hd__tap_1 TAP_13225 (  );
sky130_fd_sc_hd__tap_1 TAP_13226 (  );
sky130_fd_sc_hd__tap_1 TAP_13227 (  );
sky130_fd_sc_hd__tap_1 TAP_13228 (  );
sky130_fd_sc_hd__tap_1 TAP_13229 (  );
sky130_fd_sc_hd__tap_1 TAP_1323 (  );
sky130_fd_sc_hd__tap_1 TAP_13230 (  );
sky130_fd_sc_hd__tap_1 TAP_13231 (  );
sky130_fd_sc_hd__tap_1 TAP_13232 (  );
sky130_fd_sc_hd__tap_1 TAP_13233 (  );
sky130_fd_sc_hd__tap_1 TAP_13234 (  );
sky130_fd_sc_hd__tap_1 TAP_13235 (  );
sky130_fd_sc_hd__tap_1 TAP_13236 (  );
sky130_fd_sc_hd__tap_1 TAP_13237 (  );
sky130_fd_sc_hd__tap_1 TAP_13238 (  );
sky130_fd_sc_hd__tap_1 TAP_13239 (  );
sky130_fd_sc_hd__tap_1 TAP_1324 (  );
sky130_fd_sc_hd__tap_1 TAP_13240 (  );
sky130_fd_sc_hd__tap_1 TAP_13241 (  );
sky130_fd_sc_hd__tap_1 TAP_13242 (  );
sky130_fd_sc_hd__tap_1 TAP_13243 (  );
sky130_fd_sc_hd__tap_1 TAP_13244 (  );
sky130_fd_sc_hd__tap_1 TAP_13245 (  );
sky130_fd_sc_hd__tap_1 TAP_13246 (  );
sky130_fd_sc_hd__tap_1 TAP_13247 (  );
sky130_fd_sc_hd__tap_1 TAP_13248 (  );
sky130_fd_sc_hd__tap_1 TAP_13249 (  );
sky130_fd_sc_hd__tap_1 TAP_1325 (  );
sky130_fd_sc_hd__tap_1 TAP_13250 (  );
sky130_fd_sc_hd__tap_1 TAP_13251 (  );
sky130_fd_sc_hd__tap_1 TAP_13252 (  );
sky130_fd_sc_hd__tap_1 TAP_13253 (  );
sky130_fd_sc_hd__tap_1 TAP_13254 (  );
sky130_fd_sc_hd__tap_1 TAP_13255 (  );
sky130_fd_sc_hd__tap_1 TAP_13256 (  );
sky130_fd_sc_hd__tap_1 TAP_13257 (  );
sky130_fd_sc_hd__tap_1 TAP_13258 (  );
sky130_fd_sc_hd__tap_1 TAP_13259 (  );
sky130_fd_sc_hd__tap_1 TAP_1326 (  );
sky130_fd_sc_hd__tap_1 TAP_13260 (  );
sky130_fd_sc_hd__tap_1 TAP_13261 (  );
sky130_fd_sc_hd__tap_1 TAP_13262 (  );
sky130_fd_sc_hd__tap_1 TAP_13263 (  );
sky130_fd_sc_hd__tap_1 TAP_13264 (  );
sky130_fd_sc_hd__tap_1 TAP_13265 (  );
sky130_fd_sc_hd__tap_1 TAP_13266 (  );
sky130_fd_sc_hd__tap_1 TAP_13267 (  );
sky130_fd_sc_hd__tap_1 TAP_13268 (  );
sky130_fd_sc_hd__tap_1 TAP_13269 (  );
sky130_fd_sc_hd__tap_1 TAP_1327 (  );
sky130_fd_sc_hd__tap_1 TAP_13270 (  );
sky130_fd_sc_hd__tap_1 TAP_13271 (  );
sky130_fd_sc_hd__tap_1 TAP_13272 (  );
sky130_fd_sc_hd__tap_1 TAP_13273 (  );
sky130_fd_sc_hd__tap_1 TAP_13274 (  );
sky130_fd_sc_hd__tap_1 TAP_13275 (  );
sky130_fd_sc_hd__tap_1 TAP_13276 (  );
sky130_fd_sc_hd__tap_1 TAP_13277 (  );
sky130_fd_sc_hd__tap_1 TAP_13278 (  );
sky130_fd_sc_hd__tap_1 TAP_13279 (  );
sky130_fd_sc_hd__tap_1 TAP_1328 (  );
sky130_fd_sc_hd__tap_1 TAP_13280 (  );
sky130_fd_sc_hd__tap_1 TAP_13281 (  );
sky130_fd_sc_hd__tap_1 TAP_13282 (  );
sky130_fd_sc_hd__tap_1 TAP_13283 (  );
sky130_fd_sc_hd__tap_1 TAP_13284 (  );
sky130_fd_sc_hd__tap_1 TAP_13285 (  );
sky130_fd_sc_hd__tap_1 TAP_13286 (  );
sky130_fd_sc_hd__tap_1 TAP_13287 (  );
sky130_fd_sc_hd__tap_1 TAP_13288 (  );
sky130_fd_sc_hd__tap_1 TAP_13289 (  );
sky130_fd_sc_hd__tap_1 TAP_1329 (  );
sky130_fd_sc_hd__tap_1 TAP_13290 (  );
sky130_fd_sc_hd__tap_1 TAP_13291 (  );
sky130_fd_sc_hd__tap_1 TAP_13292 (  );
sky130_fd_sc_hd__tap_1 TAP_13293 (  );
sky130_fd_sc_hd__tap_1 TAP_13294 (  );
sky130_fd_sc_hd__tap_1 TAP_13295 (  );
sky130_fd_sc_hd__tap_1 TAP_13296 (  );
sky130_fd_sc_hd__tap_1 TAP_13297 (  );
sky130_fd_sc_hd__tap_1 TAP_13298 (  );
sky130_fd_sc_hd__tap_1 TAP_13299 (  );
sky130_fd_sc_hd__tap_1 TAP_1330 (  );
sky130_fd_sc_hd__tap_1 TAP_13300 (  );
sky130_fd_sc_hd__tap_1 TAP_13301 (  );
sky130_fd_sc_hd__tap_1 TAP_13302 (  );
sky130_fd_sc_hd__tap_1 TAP_13303 (  );
sky130_fd_sc_hd__tap_1 TAP_13304 (  );
sky130_fd_sc_hd__tap_1 TAP_13305 (  );
sky130_fd_sc_hd__tap_1 TAP_13306 (  );
sky130_fd_sc_hd__tap_1 TAP_13307 (  );
sky130_fd_sc_hd__tap_1 TAP_13308 (  );
sky130_fd_sc_hd__tap_1 TAP_13309 (  );
sky130_fd_sc_hd__tap_1 TAP_1331 (  );
sky130_fd_sc_hd__tap_1 TAP_13310 (  );
sky130_fd_sc_hd__tap_1 TAP_13311 (  );
sky130_fd_sc_hd__tap_1 TAP_13312 (  );
sky130_fd_sc_hd__tap_1 TAP_13313 (  );
sky130_fd_sc_hd__tap_1 TAP_13314 (  );
sky130_fd_sc_hd__tap_1 TAP_13315 (  );
sky130_fd_sc_hd__tap_1 TAP_13316 (  );
sky130_fd_sc_hd__tap_1 TAP_13317 (  );
sky130_fd_sc_hd__tap_1 TAP_13318 (  );
sky130_fd_sc_hd__tap_1 TAP_13319 (  );
sky130_fd_sc_hd__tap_1 TAP_1332 (  );
sky130_fd_sc_hd__tap_1 TAP_13320 (  );
sky130_fd_sc_hd__tap_1 TAP_13321 (  );
sky130_fd_sc_hd__tap_1 TAP_13322 (  );
sky130_fd_sc_hd__tap_1 TAP_13323 (  );
sky130_fd_sc_hd__tap_1 TAP_13324 (  );
sky130_fd_sc_hd__tap_1 TAP_13325 (  );
sky130_fd_sc_hd__tap_1 TAP_13326 (  );
sky130_fd_sc_hd__tap_1 TAP_13327 (  );
sky130_fd_sc_hd__tap_1 TAP_13328 (  );
sky130_fd_sc_hd__tap_1 TAP_13329 (  );
sky130_fd_sc_hd__tap_1 TAP_1333 (  );
sky130_fd_sc_hd__tap_1 TAP_13330 (  );
sky130_fd_sc_hd__tap_1 TAP_13331 (  );
sky130_fd_sc_hd__tap_1 TAP_13332 (  );
sky130_fd_sc_hd__tap_1 TAP_13333 (  );
sky130_fd_sc_hd__tap_1 TAP_13334 (  );
sky130_fd_sc_hd__tap_1 TAP_13335 (  );
sky130_fd_sc_hd__tap_1 TAP_13336 (  );
sky130_fd_sc_hd__tap_1 TAP_13337 (  );
sky130_fd_sc_hd__tap_1 TAP_13338 (  );
sky130_fd_sc_hd__tap_1 TAP_13339 (  );
sky130_fd_sc_hd__tap_1 TAP_1334 (  );
sky130_fd_sc_hd__tap_1 TAP_13340 (  );
sky130_fd_sc_hd__tap_1 TAP_13341 (  );
sky130_fd_sc_hd__tap_1 TAP_13342 (  );
sky130_fd_sc_hd__tap_1 TAP_13343 (  );
sky130_fd_sc_hd__tap_1 TAP_13344 (  );
sky130_fd_sc_hd__tap_1 TAP_13345 (  );
sky130_fd_sc_hd__tap_1 TAP_13346 (  );
sky130_fd_sc_hd__tap_1 TAP_13347 (  );
sky130_fd_sc_hd__tap_1 TAP_13348 (  );
sky130_fd_sc_hd__tap_1 TAP_13349 (  );
sky130_fd_sc_hd__tap_1 TAP_1335 (  );
sky130_fd_sc_hd__tap_1 TAP_13350 (  );
sky130_fd_sc_hd__tap_1 TAP_13351 (  );
sky130_fd_sc_hd__tap_1 TAP_13352 (  );
sky130_fd_sc_hd__tap_1 TAP_13353 (  );
sky130_fd_sc_hd__tap_1 TAP_13354 (  );
sky130_fd_sc_hd__tap_1 TAP_13355 (  );
sky130_fd_sc_hd__tap_1 TAP_13356 (  );
sky130_fd_sc_hd__tap_1 TAP_13357 (  );
sky130_fd_sc_hd__tap_1 TAP_13358 (  );
sky130_fd_sc_hd__tap_1 TAP_13359 (  );
sky130_fd_sc_hd__tap_1 TAP_1336 (  );
sky130_fd_sc_hd__tap_1 TAP_13360 (  );
sky130_fd_sc_hd__tap_1 TAP_13361 (  );
sky130_fd_sc_hd__tap_1 TAP_13362 (  );
sky130_fd_sc_hd__tap_1 TAP_13363 (  );
sky130_fd_sc_hd__tap_1 TAP_13364 (  );
sky130_fd_sc_hd__tap_1 TAP_13365 (  );
sky130_fd_sc_hd__tap_1 TAP_13366 (  );
sky130_fd_sc_hd__tap_1 TAP_13367 (  );
sky130_fd_sc_hd__tap_1 TAP_13368 (  );
sky130_fd_sc_hd__tap_1 TAP_13369 (  );
sky130_fd_sc_hd__tap_1 TAP_1337 (  );
sky130_fd_sc_hd__tap_1 TAP_13370 (  );
sky130_fd_sc_hd__tap_1 TAP_13371 (  );
sky130_fd_sc_hd__tap_1 TAP_13372 (  );
sky130_fd_sc_hd__tap_1 TAP_13373 (  );
sky130_fd_sc_hd__tap_1 TAP_13374 (  );
sky130_fd_sc_hd__tap_1 TAP_13375 (  );
sky130_fd_sc_hd__tap_1 TAP_13376 (  );
sky130_fd_sc_hd__tap_1 TAP_13377 (  );
sky130_fd_sc_hd__tap_1 TAP_13378 (  );
sky130_fd_sc_hd__tap_1 TAP_13379 (  );
sky130_fd_sc_hd__tap_1 TAP_1338 (  );
sky130_fd_sc_hd__tap_1 TAP_13380 (  );
sky130_fd_sc_hd__tap_1 TAP_13381 (  );
sky130_fd_sc_hd__tap_1 TAP_13382 (  );
sky130_fd_sc_hd__tap_1 TAP_13383 (  );
sky130_fd_sc_hd__tap_1 TAP_13384 (  );
sky130_fd_sc_hd__tap_1 TAP_13385 (  );
sky130_fd_sc_hd__tap_1 TAP_13386 (  );
sky130_fd_sc_hd__tap_1 TAP_13387 (  );
sky130_fd_sc_hd__tap_1 TAP_13388 (  );
sky130_fd_sc_hd__tap_1 TAP_13389 (  );
sky130_fd_sc_hd__tap_1 TAP_1339 (  );
sky130_fd_sc_hd__tap_1 TAP_13390 (  );
sky130_fd_sc_hd__tap_1 TAP_13391 (  );
sky130_fd_sc_hd__tap_1 TAP_13392 (  );
sky130_fd_sc_hd__tap_1 TAP_13393 (  );
sky130_fd_sc_hd__tap_1 TAP_13394 (  );
sky130_fd_sc_hd__tap_1 TAP_13395 (  );
sky130_fd_sc_hd__tap_1 TAP_13396 (  );
sky130_fd_sc_hd__tap_1 TAP_13397 (  );
sky130_fd_sc_hd__tap_1 TAP_13398 (  );
sky130_fd_sc_hd__tap_1 TAP_13399 (  );
sky130_fd_sc_hd__tap_1 TAP_1340 (  );
sky130_fd_sc_hd__tap_1 TAP_13400 (  );
sky130_fd_sc_hd__tap_1 TAP_13401 (  );
sky130_fd_sc_hd__tap_1 TAP_13402 (  );
sky130_fd_sc_hd__tap_1 TAP_13403 (  );
sky130_fd_sc_hd__tap_1 TAP_13404 (  );
sky130_fd_sc_hd__tap_1 TAP_13405 (  );
sky130_fd_sc_hd__tap_1 TAP_13406 (  );
sky130_fd_sc_hd__tap_1 TAP_13407 (  );
sky130_fd_sc_hd__tap_1 TAP_13408 (  );
sky130_fd_sc_hd__tap_1 TAP_13409 (  );
sky130_fd_sc_hd__tap_1 TAP_1341 (  );
sky130_fd_sc_hd__tap_1 TAP_13410 (  );
sky130_fd_sc_hd__tap_1 TAP_13411 (  );
sky130_fd_sc_hd__tap_1 TAP_13412 (  );
sky130_fd_sc_hd__tap_1 TAP_13413 (  );
sky130_fd_sc_hd__tap_1 TAP_13414 (  );
sky130_fd_sc_hd__tap_1 TAP_13415 (  );
sky130_fd_sc_hd__tap_1 TAP_13416 (  );
sky130_fd_sc_hd__tap_1 TAP_13417 (  );
sky130_fd_sc_hd__tap_1 TAP_13418 (  );
sky130_fd_sc_hd__tap_1 TAP_13419 (  );
sky130_fd_sc_hd__tap_1 TAP_1342 (  );
sky130_fd_sc_hd__tap_1 TAP_13420 (  );
sky130_fd_sc_hd__tap_1 TAP_13421 (  );
sky130_fd_sc_hd__tap_1 TAP_13422 (  );
sky130_fd_sc_hd__tap_1 TAP_13423 (  );
sky130_fd_sc_hd__tap_1 TAP_13424 (  );
sky130_fd_sc_hd__tap_1 TAP_13425 (  );
sky130_fd_sc_hd__tap_1 TAP_13426 (  );
sky130_fd_sc_hd__tap_1 TAP_13427 (  );
sky130_fd_sc_hd__tap_1 TAP_13428 (  );
sky130_fd_sc_hd__tap_1 TAP_13429 (  );
sky130_fd_sc_hd__tap_1 TAP_1343 (  );
sky130_fd_sc_hd__tap_1 TAP_13430 (  );
sky130_fd_sc_hd__tap_1 TAP_13431 (  );
sky130_fd_sc_hd__tap_1 TAP_13432 (  );
sky130_fd_sc_hd__tap_1 TAP_13433 (  );
sky130_fd_sc_hd__tap_1 TAP_13434 (  );
sky130_fd_sc_hd__tap_1 TAP_13435 (  );
sky130_fd_sc_hd__tap_1 TAP_13436 (  );
sky130_fd_sc_hd__tap_1 TAP_13437 (  );
sky130_fd_sc_hd__tap_1 TAP_13438 (  );
sky130_fd_sc_hd__tap_1 TAP_13439 (  );
sky130_fd_sc_hd__tap_1 TAP_1344 (  );
sky130_fd_sc_hd__tap_1 TAP_13440 (  );
sky130_fd_sc_hd__tap_1 TAP_13441 (  );
sky130_fd_sc_hd__tap_1 TAP_13442 (  );
sky130_fd_sc_hd__tap_1 TAP_13443 (  );
sky130_fd_sc_hd__tap_1 TAP_13444 (  );
sky130_fd_sc_hd__tap_1 TAP_13445 (  );
sky130_fd_sc_hd__tap_1 TAP_13446 (  );
sky130_fd_sc_hd__tap_1 TAP_13447 (  );
sky130_fd_sc_hd__tap_1 TAP_13448 (  );
sky130_fd_sc_hd__tap_1 TAP_13449 (  );
sky130_fd_sc_hd__tap_1 TAP_1345 (  );
sky130_fd_sc_hd__tap_1 TAP_13450 (  );
sky130_fd_sc_hd__tap_1 TAP_13451 (  );
sky130_fd_sc_hd__tap_1 TAP_13452 (  );
sky130_fd_sc_hd__tap_1 TAP_13453 (  );
sky130_fd_sc_hd__tap_1 TAP_13454 (  );
sky130_fd_sc_hd__tap_1 TAP_13455 (  );
sky130_fd_sc_hd__tap_1 TAP_13456 (  );
sky130_fd_sc_hd__tap_1 TAP_13457 (  );
sky130_fd_sc_hd__tap_1 TAP_13458 (  );
sky130_fd_sc_hd__tap_1 TAP_13459 (  );
sky130_fd_sc_hd__tap_1 TAP_1346 (  );
sky130_fd_sc_hd__tap_1 TAP_13460 (  );
sky130_fd_sc_hd__tap_1 TAP_13461 (  );
sky130_fd_sc_hd__tap_1 TAP_13462 (  );
sky130_fd_sc_hd__tap_1 TAP_13463 (  );
sky130_fd_sc_hd__tap_1 TAP_13464 (  );
sky130_fd_sc_hd__tap_1 TAP_13465 (  );
sky130_fd_sc_hd__tap_1 TAP_13466 (  );
sky130_fd_sc_hd__tap_1 TAP_13467 (  );
sky130_fd_sc_hd__tap_1 TAP_13468 (  );
sky130_fd_sc_hd__tap_1 TAP_13469 (  );
sky130_fd_sc_hd__tap_1 TAP_1347 (  );
sky130_fd_sc_hd__tap_1 TAP_13470 (  );
sky130_fd_sc_hd__tap_1 TAP_13471 (  );
sky130_fd_sc_hd__tap_1 TAP_13472 (  );
sky130_fd_sc_hd__tap_1 TAP_13473 (  );
sky130_fd_sc_hd__tap_1 TAP_13474 (  );
sky130_fd_sc_hd__tap_1 TAP_13475 (  );
sky130_fd_sc_hd__tap_1 TAP_13476 (  );
sky130_fd_sc_hd__tap_1 TAP_13477 (  );
sky130_fd_sc_hd__tap_1 TAP_13478 (  );
sky130_fd_sc_hd__tap_1 TAP_13479 (  );
sky130_fd_sc_hd__tap_1 TAP_1348 (  );
sky130_fd_sc_hd__tap_1 TAP_13480 (  );
sky130_fd_sc_hd__tap_1 TAP_13481 (  );
sky130_fd_sc_hd__tap_1 TAP_13482 (  );
sky130_fd_sc_hd__tap_1 TAP_13483 (  );
sky130_fd_sc_hd__tap_1 TAP_13484 (  );
sky130_fd_sc_hd__tap_1 TAP_13485 (  );
sky130_fd_sc_hd__tap_1 TAP_13486 (  );
sky130_fd_sc_hd__tap_1 TAP_13487 (  );
sky130_fd_sc_hd__tap_1 TAP_13488 (  );
sky130_fd_sc_hd__tap_1 TAP_13489 (  );
sky130_fd_sc_hd__tap_1 TAP_1349 (  );
sky130_fd_sc_hd__tap_1 TAP_13490 (  );
sky130_fd_sc_hd__tap_1 TAP_13491 (  );
sky130_fd_sc_hd__tap_1 TAP_13492 (  );
sky130_fd_sc_hd__tap_1 TAP_13493 (  );
sky130_fd_sc_hd__tap_1 TAP_13494 (  );
sky130_fd_sc_hd__tap_1 TAP_13495 (  );
sky130_fd_sc_hd__tap_1 TAP_13496 (  );
sky130_fd_sc_hd__tap_1 TAP_13497 (  );
sky130_fd_sc_hd__tap_1 TAP_13498 (  );
sky130_fd_sc_hd__tap_1 TAP_13499 (  );
sky130_fd_sc_hd__tap_1 TAP_1350 (  );
sky130_fd_sc_hd__tap_1 TAP_13500 (  );
sky130_fd_sc_hd__tap_1 TAP_13501 (  );
sky130_fd_sc_hd__tap_1 TAP_13502 (  );
sky130_fd_sc_hd__tap_1 TAP_13503 (  );
sky130_fd_sc_hd__tap_1 TAP_13504 (  );
sky130_fd_sc_hd__tap_1 TAP_13505 (  );
sky130_fd_sc_hd__tap_1 TAP_13506 (  );
sky130_fd_sc_hd__tap_1 TAP_13507 (  );
sky130_fd_sc_hd__tap_1 TAP_13508 (  );
sky130_fd_sc_hd__tap_1 TAP_13509 (  );
sky130_fd_sc_hd__tap_1 TAP_1351 (  );
sky130_fd_sc_hd__tap_1 TAP_13510 (  );
sky130_fd_sc_hd__tap_1 TAP_13511 (  );
sky130_fd_sc_hd__tap_1 TAP_13512 (  );
sky130_fd_sc_hd__tap_1 TAP_13513 (  );
sky130_fd_sc_hd__tap_1 TAP_13514 (  );
sky130_fd_sc_hd__tap_1 TAP_13515 (  );
sky130_fd_sc_hd__tap_1 TAP_13516 (  );
sky130_fd_sc_hd__tap_1 TAP_13517 (  );
sky130_fd_sc_hd__tap_1 TAP_13518 (  );
sky130_fd_sc_hd__tap_1 TAP_13519 (  );
sky130_fd_sc_hd__tap_1 TAP_1352 (  );
sky130_fd_sc_hd__tap_1 TAP_13520 (  );
sky130_fd_sc_hd__tap_1 TAP_13521 (  );
sky130_fd_sc_hd__tap_1 TAP_13522 (  );
sky130_fd_sc_hd__tap_1 TAP_13523 (  );
sky130_fd_sc_hd__tap_1 TAP_13524 (  );
sky130_fd_sc_hd__tap_1 TAP_13525 (  );
sky130_fd_sc_hd__tap_1 TAP_13526 (  );
sky130_fd_sc_hd__tap_1 TAP_13527 (  );
sky130_fd_sc_hd__tap_1 TAP_13528 (  );
sky130_fd_sc_hd__tap_1 TAP_13529 (  );
sky130_fd_sc_hd__tap_1 TAP_1353 (  );
sky130_fd_sc_hd__tap_1 TAP_13530 (  );
sky130_fd_sc_hd__tap_1 TAP_13531 (  );
sky130_fd_sc_hd__tap_1 TAP_13532 (  );
sky130_fd_sc_hd__tap_1 TAP_13533 (  );
sky130_fd_sc_hd__tap_1 TAP_13534 (  );
sky130_fd_sc_hd__tap_1 TAP_13535 (  );
sky130_fd_sc_hd__tap_1 TAP_13536 (  );
sky130_fd_sc_hd__tap_1 TAP_13537 (  );
sky130_fd_sc_hd__tap_1 TAP_13538 (  );
sky130_fd_sc_hd__tap_1 TAP_13539 (  );
sky130_fd_sc_hd__tap_1 TAP_1354 (  );
sky130_fd_sc_hd__tap_1 TAP_13540 (  );
sky130_fd_sc_hd__tap_1 TAP_13541 (  );
sky130_fd_sc_hd__tap_1 TAP_13542 (  );
sky130_fd_sc_hd__tap_1 TAP_13543 (  );
sky130_fd_sc_hd__tap_1 TAP_13544 (  );
sky130_fd_sc_hd__tap_1 TAP_13545 (  );
sky130_fd_sc_hd__tap_1 TAP_13546 (  );
sky130_fd_sc_hd__tap_1 TAP_13547 (  );
sky130_fd_sc_hd__tap_1 TAP_13548 (  );
sky130_fd_sc_hd__tap_1 TAP_13549 (  );
sky130_fd_sc_hd__tap_1 TAP_1355 (  );
sky130_fd_sc_hd__tap_1 TAP_13550 (  );
sky130_fd_sc_hd__tap_1 TAP_13551 (  );
sky130_fd_sc_hd__tap_1 TAP_13552 (  );
sky130_fd_sc_hd__tap_1 TAP_13553 (  );
sky130_fd_sc_hd__tap_1 TAP_13554 (  );
sky130_fd_sc_hd__tap_1 TAP_13555 (  );
sky130_fd_sc_hd__tap_1 TAP_13556 (  );
sky130_fd_sc_hd__tap_1 TAP_13557 (  );
sky130_fd_sc_hd__tap_1 TAP_13558 (  );
sky130_fd_sc_hd__tap_1 TAP_13559 (  );
sky130_fd_sc_hd__tap_1 TAP_1356 (  );
sky130_fd_sc_hd__tap_1 TAP_13560 (  );
sky130_fd_sc_hd__tap_1 TAP_13561 (  );
sky130_fd_sc_hd__tap_1 TAP_13562 (  );
sky130_fd_sc_hd__tap_1 TAP_13563 (  );
sky130_fd_sc_hd__tap_1 TAP_13564 (  );
sky130_fd_sc_hd__tap_1 TAP_13565 (  );
sky130_fd_sc_hd__tap_1 TAP_13566 (  );
sky130_fd_sc_hd__tap_1 TAP_13567 (  );
sky130_fd_sc_hd__tap_1 TAP_13568 (  );
sky130_fd_sc_hd__tap_1 TAP_13569 (  );
sky130_fd_sc_hd__tap_1 TAP_1357 (  );
sky130_fd_sc_hd__tap_1 TAP_13570 (  );
sky130_fd_sc_hd__tap_1 TAP_13571 (  );
sky130_fd_sc_hd__tap_1 TAP_13572 (  );
sky130_fd_sc_hd__tap_1 TAP_13573 (  );
sky130_fd_sc_hd__tap_1 TAP_13574 (  );
sky130_fd_sc_hd__tap_1 TAP_13575 (  );
sky130_fd_sc_hd__tap_1 TAP_13576 (  );
sky130_fd_sc_hd__tap_1 TAP_13577 (  );
sky130_fd_sc_hd__tap_1 TAP_13578 (  );
sky130_fd_sc_hd__tap_1 TAP_13579 (  );
sky130_fd_sc_hd__tap_1 TAP_1358 (  );
sky130_fd_sc_hd__tap_1 TAP_13580 (  );
sky130_fd_sc_hd__tap_1 TAP_13581 (  );
sky130_fd_sc_hd__tap_1 TAP_13582 (  );
sky130_fd_sc_hd__tap_1 TAP_13583 (  );
sky130_fd_sc_hd__tap_1 TAP_13584 (  );
sky130_fd_sc_hd__tap_1 TAP_13585 (  );
sky130_fd_sc_hd__tap_1 TAP_13586 (  );
sky130_fd_sc_hd__tap_1 TAP_13587 (  );
sky130_fd_sc_hd__tap_1 TAP_13588 (  );
sky130_fd_sc_hd__tap_1 TAP_13589 (  );
sky130_fd_sc_hd__tap_1 TAP_1359 (  );
sky130_fd_sc_hd__tap_1 TAP_13590 (  );
sky130_fd_sc_hd__tap_1 TAP_13591 (  );
sky130_fd_sc_hd__tap_1 TAP_13592 (  );
sky130_fd_sc_hd__tap_1 TAP_13593 (  );
sky130_fd_sc_hd__tap_1 TAP_13594 (  );
sky130_fd_sc_hd__tap_1 TAP_13595 (  );
sky130_fd_sc_hd__tap_1 TAP_13596 (  );
sky130_fd_sc_hd__tap_1 TAP_13597 (  );
sky130_fd_sc_hd__tap_1 TAP_13598 (  );
sky130_fd_sc_hd__tap_1 TAP_13599 (  );
sky130_fd_sc_hd__tap_1 TAP_1360 (  );
sky130_fd_sc_hd__tap_1 TAP_13600 (  );
sky130_fd_sc_hd__tap_1 TAP_13601 (  );
sky130_fd_sc_hd__tap_1 TAP_13602 (  );
sky130_fd_sc_hd__tap_1 TAP_13603 (  );
sky130_fd_sc_hd__tap_1 TAP_13604 (  );
sky130_fd_sc_hd__tap_1 TAP_13605 (  );
sky130_fd_sc_hd__tap_1 TAP_13606 (  );
sky130_fd_sc_hd__tap_1 TAP_13607 (  );
sky130_fd_sc_hd__tap_1 TAP_13608 (  );
sky130_fd_sc_hd__tap_1 TAP_13609 (  );
sky130_fd_sc_hd__tap_1 TAP_1361 (  );
sky130_fd_sc_hd__tap_1 TAP_13610 (  );
sky130_fd_sc_hd__tap_1 TAP_13611 (  );
sky130_fd_sc_hd__tap_1 TAP_13612 (  );
sky130_fd_sc_hd__tap_1 TAP_13613 (  );
sky130_fd_sc_hd__tap_1 TAP_13614 (  );
sky130_fd_sc_hd__tap_1 TAP_13615 (  );
sky130_fd_sc_hd__tap_1 TAP_13616 (  );
sky130_fd_sc_hd__tap_1 TAP_13617 (  );
sky130_fd_sc_hd__tap_1 TAP_13618 (  );
sky130_fd_sc_hd__tap_1 TAP_13619 (  );
sky130_fd_sc_hd__tap_1 TAP_1362 (  );
sky130_fd_sc_hd__tap_1 TAP_13620 (  );
sky130_fd_sc_hd__tap_1 TAP_13621 (  );
sky130_fd_sc_hd__tap_1 TAP_13622 (  );
sky130_fd_sc_hd__tap_1 TAP_13623 (  );
sky130_fd_sc_hd__tap_1 TAP_13624 (  );
sky130_fd_sc_hd__tap_1 TAP_13625 (  );
sky130_fd_sc_hd__tap_1 TAP_13626 (  );
sky130_fd_sc_hd__tap_1 TAP_13627 (  );
sky130_fd_sc_hd__tap_1 TAP_13628 (  );
sky130_fd_sc_hd__tap_1 TAP_13629 (  );
sky130_fd_sc_hd__tap_1 TAP_1363 (  );
sky130_fd_sc_hd__tap_1 TAP_13630 (  );
sky130_fd_sc_hd__tap_1 TAP_13631 (  );
sky130_fd_sc_hd__tap_1 TAP_13632 (  );
sky130_fd_sc_hd__tap_1 TAP_13633 (  );
sky130_fd_sc_hd__tap_1 TAP_13634 (  );
sky130_fd_sc_hd__tap_1 TAP_13635 (  );
sky130_fd_sc_hd__tap_1 TAP_13636 (  );
sky130_fd_sc_hd__tap_1 TAP_13637 (  );
sky130_fd_sc_hd__tap_1 TAP_13638 (  );
sky130_fd_sc_hd__tap_1 TAP_13639 (  );
sky130_fd_sc_hd__tap_1 TAP_1364 (  );
sky130_fd_sc_hd__tap_1 TAP_13640 (  );
sky130_fd_sc_hd__tap_1 TAP_13641 (  );
sky130_fd_sc_hd__tap_1 TAP_13642 (  );
sky130_fd_sc_hd__tap_1 TAP_13643 (  );
sky130_fd_sc_hd__tap_1 TAP_13644 (  );
sky130_fd_sc_hd__tap_1 TAP_13645 (  );
sky130_fd_sc_hd__tap_1 TAP_13646 (  );
sky130_fd_sc_hd__tap_1 TAP_13647 (  );
sky130_fd_sc_hd__tap_1 TAP_13648 (  );
sky130_fd_sc_hd__tap_1 TAP_13649 (  );
sky130_fd_sc_hd__tap_1 TAP_1365 (  );
sky130_fd_sc_hd__tap_1 TAP_13650 (  );
sky130_fd_sc_hd__tap_1 TAP_13651 (  );
sky130_fd_sc_hd__tap_1 TAP_13652 (  );
sky130_fd_sc_hd__tap_1 TAP_13653 (  );
sky130_fd_sc_hd__tap_1 TAP_13654 (  );
sky130_fd_sc_hd__tap_1 TAP_13655 (  );
sky130_fd_sc_hd__tap_1 TAP_13656 (  );
sky130_fd_sc_hd__tap_1 TAP_13657 (  );
sky130_fd_sc_hd__tap_1 TAP_13658 (  );
sky130_fd_sc_hd__tap_1 TAP_13659 (  );
sky130_fd_sc_hd__tap_1 TAP_1366 (  );
sky130_fd_sc_hd__tap_1 TAP_13660 (  );
sky130_fd_sc_hd__tap_1 TAP_13661 (  );
sky130_fd_sc_hd__tap_1 TAP_13662 (  );
sky130_fd_sc_hd__tap_1 TAP_13663 (  );
sky130_fd_sc_hd__tap_1 TAP_13664 (  );
sky130_fd_sc_hd__tap_1 TAP_13665 (  );
sky130_fd_sc_hd__tap_1 TAP_13666 (  );
sky130_fd_sc_hd__tap_1 TAP_13667 (  );
sky130_fd_sc_hd__tap_1 TAP_13668 (  );
sky130_fd_sc_hd__tap_1 TAP_13669 (  );
sky130_fd_sc_hd__tap_1 TAP_1367 (  );
sky130_fd_sc_hd__tap_1 TAP_13670 (  );
sky130_fd_sc_hd__tap_1 TAP_13671 (  );
sky130_fd_sc_hd__tap_1 TAP_13672 (  );
sky130_fd_sc_hd__tap_1 TAP_13673 (  );
sky130_fd_sc_hd__tap_1 TAP_13674 (  );
sky130_fd_sc_hd__tap_1 TAP_13675 (  );
sky130_fd_sc_hd__tap_1 TAP_13676 (  );
sky130_fd_sc_hd__tap_1 TAP_13677 (  );
sky130_fd_sc_hd__tap_1 TAP_13678 (  );
sky130_fd_sc_hd__tap_1 TAP_13679 (  );
sky130_fd_sc_hd__tap_1 TAP_1368 (  );
sky130_fd_sc_hd__tap_1 TAP_13680 (  );
sky130_fd_sc_hd__tap_1 TAP_13681 (  );
sky130_fd_sc_hd__tap_1 TAP_13682 (  );
sky130_fd_sc_hd__tap_1 TAP_13683 (  );
sky130_fd_sc_hd__tap_1 TAP_13684 (  );
sky130_fd_sc_hd__tap_1 TAP_13685 (  );
sky130_fd_sc_hd__tap_1 TAP_13686 (  );
sky130_fd_sc_hd__tap_1 TAP_13687 (  );
sky130_fd_sc_hd__tap_1 TAP_13688 (  );
sky130_fd_sc_hd__tap_1 TAP_13689 (  );
sky130_fd_sc_hd__tap_1 TAP_1369 (  );
sky130_fd_sc_hd__tap_1 TAP_13690 (  );
sky130_fd_sc_hd__tap_1 TAP_13691 (  );
sky130_fd_sc_hd__tap_1 TAP_13692 (  );
sky130_fd_sc_hd__tap_1 TAP_13693 (  );
sky130_fd_sc_hd__tap_1 TAP_13694 (  );
sky130_fd_sc_hd__tap_1 TAP_13695 (  );
sky130_fd_sc_hd__tap_1 TAP_13696 (  );
sky130_fd_sc_hd__tap_1 TAP_13697 (  );
sky130_fd_sc_hd__tap_1 TAP_13698 (  );
sky130_fd_sc_hd__tap_1 TAP_13699 (  );
sky130_fd_sc_hd__tap_1 TAP_1370 (  );
sky130_fd_sc_hd__tap_1 TAP_13700 (  );
sky130_fd_sc_hd__tap_1 TAP_13701 (  );
sky130_fd_sc_hd__tap_1 TAP_13702 (  );
sky130_fd_sc_hd__tap_1 TAP_13703 (  );
sky130_fd_sc_hd__tap_1 TAP_13704 (  );
sky130_fd_sc_hd__tap_1 TAP_13705 (  );
sky130_fd_sc_hd__tap_1 TAP_13706 (  );
sky130_fd_sc_hd__tap_1 TAP_13707 (  );
sky130_fd_sc_hd__tap_1 TAP_13708 (  );
sky130_fd_sc_hd__tap_1 TAP_13709 (  );
sky130_fd_sc_hd__tap_1 TAP_1371 (  );
sky130_fd_sc_hd__tap_1 TAP_13710 (  );
sky130_fd_sc_hd__tap_1 TAP_13711 (  );
sky130_fd_sc_hd__tap_1 TAP_13712 (  );
sky130_fd_sc_hd__tap_1 TAP_13713 (  );
sky130_fd_sc_hd__tap_1 TAP_13714 (  );
sky130_fd_sc_hd__tap_1 TAP_13715 (  );
sky130_fd_sc_hd__tap_1 TAP_13716 (  );
sky130_fd_sc_hd__tap_1 TAP_13717 (  );
sky130_fd_sc_hd__tap_1 TAP_13718 (  );
sky130_fd_sc_hd__tap_1 TAP_13719 (  );
sky130_fd_sc_hd__tap_1 TAP_1372 (  );
sky130_fd_sc_hd__tap_1 TAP_13720 (  );
sky130_fd_sc_hd__tap_1 TAP_13721 (  );
sky130_fd_sc_hd__tap_1 TAP_13722 (  );
sky130_fd_sc_hd__tap_1 TAP_13723 (  );
sky130_fd_sc_hd__tap_1 TAP_13724 (  );
sky130_fd_sc_hd__tap_1 TAP_13725 (  );
sky130_fd_sc_hd__tap_1 TAP_13726 (  );
sky130_fd_sc_hd__tap_1 TAP_13727 (  );
sky130_fd_sc_hd__tap_1 TAP_13728 (  );
sky130_fd_sc_hd__tap_1 TAP_13729 (  );
sky130_fd_sc_hd__tap_1 TAP_1373 (  );
sky130_fd_sc_hd__tap_1 TAP_13730 (  );
sky130_fd_sc_hd__tap_1 TAP_13731 (  );
sky130_fd_sc_hd__tap_1 TAP_13732 (  );
sky130_fd_sc_hd__tap_1 TAP_13733 (  );
sky130_fd_sc_hd__tap_1 TAP_13734 (  );
sky130_fd_sc_hd__tap_1 TAP_13735 (  );
sky130_fd_sc_hd__tap_1 TAP_13736 (  );
sky130_fd_sc_hd__tap_1 TAP_13737 (  );
sky130_fd_sc_hd__tap_1 TAP_13738 (  );
sky130_fd_sc_hd__tap_1 TAP_13739 (  );
sky130_fd_sc_hd__tap_1 TAP_1374 (  );
sky130_fd_sc_hd__tap_1 TAP_13740 (  );
sky130_fd_sc_hd__tap_1 TAP_13741 (  );
sky130_fd_sc_hd__tap_1 TAP_13742 (  );
sky130_fd_sc_hd__tap_1 TAP_13743 (  );
sky130_fd_sc_hd__tap_1 TAP_13744 (  );
sky130_fd_sc_hd__tap_1 TAP_13745 (  );
sky130_fd_sc_hd__tap_1 TAP_13746 (  );
sky130_fd_sc_hd__tap_1 TAP_13747 (  );
sky130_fd_sc_hd__tap_1 TAP_13748 (  );
sky130_fd_sc_hd__tap_1 TAP_13749 (  );
sky130_fd_sc_hd__tap_1 TAP_1375 (  );
sky130_fd_sc_hd__tap_1 TAP_13750 (  );
sky130_fd_sc_hd__tap_1 TAP_13751 (  );
sky130_fd_sc_hd__tap_1 TAP_13752 (  );
sky130_fd_sc_hd__tap_1 TAP_13753 (  );
sky130_fd_sc_hd__tap_1 TAP_13754 (  );
sky130_fd_sc_hd__tap_1 TAP_13755 (  );
sky130_fd_sc_hd__tap_1 TAP_13756 (  );
sky130_fd_sc_hd__tap_1 TAP_13757 (  );
sky130_fd_sc_hd__tap_1 TAP_13758 (  );
sky130_fd_sc_hd__tap_1 TAP_13759 (  );
sky130_fd_sc_hd__tap_1 TAP_1376 (  );
sky130_fd_sc_hd__tap_1 TAP_13760 (  );
sky130_fd_sc_hd__tap_1 TAP_13761 (  );
sky130_fd_sc_hd__tap_1 TAP_13762 (  );
sky130_fd_sc_hd__tap_1 TAP_13763 (  );
sky130_fd_sc_hd__tap_1 TAP_13764 (  );
sky130_fd_sc_hd__tap_1 TAP_13765 (  );
sky130_fd_sc_hd__tap_1 TAP_13766 (  );
sky130_fd_sc_hd__tap_1 TAP_13767 (  );
sky130_fd_sc_hd__tap_1 TAP_13768 (  );
sky130_fd_sc_hd__tap_1 TAP_13769 (  );
sky130_fd_sc_hd__tap_1 TAP_1377 (  );
sky130_fd_sc_hd__tap_1 TAP_13770 (  );
sky130_fd_sc_hd__tap_1 TAP_13771 (  );
sky130_fd_sc_hd__tap_1 TAP_13772 (  );
sky130_fd_sc_hd__tap_1 TAP_13773 (  );
sky130_fd_sc_hd__tap_1 TAP_13774 (  );
sky130_fd_sc_hd__tap_1 TAP_13775 (  );
sky130_fd_sc_hd__tap_1 TAP_13776 (  );
sky130_fd_sc_hd__tap_1 TAP_13777 (  );
sky130_fd_sc_hd__tap_1 TAP_13778 (  );
sky130_fd_sc_hd__tap_1 TAP_13779 (  );
sky130_fd_sc_hd__tap_1 TAP_1378 (  );
sky130_fd_sc_hd__tap_1 TAP_13780 (  );
sky130_fd_sc_hd__tap_1 TAP_13781 (  );
sky130_fd_sc_hd__tap_1 TAP_13782 (  );
sky130_fd_sc_hd__tap_1 TAP_13783 (  );
sky130_fd_sc_hd__tap_1 TAP_13784 (  );
sky130_fd_sc_hd__tap_1 TAP_13785 (  );
sky130_fd_sc_hd__tap_1 TAP_13786 (  );
sky130_fd_sc_hd__tap_1 TAP_13787 (  );
sky130_fd_sc_hd__tap_1 TAP_13788 (  );
sky130_fd_sc_hd__tap_1 TAP_13789 (  );
sky130_fd_sc_hd__tap_1 TAP_1379 (  );
sky130_fd_sc_hd__tap_1 TAP_13790 (  );
sky130_fd_sc_hd__tap_1 TAP_13791 (  );
sky130_fd_sc_hd__tap_1 TAP_13792 (  );
sky130_fd_sc_hd__tap_1 TAP_13793 (  );
sky130_fd_sc_hd__tap_1 TAP_13794 (  );
sky130_fd_sc_hd__tap_1 TAP_13795 (  );
sky130_fd_sc_hd__tap_1 TAP_13796 (  );
sky130_fd_sc_hd__tap_1 TAP_13797 (  );
sky130_fd_sc_hd__tap_1 TAP_13798 (  );
sky130_fd_sc_hd__tap_1 TAP_13799 (  );
sky130_fd_sc_hd__tap_1 TAP_1380 (  );
sky130_fd_sc_hd__tap_1 TAP_13800 (  );
sky130_fd_sc_hd__tap_1 TAP_13801 (  );
sky130_fd_sc_hd__tap_1 TAP_13802 (  );
sky130_fd_sc_hd__tap_1 TAP_13803 (  );
sky130_fd_sc_hd__tap_1 TAP_13804 (  );
sky130_fd_sc_hd__tap_1 TAP_13805 (  );
sky130_fd_sc_hd__tap_1 TAP_13806 (  );
sky130_fd_sc_hd__tap_1 TAP_13807 (  );
sky130_fd_sc_hd__tap_1 TAP_13808 (  );
sky130_fd_sc_hd__tap_1 TAP_13809 (  );
sky130_fd_sc_hd__tap_1 TAP_1381 (  );
sky130_fd_sc_hd__tap_1 TAP_13810 (  );
sky130_fd_sc_hd__tap_1 TAP_13811 (  );
sky130_fd_sc_hd__tap_1 TAP_13812 (  );
sky130_fd_sc_hd__tap_1 TAP_13813 (  );
sky130_fd_sc_hd__tap_1 TAP_13814 (  );
sky130_fd_sc_hd__tap_1 TAP_13815 (  );
sky130_fd_sc_hd__tap_1 TAP_13816 (  );
sky130_fd_sc_hd__tap_1 TAP_13817 (  );
sky130_fd_sc_hd__tap_1 TAP_13818 (  );
sky130_fd_sc_hd__tap_1 TAP_13819 (  );
sky130_fd_sc_hd__tap_1 TAP_1382 (  );
sky130_fd_sc_hd__tap_1 TAP_13820 (  );
sky130_fd_sc_hd__tap_1 TAP_13821 (  );
sky130_fd_sc_hd__tap_1 TAP_13822 (  );
sky130_fd_sc_hd__tap_1 TAP_13823 (  );
sky130_fd_sc_hd__tap_1 TAP_13824 (  );
sky130_fd_sc_hd__tap_1 TAP_13825 (  );
sky130_fd_sc_hd__tap_1 TAP_13826 (  );
sky130_fd_sc_hd__tap_1 TAP_13827 (  );
sky130_fd_sc_hd__tap_1 TAP_13828 (  );
sky130_fd_sc_hd__tap_1 TAP_13829 (  );
sky130_fd_sc_hd__tap_1 TAP_1383 (  );
sky130_fd_sc_hd__tap_1 TAP_13830 (  );
sky130_fd_sc_hd__tap_1 TAP_13831 (  );
sky130_fd_sc_hd__tap_1 TAP_13832 (  );
sky130_fd_sc_hd__tap_1 TAP_13833 (  );
sky130_fd_sc_hd__tap_1 TAP_13834 (  );
sky130_fd_sc_hd__tap_1 TAP_13835 (  );
sky130_fd_sc_hd__tap_1 TAP_13836 (  );
sky130_fd_sc_hd__tap_1 TAP_13837 (  );
sky130_fd_sc_hd__tap_1 TAP_13838 (  );
sky130_fd_sc_hd__tap_1 TAP_13839 (  );
sky130_fd_sc_hd__tap_1 TAP_1384 (  );
sky130_fd_sc_hd__tap_1 TAP_13840 (  );
sky130_fd_sc_hd__tap_1 TAP_13841 (  );
sky130_fd_sc_hd__tap_1 TAP_13842 (  );
sky130_fd_sc_hd__tap_1 TAP_13843 (  );
sky130_fd_sc_hd__tap_1 TAP_13844 (  );
sky130_fd_sc_hd__tap_1 TAP_13845 (  );
sky130_fd_sc_hd__tap_1 TAP_13846 (  );
sky130_fd_sc_hd__tap_1 TAP_13847 (  );
sky130_fd_sc_hd__tap_1 TAP_13848 (  );
sky130_fd_sc_hd__tap_1 TAP_13849 (  );
sky130_fd_sc_hd__tap_1 TAP_1385 (  );
sky130_fd_sc_hd__tap_1 TAP_13850 (  );
sky130_fd_sc_hd__tap_1 TAP_13851 (  );
sky130_fd_sc_hd__tap_1 TAP_13852 (  );
sky130_fd_sc_hd__tap_1 TAP_13853 (  );
sky130_fd_sc_hd__tap_1 TAP_13854 (  );
sky130_fd_sc_hd__tap_1 TAP_13855 (  );
sky130_fd_sc_hd__tap_1 TAP_13856 (  );
sky130_fd_sc_hd__tap_1 TAP_13857 (  );
sky130_fd_sc_hd__tap_1 TAP_13858 (  );
sky130_fd_sc_hd__tap_1 TAP_13859 (  );
sky130_fd_sc_hd__tap_1 TAP_1386 (  );
sky130_fd_sc_hd__tap_1 TAP_13860 (  );
sky130_fd_sc_hd__tap_1 TAP_13861 (  );
sky130_fd_sc_hd__tap_1 TAP_13862 (  );
sky130_fd_sc_hd__tap_1 TAP_13863 (  );
sky130_fd_sc_hd__tap_1 TAP_13864 (  );
sky130_fd_sc_hd__tap_1 TAP_13865 (  );
sky130_fd_sc_hd__tap_1 TAP_13866 (  );
sky130_fd_sc_hd__tap_1 TAP_13867 (  );
sky130_fd_sc_hd__tap_1 TAP_13868 (  );
sky130_fd_sc_hd__tap_1 TAP_13869 (  );
sky130_fd_sc_hd__tap_1 TAP_1387 (  );
sky130_fd_sc_hd__tap_1 TAP_13870 (  );
sky130_fd_sc_hd__tap_1 TAP_13871 (  );
sky130_fd_sc_hd__tap_1 TAP_13872 (  );
sky130_fd_sc_hd__tap_1 TAP_13873 (  );
sky130_fd_sc_hd__tap_1 TAP_13874 (  );
sky130_fd_sc_hd__tap_1 TAP_13875 (  );
sky130_fd_sc_hd__tap_1 TAP_13876 (  );
sky130_fd_sc_hd__tap_1 TAP_13877 (  );
sky130_fd_sc_hd__tap_1 TAP_13878 (  );
sky130_fd_sc_hd__tap_1 TAP_13879 (  );
sky130_fd_sc_hd__tap_1 TAP_1388 (  );
sky130_fd_sc_hd__tap_1 TAP_13880 (  );
sky130_fd_sc_hd__tap_1 TAP_13881 (  );
sky130_fd_sc_hd__tap_1 TAP_13882 (  );
sky130_fd_sc_hd__tap_1 TAP_13883 (  );
sky130_fd_sc_hd__tap_1 TAP_13884 (  );
sky130_fd_sc_hd__tap_1 TAP_13885 (  );
sky130_fd_sc_hd__tap_1 TAP_13886 (  );
sky130_fd_sc_hd__tap_1 TAP_13887 (  );
sky130_fd_sc_hd__tap_1 TAP_13888 (  );
sky130_fd_sc_hd__tap_1 TAP_13889 (  );
sky130_fd_sc_hd__tap_1 TAP_1389 (  );
sky130_fd_sc_hd__tap_1 TAP_13890 (  );
sky130_fd_sc_hd__tap_1 TAP_13891 (  );
sky130_fd_sc_hd__tap_1 TAP_13892 (  );
sky130_fd_sc_hd__tap_1 TAP_13893 (  );
sky130_fd_sc_hd__tap_1 TAP_13894 (  );
sky130_fd_sc_hd__tap_1 TAP_13895 (  );
sky130_fd_sc_hd__tap_1 TAP_13896 (  );
sky130_fd_sc_hd__tap_1 TAP_13897 (  );
sky130_fd_sc_hd__tap_1 TAP_13898 (  );
sky130_fd_sc_hd__tap_1 TAP_13899 (  );
sky130_fd_sc_hd__tap_1 TAP_1390 (  );
sky130_fd_sc_hd__tap_1 TAP_13900 (  );
sky130_fd_sc_hd__tap_1 TAP_13901 (  );
sky130_fd_sc_hd__tap_1 TAP_13902 (  );
sky130_fd_sc_hd__tap_1 TAP_13903 (  );
sky130_fd_sc_hd__tap_1 TAP_13904 (  );
sky130_fd_sc_hd__tap_1 TAP_13905 (  );
sky130_fd_sc_hd__tap_1 TAP_13906 (  );
sky130_fd_sc_hd__tap_1 TAP_13907 (  );
sky130_fd_sc_hd__tap_1 TAP_13908 (  );
sky130_fd_sc_hd__tap_1 TAP_13909 (  );
sky130_fd_sc_hd__tap_1 TAP_1391 (  );
sky130_fd_sc_hd__tap_1 TAP_13910 (  );
sky130_fd_sc_hd__tap_1 TAP_13911 (  );
sky130_fd_sc_hd__tap_1 TAP_13912 (  );
sky130_fd_sc_hd__tap_1 TAP_13913 (  );
sky130_fd_sc_hd__tap_1 TAP_13914 (  );
sky130_fd_sc_hd__tap_1 TAP_13915 (  );
sky130_fd_sc_hd__tap_1 TAP_13916 (  );
sky130_fd_sc_hd__tap_1 TAP_13917 (  );
sky130_fd_sc_hd__tap_1 TAP_13918 (  );
sky130_fd_sc_hd__tap_1 TAP_13919 (  );
sky130_fd_sc_hd__tap_1 TAP_1392 (  );
sky130_fd_sc_hd__tap_1 TAP_13920 (  );
sky130_fd_sc_hd__tap_1 TAP_13921 (  );
sky130_fd_sc_hd__tap_1 TAP_13922 (  );
sky130_fd_sc_hd__tap_1 TAP_13923 (  );
sky130_fd_sc_hd__tap_1 TAP_13924 (  );
sky130_fd_sc_hd__tap_1 TAP_13925 (  );
sky130_fd_sc_hd__tap_1 TAP_13926 (  );
sky130_fd_sc_hd__tap_1 TAP_13927 (  );
sky130_fd_sc_hd__tap_1 TAP_13928 (  );
sky130_fd_sc_hd__tap_1 TAP_13929 (  );
sky130_fd_sc_hd__tap_1 TAP_1393 (  );
sky130_fd_sc_hd__tap_1 TAP_13930 (  );
sky130_fd_sc_hd__tap_1 TAP_13931 (  );
sky130_fd_sc_hd__tap_1 TAP_13932 (  );
sky130_fd_sc_hd__tap_1 TAP_13933 (  );
sky130_fd_sc_hd__tap_1 TAP_13934 (  );
sky130_fd_sc_hd__tap_1 TAP_13935 (  );
sky130_fd_sc_hd__tap_1 TAP_13936 (  );
sky130_fd_sc_hd__tap_1 TAP_13937 (  );
sky130_fd_sc_hd__tap_1 TAP_13938 (  );
sky130_fd_sc_hd__tap_1 TAP_13939 (  );
sky130_fd_sc_hd__tap_1 TAP_1394 (  );
sky130_fd_sc_hd__tap_1 TAP_13940 (  );
sky130_fd_sc_hd__tap_1 TAP_13941 (  );
sky130_fd_sc_hd__tap_1 TAP_13942 (  );
sky130_fd_sc_hd__tap_1 TAP_13943 (  );
sky130_fd_sc_hd__tap_1 TAP_13944 (  );
sky130_fd_sc_hd__tap_1 TAP_13945 (  );
sky130_fd_sc_hd__tap_1 TAP_13946 (  );
sky130_fd_sc_hd__tap_1 TAP_13947 (  );
sky130_fd_sc_hd__tap_1 TAP_13948 (  );
sky130_fd_sc_hd__tap_1 TAP_13949 (  );
sky130_fd_sc_hd__tap_1 TAP_1395 (  );
sky130_fd_sc_hd__tap_1 TAP_13950 (  );
sky130_fd_sc_hd__tap_1 TAP_13951 (  );
sky130_fd_sc_hd__tap_1 TAP_13952 (  );
sky130_fd_sc_hd__tap_1 TAP_13953 (  );
sky130_fd_sc_hd__tap_1 TAP_13954 (  );
sky130_fd_sc_hd__tap_1 TAP_13955 (  );
sky130_fd_sc_hd__tap_1 TAP_13956 (  );
sky130_fd_sc_hd__tap_1 TAP_13957 (  );
sky130_fd_sc_hd__tap_1 TAP_13958 (  );
sky130_fd_sc_hd__tap_1 TAP_13959 (  );
sky130_fd_sc_hd__tap_1 TAP_1396 (  );
sky130_fd_sc_hd__tap_1 TAP_13960 (  );
sky130_fd_sc_hd__tap_1 TAP_13961 (  );
sky130_fd_sc_hd__tap_1 TAP_13962 (  );
sky130_fd_sc_hd__tap_1 TAP_13963 (  );
sky130_fd_sc_hd__tap_1 TAP_13964 (  );
sky130_fd_sc_hd__tap_1 TAP_13965 (  );
sky130_fd_sc_hd__tap_1 TAP_13966 (  );
sky130_fd_sc_hd__tap_1 TAP_13967 (  );
sky130_fd_sc_hd__tap_1 TAP_13968 (  );
sky130_fd_sc_hd__tap_1 TAP_13969 (  );
sky130_fd_sc_hd__tap_1 TAP_1397 (  );
sky130_fd_sc_hd__tap_1 TAP_13970 (  );
sky130_fd_sc_hd__tap_1 TAP_13971 (  );
sky130_fd_sc_hd__tap_1 TAP_13972 (  );
sky130_fd_sc_hd__tap_1 TAP_13973 (  );
sky130_fd_sc_hd__tap_1 TAP_13974 (  );
sky130_fd_sc_hd__tap_1 TAP_13975 (  );
sky130_fd_sc_hd__tap_1 TAP_13976 (  );
sky130_fd_sc_hd__tap_1 TAP_13977 (  );
sky130_fd_sc_hd__tap_1 TAP_13978 (  );
sky130_fd_sc_hd__tap_1 TAP_13979 (  );
sky130_fd_sc_hd__tap_1 TAP_1398 (  );
sky130_fd_sc_hd__tap_1 TAP_13980 (  );
sky130_fd_sc_hd__tap_1 TAP_13981 (  );
sky130_fd_sc_hd__tap_1 TAP_13982 (  );
sky130_fd_sc_hd__tap_1 TAP_13983 (  );
sky130_fd_sc_hd__tap_1 TAP_13984 (  );
sky130_fd_sc_hd__tap_1 TAP_13985 (  );
sky130_fd_sc_hd__tap_1 TAP_13986 (  );
sky130_fd_sc_hd__tap_1 TAP_13987 (  );
sky130_fd_sc_hd__tap_1 TAP_13988 (  );
sky130_fd_sc_hd__tap_1 TAP_13989 (  );
sky130_fd_sc_hd__tap_1 TAP_1399 (  );
sky130_fd_sc_hd__tap_1 TAP_13990 (  );
sky130_fd_sc_hd__tap_1 TAP_13991 (  );
sky130_fd_sc_hd__tap_1 TAP_13992 (  );
sky130_fd_sc_hd__tap_1 TAP_13993 (  );
sky130_fd_sc_hd__tap_1 TAP_13994 (  );
sky130_fd_sc_hd__tap_1 TAP_13995 (  );
sky130_fd_sc_hd__tap_1 TAP_13996 (  );
sky130_fd_sc_hd__tap_1 TAP_13997 (  );
sky130_fd_sc_hd__tap_1 TAP_13998 (  );
sky130_fd_sc_hd__tap_1 TAP_13999 (  );
sky130_fd_sc_hd__tap_1 TAP_1400 (  );
sky130_fd_sc_hd__tap_1 TAP_14000 (  );
sky130_fd_sc_hd__tap_1 TAP_14001 (  );
sky130_fd_sc_hd__tap_1 TAP_14002 (  );
sky130_fd_sc_hd__tap_1 TAP_14003 (  );
sky130_fd_sc_hd__tap_1 TAP_14004 (  );
sky130_fd_sc_hd__tap_1 TAP_14005 (  );
sky130_fd_sc_hd__tap_1 TAP_14006 (  );
sky130_fd_sc_hd__tap_1 TAP_14007 (  );
sky130_fd_sc_hd__tap_1 TAP_14008 (  );
sky130_fd_sc_hd__tap_1 TAP_14009 (  );
sky130_fd_sc_hd__tap_1 TAP_1401 (  );
sky130_fd_sc_hd__tap_1 TAP_14010 (  );
sky130_fd_sc_hd__tap_1 TAP_14011 (  );
sky130_fd_sc_hd__tap_1 TAP_14012 (  );
sky130_fd_sc_hd__tap_1 TAP_14013 (  );
sky130_fd_sc_hd__tap_1 TAP_14014 (  );
sky130_fd_sc_hd__tap_1 TAP_14015 (  );
sky130_fd_sc_hd__tap_1 TAP_14016 (  );
sky130_fd_sc_hd__tap_1 TAP_14017 (  );
sky130_fd_sc_hd__tap_1 TAP_14018 (  );
sky130_fd_sc_hd__tap_1 TAP_14019 (  );
sky130_fd_sc_hd__tap_1 TAP_1402 (  );
sky130_fd_sc_hd__tap_1 TAP_14020 (  );
sky130_fd_sc_hd__tap_1 TAP_14021 (  );
sky130_fd_sc_hd__tap_1 TAP_14022 (  );
sky130_fd_sc_hd__tap_1 TAP_14023 (  );
sky130_fd_sc_hd__tap_1 TAP_14024 (  );
sky130_fd_sc_hd__tap_1 TAP_14025 (  );
sky130_fd_sc_hd__tap_1 TAP_14026 (  );
sky130_fd_sc_hd__tap_1 TAP_14027 (  );
sky130_fd_sc_hd__tap_1 TAP_14028 (  );
sky130_fd_sc_hd__tap_1 TAP_14029 (  );
sky130_fd_sc_hd__tap_1 TAP_1403 (  );
sky130_fd_sc_hd__tap_1 TAP_14030 (  );
sky130_fd_sc_hd__tap_1 TAP_14031 (  );
sky130_fd_sc_hd__tap_1 TAP_14032 (  );
sky130_fd_sc_hd__tap_1 TAP_14033 (  );
sky130_fd_sc_hd__tap_1 TAP_14034 (  );
sky130_fd_sc_hd__tap_1 TAP_14035 (  );
sky130_fd_sc_hd__tap_1 TAP_14036 (  );
sky130_fd_sc_hd__tap_1 TAP_14037 (  );
sky130_fd_sc_hd__tap_1 TAP_14038 (  );
sky130_fd_sc_hd__tap_1 TAP_14039 (  );
sky130_fd_sc_hd__tap_1 TAP_1404 (  );
sky130_fd_sc_hd__tap_1 TAP_14040 (  );
sky130_fd_sc_hd__tap_1 TAP_14041 (  );
sky130_fd_sc_hd__tap_1 TAP_14042 (  );
sky130_fd_sc_hd__tap_1 TAP_14043 (  );
sky130_fd_sc_hd__tap_1 TAP_14044 (  );
sky130_fd_sc_hd__tap_1 TAP_14045 (  );
sky130_fd_sc_hd__tap_1 TAP_14046 (  );
sky130_fd_sc_hd__tap_1 TAP_14047 (  );
sky130_fd_sc_hd__tap_1 TAP_14048 (  );
sky130_fd_sc_hd__tap_1 TAP_14049 (  );
sky130_fd_sc_hd__tap_1 TAP_1405 (  );
sky130_fd_sc_hd__tap_1 TAP_14050 (  );
sky130_fd_sc_hd__tap_1 TAP_14051 (  );
sky130_fd_sc_hd__tap_1 TAP_14052 (  );
sky130_fd_sc_hd__tap_1 TAP_14053 (  );
sky130_fd_sc_hd__tap_1 TAP_14054 (  );
sky130_fd_sc_hd__tap_1 TAP_14055 (  );
sky130_fd_sc_hd__tap_1 TAP_14056 (  );
sky130_fd_sc_hd__tap_1 TAP_14057 (  );
sky130_fd_sc_hd__tap_1 TAP_14058 (  );
sky130_fd_sc_hd__tap_1 TAP_14059 (  );
sky130_fd_sc_hd__tap_1 TAP_1406 (  );
sky130_fd_sc_hd__tap_1 TAP_14060 (  );
sky130_fd_sc_hd__tap_1 TAP_14061 (  );
sky130_fd_sc_hd__tap_1 TAP_14062 (  );
sky130_fd_sc_hd__tap_1 TAP_14063 (  );
sky130_fd_sc_hd__tap_1 TAP_14064 (  );
sky130_fd_sc_hd__tap_1 TAP_14065 (  );
sky130_fd_sc_hd__tap_1 TAP_14066 (  );
sky130_fd_sc_hd__tap_1 TAP_14067 (  );
sky130_fd_sc_hd__tap_1 TAP_14068 (  );
sky130_fd_sc_hd__tap_1 TAP_14069 (  );
sky130_fd_sc_hd__tap_1 TAP_1407 (  );
sky130_fd_sc_hd__tap_1 TAP_14070 (  );
sky130_fd_sc_hd__tap_1 TAP_14071 (  );
sky130_fd_sc_hd__tap_1 TAP_14072 (  );
sky130_fd_sc_hd__tap_1 TAP_14073 (  );
sky130_fd_sc_hd__tap_1 TAP_14074 (  );
sky130_fd_sc_hd__tap_1 TAP_14075 (  );
sky130_fd_sc_hd__tap_1 TAP_14076 (  );
sky130_fd_sc_hd__tap_1 TAP_14077 (  );
sky130_fd_sc_hd__tap_1 TAP_14078 (  );
sky130_fd_sc_hd__tap_1 TAP_14079 (  );
sky130_fd_sc_hd__tap_1 TAP_1408 (  );
sky130_fd_sc_hd__tap_1 TAP_14080 (  );
sky130_fd_sc_hd__tap_1 TAP_14081 (  );
sky130_fd_sc_hd__tap_1 TAP_14082 (  );
sky130_fd_sc_hd__tap_1 TAP_14083 (  );
sky130_fd_sc_hd__tap_1 TAP_14084 (  );
sky130_fd_sc_hd__tap_1 TAP_14085 (  );
sky130_fd_sc_hd__tap_1 TAP_14086 (  );
sky130_fd_sc_hd__tap_1 TAP_14087 (  );
sky130_fd_sc_hd__tap_1 TAP_14088 (  );
sky130_fd_sc_hd__tap_1 TAP_14089 (  );
sky130_fd_sc_hd__tap_1 TAP_1409 (  );
sky130_fd_sc_hd__tap_1 TAP_14090 (  );
sky130_fd_sc_hd__tap_1 TAP_14091 (  );
sky130_fd_sc_hd__tap_1 TAP_14092 (  );
sky130_fd_sc_hd__tap_1 TAP_14093 (  );
sky130_fd_sc_hd__tap_1 TAP_14094 (  );
sky130_fd_sc_hd__tap_1 TAP_14095 (  );
sky130_fd_sc_hd__tap_1 TAP_14096 (  );
sky130_fd_sc_hd__tap_1 TAP_14097 (  );
sky130_fd_sc_hd__tap_1 TAP_14098 (  );
sky130_fd_sc_hd__tap_1 TAP_14099 (  );
sky130_fd_sc_hd__tap_1 TAP_1410 (  );
sky130_fd_sc_hd__tap_1 TAP_14100 (  );
sky130_fd_sc_hd__tap_1 TAP_14101 (  );
sky130_fd_sc_hd__tap_1 TAP_14102 (  );
sky130_fd_sc_hd__tap_1 TAP_14103 (  );
sky130_fd_sc_hd__tap_1 TAP_14104 (  );
sky130_fd_sc_hd__tap_1 TAP_14105 (  );
sky130_fd_sc_hd__tap_1 TAP_14106 (  );
sky130_fd_sc_hd__tap_1 TAP_14107 (  );
sky130_fd_sc_hd__tap_1 TAP_14108 (  );
sky130_fd_sc_hd__tap_1 TAP_14109 (  );
sky130_fd_sc_hd__tap_1 TAP_1411 (  );
sky130_fd_sc_hd__tap_1 TAP_14110 (  );
sky130_fd_sc_hd__tap_1 TAP_14111 (  );
sky130_fd_sc_hd__tap_1 TAP_14112 (  );
sky130_fd_sc_hd__tap_1 TAP_14113 (  );
sky130_fd_sc_hd__tap_1 TAP_14114 (  );
sky130_fd_sc_hd__tap_1 TAP_14115 (  );
sky130_fd_sc_hd__tap_1 TAP_14116 (  );
sky130_fd_sc_hd__tap_1 TAP_14117 (  );
sky130_fd_sc_hd__tap_1 TAP_14118 (  );
sky130_fd_sc_hd__tap_1 TAP_14119 (  );
sky130_fd_sc_hd__tap_1 TAP_1412 (  );
sky130_fd_sc_hd__tap_1 TAP_14120 (  );
sky130_fd_sc_hd__tap_1 TAP_14121 (  );
sky130_fd_sc_hd__tap_1 TAP_14122 (  );
sky130_fd_sc_hd__tap_1 TAP_14123 (  );
sky130_fd_sc_hd__tap_1 TAP_14124 (  );
sky130_fd_sc_hd__tap_1 TAP_14125 (  );
sky130_fd_sc_hd__tap_1 TAP_14126 (  );
sky130_fd_sc_hd__tap_1 TAP_14127 (  );
sky130_fd_sc_hd__tap_1 TAP_14128 (  );
sky130_fd_sc_hd__tap_1 TAP_14129 (  );
sky130_fd_sc_hd__tap_1 TAP_1413 (  );
sky130_fd_sc_hd__tap_1 TAP_14130 (  );
sky130_fd_sc_hd__tap_1 TAP_14131 (  );
sky130_fd_sc_hd__tap_1 TAP_14132 (  );
sky130_fd_sc_hd__tap_1 TAP_14133 (  );
sky130_fd_sc_hd__tap_1 TAP_14134 (  );
sky130_fd_sc_hd__tap_1 TAP_14135 (  );
sky130_fd_sc_hd__tap_1 TAP_14136 (  );
sky130_fd_sc_hd__tap_1 TAP_14137 (  );
sky130_fd_sc_hd__tap_1 TAP_14138 (  );
sky130_fd_sc_hd__tap_1 TAP_14139 (  );
sky130_fd_sc_hd__tap_1 TAP_1414 (  );
sky130_fd_sc_hd__tap_1 TAP_14140 (  );
sky130_fd_sc_hd__tap_1 TAP_14141 (  );
sky130_fd_sc_hd__tap_1 TAP_14142 (  );
sky130_fd_sc_hd__tap_1 TAP_14143 (  );
sky130_fd_sc_hd__tap_1 TAP_14144 (  );
sky130_fd_sc_hd__tap_1 TAP_14145 (  );
sky130_fd_sc_hd__tap_1 TAP_14146 (  );
sky130_fd_sc_hd__tap_1 TAP_14147 (  );
sky130_fd_sc_hd__tap_1 TAP_14148 (  );
sky130_fd_sc_hd__tap_1 TAP_14149 (  );
sky130_fd_sc_hd__tap_1 TAP_1415 (  );
sky130_fd_sc_hd__tap_1 TAP_14150 (  );
sky130_fd_sc_hd__tap_1 TAP_14151 (  );
sky130_fd_sc_hd__tap_1 TAP_14152 (  );
sky130_fd_sc_hd__tap_1 TAP_14153 (  );
sky130_fd_sc_hd__tap_1 TAP_14154 (  );
sky130_fd_sc_hd__tap_1 TAP_14155 (  );
sky130_fd_sc_hd__tap_1 TAP_14156 (  );
sky130_fd_sc_hd__tap_1 TAP_14157 (  );
sky130_fd_sc_hd__tap_1 TAP_14158 (  );
sky130_fd_sc_hd__tap_1 TAP_14159 (  );
sky130_fd_sc_hd__tap_1 TAP_1416 (  );
sky130_fd_sc_hd__tap_1 TAP_14160 (  );
sky130_fd_sc_hd__tap_1 TAP_14161 (  );
sky130_fd_sc_hd__tap_1 TAP_14162 (  );
sky130_fd_sc_hd__tap_1 TAP_14163 (  );
sky130_fd_sc_hd__tap_1 TAP_14164 (  );
sky130_fd_sc_hd__tap_1 TAP_14165 (  );
sky130_fd_sc_hd__tap_1 TAP_14166 (  );
sky130_fd_sc_hd__tap_1 TAP_14167 (  );
sky130_fd_sc_hd__tap_1 TAP_14168 (  );
sky130_fd_sc_hd__tap_1 TAP_14169 (  );
sky130_fd_sc_hd__tap_1 TAP_1417 (  );
sky130_fd_sc_hd__tap_1 TAP_14170 (  );
sky130_fd_sc_hd__tap_1 TAP_14171 (  );
sky130_fd_sc_hd__tap_1 TAP_14172 (  );
sky130_fd_sc_hd__tap_1 TAP_14173 (  );
sky130_fd_sc_hd__tap_1 TAP_14174 (  );
sky130_fd_sc_hd__tap_1 TAP_14175 (  );
sky130_fd_sc_hd__tap_1 TAP_14176 (  );
sky130_fd_sc_hd__tap_1 TAP_14177 (  );
sky130_fd_sc_hd__tap_1 TAP_14178 (  );
sky130_fd_sc_hd__tap_1 TAP_14179 (  );
sky130_fd_sc_hd__tap_1 TAP_1418 (  );
sky130_fd_sc_hd__tap_1 TAP_14180 (  );
sky130_fd_sc_hd__tap_1 TAP_14181 (  );
sky130_fd_sc_hd__tap_1 TAP_14182 (  );
sky130_fd_sc_hd__tap_1 TAP_14183 (  );
sky130_fd_sc_hd__tap_1 TAP_14184 (  );
sky130_fd_sc_hd__tap_1 TAP_14185 (  );
sky130_fd_sc_hd__tap_1 TAP_14186 (  );
sky130_fd_sc_hd__tap_1 TAP_14187 (  );
sky130_fd_sc_hd__tap_1 TAP_14188 (  );
sky130_fd_sc_hd__tap_1 TAP_14189 (  );
sky130_fd_sc_hd__tap_1 TAP_1419 (  );
sky130_fd_sc_hd__tap_1 TAP_14190 (  );
sky130_fd_sc_hd__tap_1 TAP_14191 (  );
sky130_fd_sc_hd__tap_1 TAP_14192 (  );
sky130_fd_sc_hd__tap_1 TAP_14193 (  );
sky130_fd_sc_hd__tap_1 TAP_14194 (  );
sky130_fd_sc_hd__tap_1 TAP_14195 (  );
sky130_fd_sc_hd__tap_1 TAP_14196 (  );
sky130_fd_sc_hd__tap_1 TAP_14197 (  );
sky130_fd_sc_hd__tap_1 TAP_14198 (  );
sky130_fd_sc_hd__tap_1 TAP_14199 (  );
sky130_fd_sc_hd__tap_1 TAP_1420 (  );
sky130_fd_sc_hd__tap_1 TAP_14200 (  );
sky130_fd_sc_hd__tap_1 TAP_14201 (  );
sky130_fd_sc_hd__tap_1 TAP_14202 (  );
sky130_fd_sc_hd__tap_1 TAP_14203 (  );
sky130_fd_sc_hd__tap_1 TAP_14204 (  );
sky130_fd_sc_hd__tap_1 TAP_14205 (  );
sky130_fd_sc_hd__tap_1 TAP_14206 (  );
sky130_fd_sc_hd__tap_1 TAP_14207 (  );
sky130_fd_sc_hd__tap_1 TAP_14208 (  );
sky130_fd_sc_hd__tap_1 TAP_14209 (  );
sky130_fd_sc_hd__tap_1 TAP_1421 (  );
sky130_fd_sc_hd__tap_1 TAP_14210 (  );
sky130_fd_sc_hd__tap_1 TAP_14211 (  );
sky130_fd_sc_hd__tap_1 TAP_14212 (  );
sky130_fd_sc_hd__tap_1 TAP_14213 (  );
sky130_fd_sc_hd__tap_1 TAP_14214 (  );
sky130_fd_sc_hd__tap_1 TAP_14215 (  );
sky130_fd_sc_hd__tap_1 TAP_14216 (  );
sky130_fd_sc_hd__tap_1 TAP_14217 (  );
sky130_fd_sc_hd__tap_1 TAP_14218 (  );
sky130_fd_sc_hd__tap_1 TAP_14219 (  );
sky130_fd_sc_hd__tap_1 TAP_1422 (  );
sky130_fd_sc_hd__tap_1 TAP_14220 (  );
sky130_fd_sc_hd__tap_1 TAP_14221 (  );
sky130_fd_sc_hd__tap_1 TAP_14222 (  );
sky130_fd_sc_hd__tap_1 TAP_14223 (  );
sky130_fd_sc_hd__tap_1 TAP_14224 (  );
sky130_fd_sc_hd__tap_1 TAP_14225 (  );
sky130_fd_sc_hd__tap_1 TAP_14226 (  );
sky130_fd_sc_hd__tap_1 TAP_14227 (  );
sky130_fd_sc_hd__tap_1 TAP_14228 (  );
sky130_fd_sc_hd__tap_1 TAP_14229 (  );
sky130_fd_sc_hd__tap_1 TAP_1423 (  );
sky130_fd_sc_hd__tap_1 TAP_14230 (  );
sky130_fd_sc_hd__tap_1 TAP_14231 (  );
sky130_fd_sc_hd__tap_1 TAP_14232 (  );
sky130_fd_sc_hd__tap_1 TAP_14233 (  );
sky130_fd_sc_hd__tap_1 TAP_14234 (  );
sky130_fd_sc_hd__tap_1 TAP_14235 (  );
sky130_fd_sc_hd__tap_1 TAP_14236 (  );
sky130_fd_sc_hd__tap_1 TAP_14237 (  );
sky130_fd_sc_hd__tap_1 TAP_14238 (  );
sky130_fd_sc_hd__tap_1 TAP_14239 (  );
sky130_fd_sc_hd__tap_1 TAP_1424 (  );
sky130_fd_sc_hd__tap_1 TAP_14240 (  );
sky130_fd_sc_hd__tap_1 TAP_14241 (  );
sky130_fd_sc_hd__tap_1 TAP_14242 (  );
sky130_fd_sc_hd__tap_1 TAP_14243 (  );
sky130_fd_sc_hd__tap_1 TAP_14244 (  );
sky130_fd_sc_hd__tap_1 TAP_14245 (  );
sky130_fd_sc_hd__tap_1 TAP_14246 (  );
sky130_fd_sc_hd__tap_1 TAP_14247 (  );
sky130_fd_sc_hd__tap_1 TAP_14248 (  );
sky130_fd_sc_hd__tap_1 TAP_14249 (  );
sky130_fd_sc_hd__tap_1 TAP_1425 (  );
sky130_fd_sc_hd__tap_1 TAP_14250 (  );
sky130_fd_sc_hd__tap_1 TAP_14251 (  );
sky130_fd_sc_hd__tap_1 TAP_14252 (  );
sky130_fd_sc_hd__tap_1 TAP_14253 (  );
sky130_fd_sc_hd__tap_1 TAP_14254 (  );
sky130_fd_sc_hd__tap_1 TAP_14255 (  );
sky130_fd_sc_hd__tap_1 TAP_14256 (  );
sky130_fd_sc_hd__tap_1 TAP_14257 (  );
sky130_fd_sc_hd__tap_1 TAP_14258 (  );
sky130_fd_sc_hd__tap_1 TAP_14259 (  );
sky130_fd_sc_hd__tap_1 TAP_1426 (  );
sky130_fd_sc_hd__tap_1 TAP_14260 (  );
sky130_fd_sc_hd__tap_1 TAP_14261 (  );
sky130_fd_sc_hd__tap_1 TAP_14262 (  );
sky130_fd_sc_hd__tap_1 TAP_14263 (  );
sky130_fd_sc_hd__tap_1 TAP_14264 (  );
sky130_fd_sc_hd__tap_1 TAP_14265 (  );
sky130_fd_sc_hd__tap_1 TAP_14266 (  );
sky130_fd_sc_hd__tap_1 TAP_14267 (  );
sky130_fd_sc_hd__tap_1 TAP_14268 (  );
sky130_fd_sc_hd__tap_1 TAP_14269 (  );
sky130_fd_sc_hd__tap_1 TAP_1427 (  );
sky130_fd_sc_hd__tap_1 TAP_14270 (  );
sky130_fd_sc_hd__tap_1 TAP_14271 (  );
sky130_fd_sc_hd__tap_1 TAP_14272 (  );
sky130_fd_sc_hd__tap_1 TAP_14273 (  );
sky130_fd_sc_hd__tap_1 TAP_14274 (  );
sky130_fd_sc_hd__tap_1 TAP_14275 (  );
sky130_fd_sc_hd__tap_1 TAP_14276 (  );
sky130_fd_sc_hd__tap_1 TAP_14277 (  );
sky130_fd_sc_hd__tap_1 TAP_14278 (  );
sky130_fd_sc_hd__tap_1 TAP_14279 (  );
sky130_fd_sc_hd__tap_1 TAP_1428 (  );
sky130_fd_sc_hd__tap_1 TAP_14280 (  );
sky130_fd_sc_hd__tap_1 TAP_14281 (  );
sky130_fd_sc_hd__tap_1 TAP_14282 (  );
sky130_fd_sc_hd__tap_1 TAP_14283 (  );
sky130_fd_sc_hd__tap_1 TAP_14284 (  );
sky130_fd_sc_hd__tap_1 TAP_14285 (  );
sky130_fd_sc_hd__tap_1 TAP_14286 (  );
sky130_fd_sc_hd__tap_1 TAP_14287 (  );
sky130_fd_sc_hd__tap_1 TAP_14288 (  );
sky130_fd_sc_hd__tap_1 TAP_14289 (  );
sky130_fd_sc_hd__tap_1 TAP_1429 (  );
sky130_fd_sc_hd__tap_1 TAP_14290 (  );
sky130_fd_sc_hd__tap_1 TAP_14291 (  );
sky130_fd_sc_hd__tap_1 TAP_14292 (  );
sky130_fd_sc_hd__tap_1 TAP_14293 (  );
sky130_fd_sc_hd__tap_1 TAP_14294 (  );
sky130_fd_sc_hd__tap_1 TAP_14295 (  );
sky130_fd_sc_hd__tap_1 TAP_14296 (  );
sky130_fd_sc_hd__tap_1 TAP_14297 (  );
sky130_fd_sc_hd__tap_1 TAP_14298 (  );
sky130_fd_sc_hd__tap_1 TAP_14299 (  );
sky130_fd_sc_hd__tap_1 TAP_1430 (  );
sky130_fd_sc_hd__tap_1 TAP_14300 (  );
sky130_fd_sc_hd__tap_1 TAP_14301 (  );
sky130_fd_sc_hd__tap_1 TAP_14302 (  );
sky130_fd_sc_hd__tap_1 TAP_14303 (  );
sky130_fd_sc_hd__tap_1 TAP_14304 (  );
sky130_fd_sc_hd__tap_1 TAP_14305 (  );
sky130_fd_sc_hd__tap_1 TAP_14306 (  );
sky130_fd_sc_hd__tap_1 TAP_14307 (  );
sky130_fd_sc_hd__tap_1 TAP_14308 (  );
sky130_fd_sc_hd__tap_1 TAP_14309 (  );
sky130_fd_sc_hd__tap_1 TAP_1431 (  );
sky130_fd_sc_hd__tap_1 TAP_14310 (  );
sky130_fd_sc_hd__tap_1 TAP_14311 (  );
sky130_fd_sc_hd__tap_1 TAP_14312 (  );
sky130_fd_sc_hd__tap_1 TAP_14313 (  );
sky130_fd_sc_hd__tap_1 TAP_14314 (  );
sky130_fd_sc_hd__tap_1 TAP_14315 (  );
sky130_fd_sc_hd__tap_1 TAP_14316 (  );
sky130_fd_sc_hd__tap_1 TAP_14317 (  );
sky130_fd_sc_hd__tap_1 TAP_14318 (  );
sky130_fd_sc_hd__tap_1 TAP_14319 (  );
sky130_fd_sc_hd__tap_1 TAP_1432 (  );
sky130_fd_sc_hd__tap_1 TAP_14320 (  );
sky130_fd_sc_hd__tap_1 TAP_14321 (  );
sky130_fd_sc_hd__tap_1 TAP_14322 (  );
sky130_fd_sc_hd__tap_1 TAP_14323 (  );
sky130_fd_sc_hd__tap_1 TAP_14324 (  );
sky130_fd_sc_hd__tap_1 TAP_14325 (  );
sky130_fd_sc_hd__tap_1 TAP_14326 (  );
sky130_fd_sc_hd__tap_1 TAP_14327 (  );
sky130_fd_sc_hd__tap_1 TAP_14328 (  );
sky130_fd_sc_hd__tap_1 TAP_14329 (  );
sky130_fd_sc_hd__tap_1 TAP_1433 (  );
sky130_fd_sc_hd__tap_1 TAP_14330 (  );
sky130_fd_sc_hd__tap_1 TAP_14331 (  );
sky130_fd_sc_hd__tap_1 TAP_14332 (  );
sky130_fd_sc_hd__tap_1 TAP_14333 (  );
sky130_fd_sc_hd__tap_1 TAP_14334 (  );
sky130_fd_sc_hd__tap_1 TAP_14335 (  );
sky130_fd_sc_hd__tap_1 TAP_14336 (  );
sky130_fd_sc_hd__tap_1 TAP_14337 (  );
sky130_fd_sc_hd__tap_1 TAP_14338 (  );
sky130_fd_sc_hd__tap_1 TAP_14339 (  );
sky130_fd_sc_hd__tap_1 TAP_1434 (  );
sky130_fd_sc_hd__tap_1 TAP_14340 (  );
sky130_fd_sc_hd__tap_1 TAP_14341 (  );
sky130_fd_sc_hd__tap_1 TAP_14342 (  );
sky130_fd_sc_hd__tap_1 TAP_14343 (  );
sky130_fd_sc_hd__tap_1 TAP_14344 (  );
sky130_fd_sc_hd__tap_1 TAP_14345 (  );
sky130_fd_sc_hd__tap_1 TAP_14346 (  );
sky130_fd_sc_hd__tap_1 TAP_14347 (  );
sky130_fd_sc_hd__tap_1 TAP_14348 (  );
sky130_fd_sc_hd__tap_1 TAP_14349 (  );
sky130_fd_sc_hd__tap_1 TAP_1435 (  );
sky130_fd_sc_hd__tap_1 TAP_14350 (  );
sky130_fd_sc_hd__tap_1 TAP_14351 (  );
sky130_fd_sc_hd__tap_1 TAP_14352 (  );
sky130_fd_sc_hd__tap_1 TAP_14353 (  );
sky130_fd_sc_hd__tap_1 TAP_14354 (  );
sky130_fd_sc_hd__tap_1 TAP_14355 (  );
sky130_fd_sc_hd__tap_1 TAP_14356 (  );
sky130_fd_sc_hd__tap_1 TAP_14357 (  );
sky130_fd_sc_hd__tap_1 TAP_14358 (  );
sky130_fd_sc_hd__tap_1 TAP_14359 (  );
sky130_fd_sc_hd__tap_1 TAP_1436 (  );
sky130_fd_sc_hd__tap_1 TAP_14360 (  );
sky130_fd_sc_hd__tap_1 TAP_14361 (  );
sky130_fd_sc_hd__tap_1 TAP_14362 (  );
sky130_fd_sc_hd__tap_1 TAP_14363 (  );
sky130_fd_sc_hd__tap_1 TAP_14364 (  );
sky130_fd_sc_hd__tap_1 TAP_14365 (  );
sky130_fd_sc_hd__tap_1 TAP_14366 (  );
sky130_fd_sc_hd__tap_1 TAP_14367 (  );
sky130_fd_sc_hd__tap_1 TAP_14368 (  );
sky130_fd_sc_hd__tap_1 TAP_14369 (  );
sky130_fd_sc_hd__tap_1 TAP_1437 (  );
sky130_fd_sc_hd__tap_1 TAP_14370 (  );
sky130_fd_sc_hd__tap_1 TAP_14371 (  );
sky130_fd_sc_hd__tap_1 TAP_14372 (  );
sky130_fd_sc_hd__tap_1 TAP_14373 (  );
sky130_fd_sc_hd__tap_1 TAP_14374 (  );
sky130_fd_sc_hd__tap_1 TAP_14375 (  );
sky130_fd_sc_hd__tap_1 TAP_14376 (  );
sky130_fd_sc_hd__tap_1 TAP_14377 (  );
sky130_fd_sc_hd__tap_1 TAP_14378 (  );
sky130_fd_sc_hd__tap_1 TAP_14379 (  );
sky130_fd_sc_hd__tap_1 TAP_1438 (  );
sky130_fd_sc_hd__tap_1 TAP_14380 (  );
sky130_fd_sc_hd__tap_1 TAP_14381 (  );
sky130_fd_sc_hd__tap_1 TAP_14382 (  );
sky130_fd_sc_hd__tap_1 TAP_14383 (  );
sky130_fd_sc_hd__tap_1 TAP_14384 (  );
sky130_fd_sc_hd__tap_1 TAP_14385 (  );
sky130_fd_sc_hd__tap_1 TAP_14386 (  );
sky130_fd_sc_hd__tap_1 TAP_14387 (  );
sky130_fd_sc_hd__tap_1 TAP_14388 (  );
sky130_fd_sc_hd__tap_1 TAP_14389 (  );
sky130_fd_sc_hd__tap_1 TAP_1439 (  );
sky130_fd_sc_hd__tap_1 TAP_14390 (  );
sky130_fd_sc_hd__tap_1 TAP_14391 (  );
sky130_fd_sc_hd__tap_1 TAP_14392 (  );
sky130_fd_sc_hd__tap_1 TAP_14393 (  );
sky130_fd_sc_hd__tap_1 TAP_14394 (  );
sky130_fd_sc_hd__tap_1 TAP_14395 (  );
sky130_fd_sc_hd__tap_1 TAP_14396 (  );
sky130_fd_sc_hd__tap_1 TAP_14397 (  );
sky130_fd_sc_hd__tap_1 TAP_14398 (  );
sky130_fd_sc_hd__tap_1 TAP_14399 (  );
sky130_fd_sc_hd__tap_1 TAP_1440 (  );
sky130_fd_sc_hd__tap_1 TAP_14400 (  );
sky130_fd_sc_hd__tap_1 TAP_14401 (  );
sky130_fd_sc_hd__tap_1 TAP_14402 (  );
sky130_fd_sc_hd__tap_1 TAP_14403 (  );
sky130_fd_sc_hd__tap_1 TAP_14404 (  );
sky130_fd_sc_hd__tap_1 TAP_14405 (  );
sky130_fd_sc_hd__tap_1 TAP_14406 (  );
sky130_fd_sc_hd__tap_1 TAP_14407 (  );
sky130_fd_sc_hd__tap_1 TAP_14408 (  );
sky130_fd_sc_hd__tap_1 TAP_14409 (  );
sky130_fd_sc_hd__tap_1 TAP_1441 (  );
sky130_fd_sc_hd__tap_1 TAP_14410 (  );
sky130_fd_sc_hd__tap_1 TAP_14411 (  );
sky130_fd_sc_hd__tap_1 TAP_14412 (  );
sky130_fd_sc_hd__tap_1 TAP_14413 (  );
sky130_fd_sc_hd__tap_1 TAP_14414 (  );
sky130_fd_sc_hd__tap_1 TAP_14415 (  );
sky130_fd_sc_hd__tap_1 TAP_14416 (  );
sky130_fd_sc_hd__tap_1 TAP_14417 (  );
sky130_fd_sc_hd__tap_1 TAP_14418 (  );
sky130_fd_sc_hd__tap_1 TAP_14419 (  );
sky130_fd_sc_hd__tap_1 TAP_1442 (  );
sky130_fd_sc_hd__tap_1 TAP_14420 (  );
sky130_fd_sc_hd__tap_1 TAP_14421 (  );
sky130_fd_sc_hd__tap_1 TAP_14422 (  );
sky130_fd_sc_hd__tap_1 TAP_14423 (  );
sky130_fd_sc_hd__tap_1 TAP_14424 (  );
sky130_fd_sc_hd__tap_1 TAP_14425 (  );
sky130_fd_sc_hd__tap_1 TAP_14426 (  );
sky130_fd_sc_hd__tap_1 TAP_14427 (  );
sky130_fd_sc_hd__tap_1 TAP_14428 (  );
sky130_fd_sc_hd__tap_1 TAP_14429 (  );
sky130_fd_sc_hd__tap_1 TAP_1443 (  );
sky130_fd_sc_hd__tap_1 TAP_14430 (  );
sky130_fd_sc_hd__tap_1 TAP_14431 (  );
sky130_fd_sc_hd__tap_1 TAP_14432 (  );
sky130_fd_sc_hd__tap_1 TAP_14433 (  );
sky130_fd_sc_hd__tap_1 TAP_14434 (  );
sky130_fd_sc_hd__tap_1 TAP_14435 (  );
sky130_fd_sc_hd__tap_1 TAP_14436 (  );
sky130_fd_sc_hd__tap_1 TAP_14437 (  );
sky130_fd_sc_hd__tap_1 TAP_14438 (  );
sky130_fd_sc_hd__tap_1 TAP_14439 (  );
sky130_fd_sc_hd__tap_1 TAP_1444 (  );
sky130_fd_sc_hd__tap_1 TAP_14440 (  );
sky130_fd_sc_hd__tap_1 TAP_14441 (  );
sky130_fd_sc_hd__tap_1 TAP_14442 (  );
sky130_fd_sc_hd__tap_1 TAP_14443 (  );
sky130_fd_sc_hd__tap_1 TAP_14444 (  );
sky130_fd_sc_hd__tap_1 TAP_14445 (  );
sky130_fd_sc_hd__tap_1 TAP_14446 (  );
sky130_fd_sc_hd__tap_1 TAP_14447 (  );
sky130_fd_sc_hd__tap_1 TAP_14448 (  );
sky130_fd_sc_hd__tap_1 TAP_14449 (  );
sky130_fd_sc_hd__tap_1 TAP_1445 (  );
sky130_fd_sc_hd__tap_1 TAP_14450 (  );
sky130_fd_sc_hd__tap_1 TAP_14451 (  );
sky130_fd_sc_hd__tap_1 TAP_14452 (  );
sky130_fd_sc_hd__tap_1 TAP_14453 (  );
sky130_fd_sc_hd__tap_1 TAP_14454 (  );
sky130_fd_sc_hd__tap_1 TAP_14455 (  );
sky130_fd_sc_hd__tap_1 TAP_14456 (  );
sky130_fd_sc_hd__tap_1 TAP_14457 (  );
sky130_fd_sc_hd__tap_1 TAP_14458 (  );
sky130_fd_sc_hd__tap_1 TAP_14459 (  );
sky130_fd_sc_hd__tap_1 TAP_1446 (  );
sky130_fd_sc_hd__tap_1 TAP_14460 (  );
sky130_fd_sc_hd__tap_1 TAP_14461 (  );
sky130_fd_sc_hd__tap_1 TAP_14462 (  );
sky130_fd_sc_hd__tap_1 TAP_14463 (  );
sky130_fd_sc_hd__tap_1 TAP_14464 (  );
sky130_fd_sc_hd__tap_1 TAP_14465 (  );
sky130_fd_sc_hd__tap_1 TAP_14466 (  );
sky130_fd_sc_hd__tap_1 TAP_14467 (  );
sky130_fd_sc_hd__tap_1 TAP_14468 (  );
sky130_fd_sc_hd__tap_1 TAP_14469 (  );
sky130_fd_sc_hd__tap_1 TAP_1447 (  );
sky130_fd_sc_hd__tap_1 TAP_14470 (  );
sky130_fd_sc_hd__tap_1 TAP_14471 (  );
sky130_fd_sc_hd__tap_1 TAP_14472 (  );
sky130_fd_sc_hd__tap_1 TAP_14473 (  );
sky130_fd_sc_hd__tap_1 TAP_14474 (  );
sky130_fd_sc_hd__tap_1 TAP_14475 (  );
sky130_fd_sc_hd__tap_1 TAP_14476 (  );
sky130_fd_sc_hd__tap_1 TAP_14477 (  );
sky130_fd_sc_hd__tap_1 TAP_14478 (  );
sky130_fd_sc_hd__tap_1 TAP_14479 (  );
sky130_fd_sc_hd__tap_1 TAP_1448 (  );
sky130_fd_sc_hd__tap_1 TAP_14480 (  );
sky130_fd_sc_hd__tap_1 TAP_14481 (  );
sky130_fd_sc_hd__tap_1 TAP_14482 (  );
sky130_fd_sc_hd__tap_1 TAP_14483 (  );
sky130_fd_sc_hd__tap_1 TAP_14484 (  );
sky130_fd_sc_hd__tap_1 TAP_14485 (  );
sky130_fd_sc_hd__tap_1 TAP_14486 (  );
sky130_fd_sc_hd__tap_1 TAP_14487 (  );
sky130_fd_sc_hd__tap_1 TAP_14488 (  );
sky130_fd_sc_hd__tap_1 TAP_14489 (  );
sky130_fd_sc_hd__tap_1 TAP_1449 (  );
sky130_fd_sc_hd__tap_1 TAP_14490 (  );
sky130_fd_sc_hd__tap_1 TAP_14491 (  );
sky130_fd_sc_hd__tap_1 TAP_14492 (  );
sky130_fd_sc_hd__tap_1 TAP_14493 (  );
sky130_fd_sc_hd__tap_1 TAP_14494 (  );
sky130_fd_sc_hd__tap_1 TAP_14495 (  );
sky130_fd_sc_hd__tap_1 TAP_14496 (  );
sky130_fd_sc_hd__tap_1 TAP_14497 (  );
sky130_fd_sc_hd__tap_1 TAP_14498 (  );
sky130_fd_sc_hd__tap_1 TAP_14499 (  );
sky130_fd_sc_hd__tap_1 TAP_1450 (  );
sky130_fd_sc_hd__tap_1 TAP_14500 (  );
sky130_fd_sc_hd__tap_1 TAP_14501 (  );
sky130_fd_sc_hd__tap_1 TAP_14502 (  );
sky130_fd_sc_hd__tap_1 TAP_14503 (  );
sky130_fd_sc_hd__tap_1 TAP_14504 (  );
sky130_fd_sc_hd__tap_1 TAP_14505 (  );
sky130_fd_sc_hd__tap_1 TAP_14506 (  );
sky130_fd_sc_hd__tap_1 TAP_14507 (  );
sky130_fd_sc_hd__tap_1 TAP_14508 (  );
sky130_fd_sc_hd__tap_1 TAP_14509 (  );
sky130_fd_sc_hd__tap_1 TAP_1451 (  );
sky130_fd_sc_hd__tap_1 TAP_14510 (  );
sky130_fd_sc_hd__tap_1 TAP_14511 (  );
sky130_fd_sc_hd__tap_1 TAP_14512 (  );
sky130_fd_sc_hd__tap_1 TAP_14513 (  );
sky130_fd_sc_hd__tap_1 TAP_14514 (  );
sky130_fd_sc_hd__tap_1 TAP_14515 (  );
sky130_fd_sc_hd__tap_1 TAP_14516 (  );
sky130_fd_sc_hd__tap_1 TAP_14517 (  );
sky130_fd_sc_hd__tap_1 TAP_14518 (  );
sky130_fd_sc_hd__tap_1 TAP_14519 (  );
sky130_fd_sc_hd__tap_1 TAP_1452 (  );
sky130_fd_sc_hd__tap_1 TAP_14520 (  );
sky130_fd_sc_hd__tap_1 TAP_14521 (  );
sky130_fd_sc_hd__tap_1 TAP_14522 (  );
sky130_fd_sc_hd__tap_1 TAP_14523 (  );
sky130_fd_sc_hd__tap_1 TAP_14524 (  );
sky130_fd_sc_hd__tap_1 TAP_14525 (  );
sky130_fd_sc_hd__tap_1 TAP_14526 (  );
sky130_fd_sc_hd__tap_1 TAP_14527 (  );
sky130_fd_sc_hd__tap_1 TAP_14528 (  );
sky130_fd_sc_hd__tap_1 TAP_14529 (  );
sky130_fd_sc_hd__tap_1 TAP_1453 (  );
sky130_fd_sc_hd__tap_1 TAP_14530 (  );
sky130_fd_sc_hd__tap_1 TAP_14531 (  );
sky130_fd_sc_hd__tap_1 TAP_14532 (  );
sky130_fd_sc_hd__tap_1 TAP_14533 (  );
sky130_fd_sc_hd__tap_1 TAP_14534 (  );
sky130_fd_sc_hd__tap_1 TAP_14535 (  );
sky130_fd_sc_hd__tap_1 TAP_14536 (  );
sky130_fd_sc_hd__tap_1 TAP_14537 (  );
sky130_fd_sc_hd__tap_1 TAP_14538 (  );
sky130_fd_sc_hd__tap_1 TAP_14539 (  );
sky130_fd_sc_hd__tap_1 TAP_1454 (  );
sky130_fd_sc_hd__tap_1 TAP_14540 (  );
sky130_fd_sc_hd__tap_1 TAP_14541 (  );
sky130_fd_sc_hd__tap_1 TAP_14542 (  );
sky130_fd_sc_hd__tap_1 TAP_14543 (  );
sky130_fd_sc_hd__tap_1 TAP_14544 (  );
sky130_fd_sc_hd__tap_1 TAP_14545 (  );
sky130_fd_sc_hd__tap_1 TAP_14546 (  );
sky130_fd_sc_hd__tap_1 TAP_14547 (  );
sky130_fd_sc_hd__tap_1 TAP_14548 (  );
sky130_fd_sc_hd__tap_1 TAP_14549 (  );
sky130_fd_sc_hd__tap_1 TAP_1455 (  );
sky130_fd_sc_hd__tap_1 TAP_14550 (  );
sky130_fd_sc_hd__tap_1 TAP_14551 (  );
sky130_fd_sc_hd__tap_1 TAP_14552 (  );
sky130_fd_sc_hd__tap_1 TAP_14553 (  );
sky130_fd_sc_hd__tap_1 TAP_14554 (  );
sky130_fd_sc_hd__tap_1 TAP_14555 (  );
sky130_fd_sc_hd__tap_1 TAP_14556 (  );
sky130_fd_sc_hd__tap_1 TAP_14557 (  );
sky130_fd_sc_hd__tap_1 TAP_14558 (  );
sky130_fd_sc_hd__tap_1 TAP_14559 (  );
sky130_fd_sc_hd__tap_1 TAP_1456 (  );
sky130_fd_sc_hd__tap_1 TAP_14560 (  );
sky130_fd_sc_hd__tap_1 TAP_14561 (  );
sky130_fd_sc_hd__tap_1 TAP_14562 (  );
sky130_fd_sc_hd__tap_1 TAP_14563 (  );
sky130_fd_sc_hd__tap_1 TAP_14564 (  );
sky130_fd_sc_hd__tap_1 TAP_14565 (  );
sky130_fd_sc_hd__tap_1 TAP_14566 (  );
sky130_fd_sc_hd__tap_1 TAP_14567 (  );
sky130_fd_sc_hd__tap_1 TAP_14568 (  );
sky130_fd_sc_hd__tap_1 TAP_14569 (  );
sky130_fd_sc_hd__tap_1 TAP_1457 (  );
sky130_fd_sc_hd__tap_1 TAP_14570 (  );
sky130_fd_sc_hd__tap_1 TAP_14571 (  );
sky130_fd_sc_hd__tap_1 TAP_14572 (  );
sky130_fd_sc_hd__tap_1 TAP_14573 (  );
sky130_fd_sc_hd__tap_1 TAP_14574 (  );
sky130_fd_sc_hd__tap_1 TAP_14575 (  );
sky130_fd_sc_hd__tap_1 TAP_14576 (  );
sky130_fd_sc_hd__tap_1 TAP_14577 (  );
sky130_fd_sc_hd__tap_1 TAP_14578 (  );
sky130_fd_sc_hd__tap_1 TAP_14579 (  );
sky130_fd_sc_hd__tap_1 TAP_1458 (  );
sky130_fd_sc_hd__tap_1 TAP_14580 (  );
sky130_fd_sc_hd__tap_1 TAP_14581 (  );
sky130_fd_sc_hd__tap_1 TAP_14582 (  );
sky130_fd_sc_hd__tap_1 TAP_14583 (  );
sky130_fd_sc_hd__tap_1 TAP_14584 (  );
sky130_fd_sc_hd__tap_1 TAP_14585 (  );
sky130_fd_sc_hd__tap_1 TAP_14586 (  );
sky130_fd_sc_hd__tap_1 TAP_14587 (  );
sky130_fd_sc_hd__tap_1 TAP_14588 (  );
sky130_fd_sc_hd__tap_1 TAP_14589 (  );
sky130_fd_sc_hd__tap_1 TAP_1459 (  );
sky130_fd_sc_hd__tap_1 TAP_14590 (  );
sky130_fd_sc_hd__tap_1 TAP_14591 (  );
sky130_fd_sc_hd__tap_1 TAP_14592 (  );
sky130_fd_sc_hd__tap_1 TAP_14593 (  );
sky130_fd_sc_hd__tap_1 TAP_14594 (  );
sky130_fd_sc_hd__tap_1 TAP_14595 (  );
sky130_fd_sc_hd__tap_1 TAP_14596 (  );
sky130_fd_sc_hd__tap_1 TAP_14597 (  );
sky130_fd_sc_hd__tap_1 TAP_14598 (  );
sky130_fd_sc_hd__tap_1 TAP_14599 (  );
sky130_fd_sc_hd__tap_1 TAP_1460 (  );
sky130_fd_sc_hd__tap_1 TAP_14600 (  );
sky130_fd_sc_hd__tap_1 TAP_14601 (  );
sky130_fd_sc_hd__tap_1 TAP_14602 (  );
sky130_fd_sc_hd__tap_1 TAP_14603 (  );
sky130_fd_sc_hd__tap_1 TAP_14604 (  );
sky130_fd_sc_hd__tap_1 TAP_14605 (  );
sky130_fd_sc_hd__tap_1 TAP_14606 (  );
sky130_fd_sc_hd__tap_1 TAP_14607 (  );
sky130_fd_sc_hd__tap_1 TAP_14608 (  );
sky130_fd_sc_hd__tap_1 TAP_14609 (  );
sky130_fd_sc_hd__tap_1 TAP_1461 (  );
sky130_fd_sc_hd__tap_1 TAP_14610 (  );
sky130_fd_sc_hd__tap_1 TAP_14611 (  );
sky130_fd_sc_hd__tap_1 TAP_14612 (  );
sky130_fd_sc_hd__tap_1 TAP_14613 (  );
sky130_fd_sc_hd__tap_1 TAP_14614 (  );
sky130_fd_sc_hd__tap_1 TAP_14615 (  );
sky130_fd_sc_hd__tap_1 TAP_14616 (  );
sky130_fd_sc_hd__tap_1 TAP_14617 (  );
sky130_fd_sc_hd__tap_1 TAP_14618 (  );
sky130_fd_sc_hd__tap_1 TAP_14619 (  );
sky130_fd_sc_hd__tap_1 TAP_1462 (  );
sky130_fd_sc_hd__tap_1 TAP_14620 (  );
sky130_fd_sc_hd__tap_1 TAP_14621 (  );
sky130_fd_sc_hd__tap_1 TAP_14622 (  );
sky130_fd_sc_hd__tap_1 TAP_14623 (  );
sky130_fd_sc_hd__tap_1 TAP_14624 (  );
sky130_fd_sc_hd__tap_1 TAP_14625 (  );
sky130_fd_sc_hd__tap_1 TAP_14626 (  );
sky130_fd_sc_hd__tap_1 TAP_14627 (  );
sky130_fd_sc_hd__tap_1 TAP_14628 (  );
sky130_fd_sc_hd__tap_1 TAP_14629 (  );
sky130_fd_sc_hd__tap_1 TAP_1463 (  );
sky130_fd_sc_hd__tap_1 TAP_14630 (  );
sky130_fd_sc_hd__tap_1 TAP_14631 (  );
sky130_fd_sc_hd__tap_1 TAP_14632 (  );
sky130_fd_sc_hd__tap_1 TAP_14633 (  );
sky130_fd_sc_hd__tap_1 TAP_14634 (  );
sky130_fd_sc_hd__tap_1 TAP_14635 (  );
sky130_fd_sc_hd__tap_1 TAP_14636 (  );
sky130_fd_sc_hd__tap_1 TAP_14637 (  );
sky130_fd_sc_hd__tap_1 TAP_14638 (  );
sky130_fd_sc_hd__tap_1 TAP_14639 (  );
sky130_fd_sc_hd__tap_1 TAP_1464 (  );
sky130_fd_sc_hd__tap_1 TAP_14640 (  );
sky130_fd_sc_hd__tap_1 TAP_14641 (  );
sky130_fd_sc_hd__tap_1 TAP_14642 (  );
sky130_fd_sc_hd__tap_1 TAP_14643 (  );
sky130_fd_sc_hd__tap_1 TAP_14644 (  );
sky130_fd_sc_hd__tap_1 TAP_14645 (  );
sky130_fd_sc_hd__tap_1 TAP_14646 (  );
sky130_fd_sc_hd__tap_1 TAP_14647 (  );
sky130_fd_sc_hd__tap_1 TAP_14648 (  );
sky130_fd_sc_hd__tap_1 TAP_14649 (  );
sky130_fd_sc_hd__tap_1 TAP_1465 (  );
sky130_fd_sc_hd__tap_1 TAP_14650 (  );
sky130_fd_sc_hd__tap_1 TAP_14651 (  );
sky130_fd_sc_hd__tap_1 TAP_14652 (  );
sky130_fd_sc_hd__tap_1 TAP_14653 (  );
sky130_fd_sc_hd__tap_1 TAP_14654 (  );
sky130_fd_sc_hd__tap_1 TAP_14655 (  );
sky130_fd_sc_hd__tap_1 TAP_14656 (  );
sky130_fd_sc_hd__tap_1 TAP_14657 (  );
sky130_fd_sc_hd__tap_1 TAP_14658 (  );
sky130_fd_sc_hd__tap_1 TAP_14659 (  );
sky130_fd_sc_hd__tap_1 TAP_1466 (  );
sky130_fd_sc_hd__tap_1 TAP_14660 (  );
sky130_fd_sc_hd__tap_1 TAP_14661 (  );
sky130_fd_sc_hd__tap_1 TAP_14662 (  );
sky130_fd_sc_hd__tap_1 TAP_14663 (  );
sky130_fd_sc_hd__tap_1 TAP_14664 (  );
sky130_fd_sc_hd__tap_1 TAP_14665 (  );
sky130_fd_sc_hd__tap_1 TAP_14666 (  );
sky130_fd_sc_hd__tap_1 TAP_14667 (  );
sky130_fd_sc_hd__tap_1 TAP_14668 (  );
sky130_fd_sc_hd__tap_1 TAP_14669 (  );
sky130_fd_sc_hd__tap_1 TAP_1467 (  );
sky130_fd_sc_hd__tap_1 TAP_14670 (  );
sky130_fd_sc_hd__tap_1 TAP_14671 (  );
sky130_fd_sc_hd__tap_1 TAP_14672 (  );
sky130_fd_sc_hd__tap_1 TAP_14673 (  );
sky130_fd_sc_hd__tap_1 TAP_14674 (  );
sky130_fd_sc_hd__tap_1 TAP_14675 (  );
sky130_fd_sc_hd__tap_1 TAP_14676 (  );
sky130_fd_sc_hd__tap_1 TAP_14677 (  );
sky130_fd_sc_hd__tap_1 TAP_14678 (  );
sky130_fd_sc_hd__tap_1 TAP_14679 (  );
sky130_fd_sc_hd__tap_1 TAP_1468 (  );
sky130_fd_sc_hd__tap_1 TAP_14680 (  );
sky130_fd_sc_hd__tap_1 TAP_14681 (  );
sky130_fd_sc_hd__tap_1 TAP_14682 (  );
sky130_fd_sc_hd__tap_1 TAP_14683 (  );
sky130_fd_sc_hd__tap_1 TAP_14684 (  );
sky130_fd_sc_hd__tap_1 TAP_14685 (  );
sky130_fd_sc_hd__tap_1 TAP_14686 (  );
sky130_fd_sc_hd__tap_1 TAP_14687 (  );
sky130_fd_sc_hd__tap_1 TAP_14688 (  );
sky130_fd_sc_hd__tap_1 TAP_14689 (  );
sky130_fd_sc_hd__tap_1 TAP_1469 (  );
sky130_fd_sc_hd__tap_1 TAP_14690 (  );
sky130_fd_sc_hd__tap_1 TAP_14691 (  );
sky130_fd_sc_hd__tap_1 TAP_14692 (  );
sky130_fd_sc_hd__tap_1 TAP_14693 (  );
sky130_fd_sc_hd__tap_1 TAP_14694 (  );
sky130_fd_sc_hd__tap_1 TAP_14695 (  );
sky130_fd_sc_hd__tap_1 TAP_14696 (  );
sky130_fd_sc_hd__tap_1 TAP_14697 (  );
sky130_fd_sc_hd__tap_1 TAP_14698 (  );
sky130_fd_sc_hd__tap_1 TAP_14699 (  );
sky130_fd_sc_hd__tap_1 TAP_1470 (  );
sky130_fd_sc_hd__tap_1 TAP_14700 (  );
sky130_fd_sc_hd__tap_1 TAP_14701 (  );
sky130_fd_sc_hd__tap_1 TAP_14702 (  );
sky130_fd_sc_hd__tap_1 TAP_14703 (  );
sky130_fd_sc_hd__tap_1 TAP_14704 (  );
sky130_fd_sc_hd__tap_1 TAP_14705 (  );
sky130_fd_sc_hd__tap_1 TAP_14706 (  );
sky130_fd_sc_hd__tap_1 TAP_14707 (  );
sky130_fd_sc_hd__tap_1 TAP_14708 (  );
sky130_fd_sc_hd__tap_1 TAP_14709 (  );
sky130_fd_sc_hd__tap_1 TAP_1471 (  );
sky130_fd_sc_hd__tap_1 TAP_14710 (  );
sky130_fd_sc_hd__tap_1 TAP_14711 (  );
sky130_fd_sc_hd__tap_1 TAP_14712 (  );
sky130_fd_sc_hd__tap_1 TAP_14713 (  );
sky130_fd_sc_hd__tap_1 TAP_14714 (  );
sky130_fd_sc_hd__tap_1 TAP_14715 (  );
sky130_fd_sc_hd__tap_1 TAP_14716 (  );
sky130_fd_sc_hd__tap_1 TAP_14717 (  );
sky130_fd_sc_hd__tap_1 TAP_14718 (  );
sky130_fd_sc_hd__tap_1 TAP_14719 (  );
sky130_fd_sc_hd__tap_1 TAP_1472 (  );
sky130_fd_sc_hd__tap_1 TAP_14720 (  );
sky130_fd_sc_hd__tap_1 TAP_14721 (  );
sky130_fd_sc_hd__tap_1 TAP_14722 (  );
sky130_fd_sc_hd__tap_1 TAP_14723 (  );
sky130_fd_sc_hd__tap_1 TAP_14724 (  );
sky130_fd_sc_hd__tap_1 TAP_14725 (  );
sky130_fd_sc_hd__tap_1 TAP_14726 (  );
sky130_fd_sc_hd__tap_1 TAP_14727 (  );
sky130_fd_sc_hd__tap_1 TAP_14728 (  );
sky130_fd_sc_hd__tap_1 TAP_14729 (  );
sky130_fd_sc_hd__tap_1 TAP_1473 (  );
sky130_fd_sc_hd__tap_1 TAP_14730 (  );
sky130_fd_sc_hd__tap_1 TAP_14731 (  );
sky130_fd_sc_hd__tap_1 TAP_14732 (  );
sky130_fd_sc_hd__tap_1 TAP_14733 (  );
sky130_fd_sc_hd__tap_1 TAP_14734 (  );
sky130_fd_sc_hd__tap_1 TAP_14735 (  );
sky130_fd_sc_hd__tap_1 TAP_14736 (  );
sky130_fd_sc_hd__tap_1 TAP_14737 (  );
sky130_fd_sc_hd__tap_1 TAP_14738 (  );
sky130_fd_sc_hd__tap_1 TAP_14739 (  );
sky130_fd_sc_hd__tap_1 TAP_1474 (  );
sky130_fd_sc_hd__tap_1 TAP_14740 (  );
sky130_fd_sc_hd__tap_1 TAP_14741 (  );
sky130_fd_sc_hd__tap_1 TAP_14742 (  );
sky130_fd_sc_hd__tap_1 TAP_14743 (  );
sky130_fd_sc_hd__tap_1 TAP_14744 (  );
sky130_fd_sc_hd__tap_1 TAP_14745 (  );
sky130_fd_sc_hd__tap_1 TAP_14746 (  );
sky130_fd_sc_hd__tap_1 TAP_14747 (  );
sky130_fd_sc_hd__tap_1 TAP_14748 (  );
sky130_fd_sc_hd__tap_1 TAP_14749 (  );
sky130_fd_sc_hd__tap_1 TAP_1475 (  );
sky130_fd_sc_hd__tap_1 TAP_14750 (  );
sky130_fd_sc_hd__tap_1 TAP_14751 (  );
sky130_fd_sc_hd__tap_1 TAP_14752 (  );
sky130_fd_sc_hd__tap_1 TAP_14753 (  );
sky130_fd_sc_hd__tap_1 TAP_14754 (  );
sky130_fd_sc_hd__tap_1 TAP_14755 (  );
sky130_fd_sc_hd__tap_1 TAP_14756 (  );
sky130_fd_sc_hd__tap_1 TAP_14757 (  );
sky130_fd_sc_hd__tap_1 TAP_14758 (  );
sky130_fd_sc_hd__tap_1 TAP_14759 (  );
sky130_fd_sc_hd__tap_1 TAP_1476 (  );
sky130_fd_sc_hd__tap_1 TAP_14760 (  );
sky130_fd_sc_hd__tap_1 TAP_14761 (  );
sky130_fd_sc_hd__tap_1 TAP_14762 (  );
sky130_fd_sc_hd__tap_1 TAP_14763 (  );
sky130_fd_sc_hd__tap_1 TAP_14764 (  );
sky130_fd_sc_hd__tap_1 TAP_14765 (  );
sky130_fd_sc_hd__tap_1 TAP_14766 (  );
sky130_fd_sc_hd__tap_1 TAP_14767 (  );
sky130_fd_sc_hd__tap_1 TAP_14768 (  );
sky130_fd_sc_hd__tap_1 TAP_14769 (  );
sky130_fd_sc_hd__tap_1 TAP_1477 (  );
sky130_fd_sc_hd__tap_1 TAP_14770 (  );
sky130_fd_sc_hd__tap_1 TAP_14771 (  );
sky130_fd_sc_hd__tap_1 TAP_14772 (  );
sky130_fd_sc_hd__tap_1 TAP_14773 (  );
sky130_fd_sc_hd__tap_1 TAP_14774 (  );
sky130_fd_sc_hd__tap_1 TAP_14775 (  );
sky130_fd_sc_hd__tap_1 TAP_14776 (  );
sky130_fd_sc_hd__tap_1 TAP_14777 (  );
sky130_fd_sc_hd__tap_1 TAP_14778 (  );
sky130_fd_sc_hd__tap_1 TAP_14779 (  );
sky130_fd_sc_hd__tap_1 TAP_1478 (  );
sky130_fd_sc_hd__tap_1 TAP_14780 (  );
sky130_fd_sc_hd__tap_1 TAP_14781 (  );
sky130_fd_sc_hd__tap_1 TAP_14782 (  );
sky130_fd_sc_hd__tap_1 TAP_14783 (  );
sky130_fd_sc_hd__tap_1 TAP_14784 (  );
sky130_fd_sc_hd__tap_1 TAP_14785 (  );
sky130_fd_sc_hd__tap_1 TAP_14786 (  );
sky130_fd_sc_hd__tap_1 TAP_14787 (  );
sky130_fd_sc_hd__tap_1 TAP_14788 (  );
sky130_fd_sc_hd__tap_1 TAP_14789 (  );
sky130_fd_sc_hd__tap_1 TAP_1479 (  );
sky130_fd_sc_hd__tap_1 TAP_14790 (  );
sky130_fd_sc_hd__tap_1 TAP_14791 (  );
sky130_fd_sc_hd__tap_1 TAP_14792 (  );
sky130_fd_sc_hd__tap_1 TAP_14793 (  );
sky130_fd_sc_hd__tap_1 TAP_14794 (  );
sky130_fd_sc_hd__tap_1 TAP_14795 (  );
sky130_fd_sc_hd__tap_1 TAP_14796 (  );
sky130_fd_sc_hd__tap_1 TAP_14797 (  );
sky130_fd_sc_hd__tap_1 TAP_14798 (  );
sky130_fd_sc_hd__tap_1 TAP_14799 (  );
sky130_fd_sc_hd__tap_1 TAP_1480 (  );
sky130_fd_sc_hd__tap_1 TAP_14800 (  );
sky130_fd_sc_hd__tap_1 TAP_14801 (  );
sky130_fd_sc_hd__tap_1 TAP_14802 (  );
sky130_fd_sc_hd__tap_1 TAP_14803 (  );
sky130_fd_sc_hd__tap_1 TAP_14804 (  );
sky130_fd_sc_hd__tap_1 TAP_14805 (  );
sky130_fd_sc_hd__tap_1 TAP_14806 (  );
sky130_fd_sc_hd__tap_1 TAP_14807 (  );
sky130_fd_sc_hd__tap_1 TAP_14808 (  );
sky130_fd_sc_hd__tap_1 TAP_14809 (  );
sky130_fd_sc_hd__tap_1 TAP_1481 (  );
sky130_fd_sc_hd__tap_1 TAP_14810 (  );
sky130_fd_sc_hd__tap_1 TAP_14811 (  );
sky130_fd_sc_hd__tap_1 TAP_14812 (  );
sky130_fd_sc_hd__tap_1 TAP_14813 (  );
sky130_fd_sc_hd__tap_1 TAP_14814 (  );
sky130_fd_sc_hd__tap_1 TAP_14815 (  );
sky130_fd_sc_hd__tap_1 TAP_14816 (  );
sky130_fd_sc_hd__tap_1 TAP_14817 (  );
sky130_fd_sc_hd__tap_1 TAP_14818 (  );
sky130_fd_sc_hd__tap_1 TAP_14819 (  );
sky130_fd_sc_hd__tap_1 TAP_1482 (  );
sky130_fd_sc_hd__tap_1 TAP_14820 (  );
sky130_fd_sc_hd__tap_1 TAP_14821 (  );
sky130_fd_sc_hd__tap_1 TAP_14822 (  );
sky130_fd_sc_hd__tap_1 TAP_14823 (  );
sky130_fd_sc_hd__tap_1 TAP_14824 (  );
sky130_fd_sc_hd__tap_1 TAP_14825 (  );
sky130_fd_sc_hd__tap_1 TAP_14826 (  );
sky130_fd_sc_hd__tap_1 TAP_14827 (  );
sky130_fd_sc_hd__tap_1 TAP_14828 (  );
sky130_fd_sc_hd__tap_1 TAP_14829 (  );
sky130_fd_sc_hd__tap_1 TAP_1483 (  );
sky130_fd_sc_hd__tap_1 TAP_14830 (  );
sky130_fd_sc_hd__tap_1 TAP_14831 (  );
sky130_fd_sc_hd__tap_1 TAP_14832 (  );
sky130_fd_sc_hd__tap_1 TAP_14833 (  );
sky130_fd_sc_hd__tap_1 TAP_14834 (  );
sky130_fd_sc_hd__tap_1 TAP_14835 (  );
sky130_fd_sc_hd__tap_1 TAP_14836 (  );
sky130_fd_sc_hd__tap_1 TAP_14837 (  );
sky130_fd_sc_hd__tap_1 TAP_14838 (  );
sky130_fd_sc_hd__tap_1 TAP_14839 (  );
sky130_fd_sc_hd__tap_1 TAP_1484 (  );
sky130_fd_sc_hd__tap_1 TAP_14840 (  );
sky130_fd_sc_hd__tap_1 TAP_14841 (  );
sky130_fd_sc_hd__tap_1 TAP_14842 (  );
sky130_fd_sc_hd__tap_1 TAP_14843 (  );
sky130_fd_sc_hd__tap_1 TAP_14844 (  );
sky130_fd_sc_hd__tap_1 TAP_14845 (  );
sky130_fd_sc_hd__tap_1 TAP_14846 (  );
sky130_fd_sc_hd__tap_1 TAP_14847 (  );
sky130_fd_sc_hd__tap_1 TAP_14848 (  );
sky130_fd_sc_hd__tap_1 TAP_14849 (  );
sky130_fd_sc_hd__tap_1 TAP_1485 (  );
sky130_fd_sc_hd__tap_1 TAP_14850 (  );
sky130_fd_sc_hd__tap_1 TAP_14851 (  );
sky130_fd_sc_hd__tap_1 TAP_14852 (  );
sky130_fd_sc_hd__tap_1 TAP_14853 (  );
sky130_fd_sc_hd__tap_1 TAP_14854 (  );
sky130_fd_sc_hd__tap_1 TAP_14855 (  );
sky130_fd_sc_hd__tap_1 TAP_14856 (  );
sky130_fd_sc_hd__tap_1 TAP_14857 (  );
sky130_fd_sc_hd__tap_1 TAP_14858 (  );
sky130_fd_sc_hd__tap_1 TAP_14859 (  );
sky130_fd_sc_hd__tap_1 TAP_1486 (  );
sky130_fd_sc_hd__tap_1 TAP_14860 (  );
sky130_fd_sc_hd__tap_1 TAP_14861 (  );
sky130_fd_sc_hd__tap_1 TAP_14862 (  );
sky130_fd_sc_hd__tap_1 TAP_14863 (  );
sky130_fd_sc_hd__tap_1 TAP_14864 (  );
sky130_fd_sc_hd__tap_1 TAP_14865 (  );
sky130_fd_sc_hd__tap_1 TAP_14866 (  );
sky130_fd_sc_hd__tap_1 TAP_14867 (  );
sky130_fd_sc_hd__tap_1 TAP_14868 (  );
sky130_fd_sc_hd__tap_1 TAP_14869 (  );
sky130_fd_sc_hd__tap_1 TAP_1487 (  );
sky130_fd_sc_hd__tap_1 TAP_14870 (  );
sky130_fd_sc_hd__tap_1 TAP_14871 (  );
sky130_fd_sc_hd__tap_1 TAP_14872 (  );
sky130_fd_sc_hd__tap_1 TAP_14873 (  );
sky130_fd_sc_hd__tap_1 TAP_14874 (  );
sky130_fd_sc_hd__tap_1 TAP_14875 (  );
sky130_fd_sc_hd__tap_1 TAP_14876 (  );
sky130_fd_sc_hd__tap_1 TAP_14877 (  );
sky130_fd_sc_hd__tap_1 TAP_14878 (  );
sky130_fd_sc_hd__tap_1 TAP_14879 (  );
sky130_fd_sc_hd__tap_1 TAP_1488 (  );
sky130_fd_sc_hd__tap_1 TAP_14880 (  );
sky130_fd_sc_hd__tap_1 TAP_14881 (  );
sky130_fd_sc_hd__tap_1 TAP_14882 (  );
sky130_fd_sc_hd__tap_1 TAP_14883 (  );
sky130_fd_sc_hd__tap_1 TAP_14884 (  );
sky130_fd_sc_hd__tap_1 TAP_14885 (  );
sky130_fd_sc_hd__tap_1 TAP_14886 (  );
sky130_fd_sc_hd__tap_1 TAP_14887 (  );
sky130_fd_sc_hd__tap_1 TAP_14888 (  );
sky130_fd_sc_hd__tap_1 TAP_14889 (  );
sky130_fd_sc_hd__tap_1 TAP_1489 (  );
sky130_fd_sc_hd__tap_1 TAP_14890 (  );
sky130_fd_sc_hd__tap_1 TAP_14891 (  );
sky130_fd_sc_hd__tap_1 TAP_14892 (  );
sky130_fd_sc_hd__tap_1 TAP_14893 (  );
sky130_fd_sc_hd__tap_1 TAP_14894 (  );
sky130_fd_sc_hd__tap_1 TAP_14895 (  );
sky130_fd_sc_hd__tap_1 TAP_14896 (  );
sky130_fd_sc_hd__tap_1 TAP_14897 (  );
sky130_fd_sc_hd__tap_1 TAP_14898 (  );
sky130_fd_sc_hd__tap_1 TAP_14899 (  );
sky130_fd_sc_hd__tap_1 TAP_1490 (  );
sky130_fd_sc_hd__tap_1 TAP_14900 (  );
sky130_fd_sc_hd__tap_1 TAP_14901 (  );
sky130_fd_sc_hd__tap_1 TAP_14902 (  );
sky130_fd_sc_hd__tap_1 TAP_14903 (  );
sky130_fd_sc_hd__tap_1 TAP_14904 (  );
sky130_fd_sc_hd__tap_1 TAP_14905 (  );
sky130_fd_sc_hd__tap_1 TAP_14906 (  );
sky130_fd_sc_hd__tap_1 TAP_14907 (  );
sky130_fd_sc_hd__tap_1 TAP_14908 (  );
sky130_fd_sc_hd__tap_1 TAP_14909 (  );
sky130_fd_sc_hd__tap_1 TAP_1491 (  );
sky130_fd_sc_hd__tap_1 TAP_14910 (  );
sky130_fd_sc_hd__tap_1 TAP_14911 (  );
sky130_fd_sc_hd__tap_1 TAP_14912 (  );
sky130_fd_sc_hd__tap_1 TAP_14913 (  );
sky130_fd_sc_hd__tap_1 TAP_14914 (  );
sky130_fd_sc_hd__tap_1 TAP_14915 (  );
sky130_fd_sc_hd__tap_1 TAP_14916 (  );
sky130_fd_sc_hd__tap_1 TAP_14917 (  );
sky130_fd_sc_hd__tap_1 TAP_14918 (  );
sky130_fd_sc_hd__tap_1 TAP_14919 (  );
sky130_fd_sc_hd__tap_1 TAP_1492 (  );
sky130_fd_sc_hd__tap_1 TAP_14920 (  );
sky130_fd_sc_hd__tap_1 TAP_14921 (  );
sky130_fd_sc_hd__tap_1 TAP_14922 (  );
sky130_fd_sc_hd__tap_1 TAP_14923 (  );
sky130_fd_sc_hd__tap_1 TAP_14924 (  );
sky130_fd_sc_hd__tap_1 TAP_14925 (  );
sky130_fd_sc_hd__tap_1 TAP_14926 (  );
sky130_fd_sc_hd__tap_1 TAP_14927 (  );
sky130_fd_sc_hd__tap_1 TAP_14928 (  );
sky130_fd_sc_hd__tap_1 TAP_14929 (  );
sky130_fd_sc_hd__tap_1 TAP_1493 (  );
sky130_fd_sc_hd__tap_1 TAP_14930 (  );
sky130_fd_sc_hd__tap_1 TAP_14931 (  );
sky130_fd_sc_hd__tap_1 TAP_14932 (  );
sky130_fd_sc_hd__tap_1 TAP_14933 (  );
sky130_fd_sc_hd__tap_1 TAP_14934 (  );
sky130_fd_sc_hd__tap_1 TAP_14935 (  );
sky130_fd_sc_hd__tap_1 TAP_14936 (  );
sky130_fd_sc_hd__tap_1 TAP_14937 (  );
sky130_fd_sc_hd__tap_1 TAP_14938 (  );
sky130_fd_sc_hd__tap_1 TAP_14939 (  );
sky130_fd_sc_hd__tap_1 TAP_1494 (  );
sky130_fd_sc_hd__tap_1 TAP_14940 (  );
sky130_fd_sc_hd__tap_1 TAP_14941 (  );
sky130_fd_sc_hd__tap_1 TAP_14942 (  );
sky130_fd_sc_hd__tap_1 TAP_14943 (  );
sky130_fd_sc_hd__tap_1 TAP_14944 (  );
sky130_fd_sc_hd__tap_1 TAP_14945 (  );
sky130_fd_sc_hd__tap_1 TAP_14946 (  );
sky130_fd_sc_hd__tap_1 TAP_14947 (  );
sky130_fd_sc_hd__tap_1 TAP_14948 (  );
sky130_fd_sc_hd__tap_1 TAP_14949 (  );
sky130_fd_sc_hd__tap_1 TAP_1495 (  );
sky130_fd_sc_hd__tap_1 TAP_14950 (  );
sky130_fd_sc_hd__tap_1 TAP_14951 (  );
sky130_fd_sc_hd__tap_1 TAP_14952 (  );
sky130_fd_sc_hd__tap_1 TAP_14953 (  );
sky130_fd_sc_hd__tap_1 TAP_14954 (  );
sky130_fd_sc_hd__tap_1 TAP_14955 (  );
sky130_fd_sc_hd__tap_1 TAP_14956 (  );
sky130_fd_sc_hd__tap_1 TAP_14957 (  );
sky130_fd_sc_hd__tap_1 TAP_14958 (  );
sky130_fd_sc_hd__tap_1 TAP_14959 (  );
sky130_fd_sc_hd__tap_1 TAP_1496 (  );
sky130_fd_sc_hd__tap_1 TAP_14960 (  );
sky130_fd_sc_hd__tap_1 TAP_14961 (  );
sky130_fd_sc_hd__tap_1 TAP_14962 (  );
sky130_fd_sc_hd__tap_1 TAP_14963 (  );
sky130_fd_sc_hd__tap_1 TAP_14964 (  );
sky130_fd_sc_hd__tap_1 TAP_14965 (  );
sky130_fd_sc_hd__tap_1 TAP_14966 (  );
sky130_fd_sc_hd__tap_1 TAP_14967 (  );
sky130_fd_sc_hd__tap_1 TAP_14968 (  );
sky130_fd_sc_hd__tap_1 TAP_14969 (  );
sky130_fd_sc_hd__tap_1 TAP_1497 (  );
sky130_fd_sc_hd__tap_1 TAP_14970 (  );
sky130_fd_sc_hd__tap_1 TAP_14971 (  );
sky130_fd_sc_hd__tap_1 TAP_14972 (  );
sky130_fd_sc_hd__tap_1 TAP_14973 (  );
sky130_fd_sc_hd__tap_1 TAP_14974 (  );
sky130_fd_sc_hd__tap_1 TAP_14975 (  );
sky130_fd_sc_hd__tap_1 TAP_14976 (  );
sky130_fd_sc_hd__tap_1 TAP_14977 (  );
sky130_fd_sc_hd__tap_1 TAP_14978 (  );
sky130_fd_sc_hd__tap_1 TAP_14979 (  );
sky130_fd_sc_hd__tap_1 TAP_1498 (  );
sky130_fd_sc_hd__tap_1 TAP_14980 (  );
sky130_fd_sc_hd__tap_1 TAP_14981 (  );
sky130_fd_sc_hd__tap_1 TAP_14982 (  );
sky130_fd_sc_hd__tap_1 TAP_14983 (  );
sky130_fd_sc_hd__tap_1 TAP_14984 (  );
sky130_fd_sc_hd__tap_1 TAP_14985 (  );
sky130_fd_sc_hd__tap_1 TAP_14986 (  );
sky130_fd_sc_hd__tap_1 TAP_14987 (  );
sky130_fd_sc_hd__tap_1 TAP_14988 (  );
sky130_fd_sc_hd__tap_1 TAP_14989 (  );
sky130_fd_sc_hd__tap_1 TAP_1499 (  );
sky130_fd_sc_hd__tap_1 TAP_14990 (  );
sky130_fd_sc_hd__tap_1 TAP_14991 (  );
sky130_fd_sc_hd__tap_1 TAP_14992 (  );
sky130_fd_sc_hd__tap_1 TAP_14993 (  );
sky130_fd_sc_hd__tap_1 TAP_14994 (  );
sky130_fd_sc_hd__tap_1 TAP_14995 (  );
sky130_fd_sc_hd__tap_1 TAP_14996 (  );
sky130_fd_sc_hd__tap_1 TAP_14997 (  );
sky130_fd_sc_hd__tap_1 TAP_14998 (  );
sky130_fd_sc_hd__tap_1 TAP_14999 (  );
sky130_fd_sc_hd__tap_1 TAP_1500 (  );
sky130_fd_sc_hd__tap_1 TAP_15000 (  );
sky130_fd_sc_hd__tap_1 TAP_15001 (  );
sky130_fd_sc_hd__tap_1 TAP_15002 (  );
sky130_fd_sc_hd__tap_1 TAP_15003 (  );
sky130_fd_sc_hd__tap_1 TAP_15004 (  );
sky130_fd_sc_hd__tap_1 TAP_15005 (  );
sky130_fd_sc_hd__tap_1 TAP_15006 (  );
sky130_fd_sc_hd__tap_1 TAP_15007 (  );
sky130_fd_sc_hd__tap_1 TAP_15008 (  );
sky130_fd_sc_hd__tap_1 TAP_15009 (  );
sky130_fd_sc_hd__tap_1 TAP_1501 (  );
sky130_fd_sc_hd__tap_1 TAP_15010 (  );
sky130_fd_sc_hd__tap_1 TAP_15011 (  );
sky130_fd_sc_hd__tap_1 TAP_15012 (  );
sky130_fd_sc_hd__tap_1 TAP_15013 (  );
sky130_fd_sc_hd__tap_1 TAP_15014 (  );
sky130_fd_sc_hd__tap_1 TAP_15015 (  );
sky130_fd_sc_hd__tap_1 TAP_15016 (  );
sky130_fd_sc_hd__tap_1 TAP_15017 (  );
sky130_fd_sc_hd__tap_1 TAP_15018 (  );
sky130_fd_sc_hd__tap_1 TAP_15019 (  );
sky130_fd_sc_hd__tap_1 TAP_1502 (  );
sky130_fd_sc_hd__tap_1 TAP_15020 (  );
sky130_fd_sc_hd__tap_1 TAP_15021 (  );
sky130_fd_sc_hd__tap_1 TAP_15022 (  );
sky130_fd_sc_hd__tap_1 TAP_15023 (  );
sky130_fd_sc_hd__tap_1 TAP_15024 (  );
sky130_fd_sc_hd__tap_1 TAP_15025 (  );
sky130_fd_sc_hd__tap_1 TAP_15026 (  );
sky130_fd_sc_hd__tap_1 TAP_15027 (  );
sky130_fd_sc_hd__tap_1 TAP_15028 (  );
sky130_fd_sc_hd__tap_1 TAP_15029 (  );
sky130_fd_sc_hd__tap_1 TAP_1503 (  );
sky130_fd_sc_hd__tap_1 TAP_15030 (  );
sky130_fd_sc_hd__tap_1 TAP_15031 (  );
sky130_fd_sc_hd__tap_1 TAP_15032 (  );
sky130_fd_sc_hd__tap_1 TAP_15033 (  );
sky130_fd_sc_hd__tap_1 TAP_15034 (  );
sky130_fd_sc_hd__tap_1 TAP_15035 (  );
sky130_fd_sc_hd__tap_1 TAP_15036 (  );
sky130_fd_sc_hd__tap_1 TAP_15037 (  );
sky130_fd_sc_hd__tap_1 TAP_15038 (  );
sky130_fd_sc_hd__tap_1 TAP_15039 (  );
sky130_fd_sc_hd__tap_1 TAP_1504 (  );
sky130_fd_sc_hd__tap_1 TAP_15040 (  );
sky130_fd_sc_hd__tap_1 TAP_15041 (  );
sky130_fd_sc_hd__tap_1 TAP_15042 (  );
sky130_fd_sc_hd__tap_1 TAP_15043 (  );
sky130_fd_sc_hd__tap_1 TAP_15044 (  );
sky130_fd_sc_hd__tap_1 TAP_15045 (  );
sky130_fd_sc_hd__tap_1 TAP_15046 (  );
sky130_fd_sc_hd__tap_1 TAP_15047 (  );
sky130_fd_sc_hd__tap_1 TAP_15048 (  );
sky130_fd_sc_hd__tap_1 TAP_15049 (  );
sky130_fd_sc_hd__tap_1 TAP_1505 (  );
sky130_fd_sc_hd__tap_1 TAP_15050 (  );
sky130_fd_sc_hd__tap_1 TAP_15051 (  );
sky130_fd_sc_hd__tap_1 TAP_15052 (  );
sky130_fd_sc_hd__tap_1 TAP_15053 (  );
sky130_fd_sc_hd__tap_1 TAP_15054 (  );
sky130_fd_sc_hd__tap_1 TAP_15055 (  );
sky130_fd_sc_hd__tap_1 TAP_15056 (  );
sky130_fd_sc_hd__tap_1 TAP_15057 (  );
sky130_fd_sc_hd__tap_1 TAP_15058 (  );
sky130_fd_sc_hd__tap_1 TAP_15059 (  );
sky130_fd_sc_hd__tap_1 TAP_1506 (  );
sky130_fd_sc_hd__tap_1 TAP_15060 (  );
sky130_fd_sc_hd__tap_1 TAP_15061 (  );
sky130_fd_sc_hd__tap_1 TAP_15062 (  );
sky130_fd_sc_hd__tap_1 TAP_15063 (  );
sky130_fd_sc_hd__tap_1 TAP_15064 (  );
sky130_fd_sc_hd__tap_1 TAP_15065 (  );
sky130_fd_sc_hd__tap_1 TAP_15066 (  );
sky130_fd_sc_hd__tap_1 TAP_15067 (  );
sky130_fd_sc_hd__tap_1 TAP_15068 (  );
sky130_fd_sc_hd__tap_1 TAP_15069 (  );
sky130_fd_sc_hd__tap_1 TAP_1507 (  );
sky130_fd_sc_hd__tap_1 TAP_15070 (  );
sky130_fd_sc_hd__tap_1 TAP_15071 (  );
sky130_fd_sc_hd__tap_1 TAP_15072 (  );
sky130_fd_sc_hd__tap_1 TAP_15073 (  );
sky130_fd_sc_hd__tap_1 TAP_15074 (  );
sky130_fd_sc_hd__tap_1 TAP_15075 (  );
sky130_fd_sc_hd__tap_1 TAP_15076 (  );
sky130_fd_sc_hd__tap_1 TAP_15077 (  );
sky130_fd_sc_hd__tap_1 TAP_15078 (  );
sky130_fd_sc_hd__tap_1 TAP_15079 (  );
sky130_fd_sc_hd__tap_1 TAP_1508 (  );
sky130_fd_sc_hd__tap_1 TAP_15080 (  );
sky130_fd_sc_hd__tap_1 TAP_15081 (  );
sky130_fd_sc_hd__tap_1 TAP_15082 (  );
sky130_fd_sc_hd__tap_1 TAP_15083 (  );
sky130_fd_sc_hd__tap_1 TAP_15084 (  );
sky130_fd_sc_hd__tap_1 TAP_15085 (  );
sky130_fd_sc_hd__tap_1 TAP_15086 (  );
sky130_fd_sc_hd__tap_1 TAP_15087 (  );
sky130_fd_sc_hd__tap_1 TAP_15088 (  );
sky130_fd_sc_hd__tap_1 TAP_15089 (  );
sky130_fd_sc_hd__tap_1 TAP_1509 (  );
sky130_fd_sc_hd__tap_1 TAP_15090 (  );
sky130_fd_sc_hd__tap_1 TAP_15091 (  );
sky130_fd_sc_hd__tap_1 TAP_15092 (  );
sky130_fd_sc_hd__tap_1 TAP_15093 (  );
sky130_fd_sc_hd__tap_1 TAP_15094 (  );
sky130_fd_sc_hd__tap_1 TAP_15095 (  );
sky130_fd_sc_hd__tap_1 TAP_15096 (  );
sky130_fd_sc_hd__tap_1 TAP_15097 (  );
sky130_fd_sc_hd__tap_1 TAP_15098 (  );
sky130_fd_sc_hd__tap_1 TAP_15099 (  );
sky130_fd_sc_hd__tap_1 TAP_1510 (  );
sky130_fd_sc_hd__tap_1 TAP_15100 (  );
sky130_fd_sc_hd__tap_1 TAP_15101 (  );
sky130_fd_sc_hd__tap_1 TAP_15102 (  );
sky130_fd_sc_hd__tap_1 TAP_15103 (  );
sky130_fd_sc_hd__tap_1 TAP_15104 (  );
sky130_fd_sc_hd__tap_1 TAP_15105 (  );
sky130_fd_sc_hd__tap_1 TAP_15106 (  );
sky130_fd_sc_hd__tap_1 TAP_15107 (  );
sky130_fd_sc_hd__tap_1 TAP_15108 (  );
sky130_fd_sc_hd__tap_1 TAP_15109 (  );
sky130_fd_sc_hd__tap_1 TAP_1511 (  );
sky130_fd_sc_hd__tap_1 TAP_15110 (  );
sky130_fd_sc_hd__tap_1 TAP_15111 (  );
sky130_fd_sc_hd__tap_1 TAP_15112 (  );
sky130_fd_sc_hd__tap_1 TAP_15113 (  );
sky130_fd_sc_hd__tap_1 TAP_15114 (  );
sky130_fd_sc_hd__tap_1 TAP_15115 (  );
sky130_fd_sc_hd__tap_1 TAP_15116 (  );
sky130_fd_sc_hd__tap_1 TAP_15117 (  );
sky130_fd_sc_hd__tap_1 TAP_15118 (  );
sky130_fd_sc_hd__tap_1 TAP_15119 (  );
sky130_fd_sc_hd__tap_1 TAP_1512 (  );
sky130_fd_sc_hd__tap_1 TAP_15120 (  );
sky130_fd_sc_hd__tap_1 TAP_15121 (  );
sky130_fd_sc_hd__tap_1 TAP_15122 (  );
sky130_fd_sc_hd__tap_1 TAP_15123 (  );
sky130_fd_sc_hd__tap_1 TAP_15124 (  );
sky130_fd_sc_hd__tap_1 TAP_15125 (  );
sky130_fd_sc_hd__tap_1 TAP_15126 (  );
sky130_fd_sc_hd__tap_1 TAP_15127 (  );
sky130_fd_sc_hd__tap_1 TAP_15128 (  );
sky130_fd_sc_hd__tap_1 TAP_15129 (  );
sky130_fd_sc_hd__tap_1 TAP_1513 (  );
sky130_fd_sc_hd__tap_1 TAP_15130 (  );
sky130_fd_sc_hd__tap_1 TAP_15131 (  );
sky130_fd_sc_hd__tap_1 TAP_15132 (  );
sky130_fd_sc_hd__tap_1 TAP_15133 (  );
sky130_fd_sc_hd__tap_1 TAP_15134 (  );
sky130_fd_sc_hd__tap_1 TAP_15135 (  );
sky130_fd_sc_hd__tap_1 TAP_15136 (  );
sky130_fd_sc_hd__tap_1 TAP_15137 (  );
sky130_fd_sc_hd__tap_1 TAP_15138 (  );
sky130_fd_sc_hd__tap_1 TAP_15139 (  );
sky130_fd_sc_hd__tap_1 TAP_1514 (  );
sky130_fd_sc_hd__tap_1 TAP_15140 (  );
sky130_fd_sc_hd__tap_1 TAP_15141 (  );
sky130_fd_sc_hd__tap_1 TAP_15142 (  );
sky130_fd_sc_hd__tap_1 TAP_15143 (  );
sky130_fd_sc_hd__tap_1 TAP_15144 (  );
sky130_fd_sc_hd__tap_1 TAP_15145 (  );
sky130_fd_sc_hd__tap_1 TAP_15146 (  );
sky130_fd_sc_hd__tap_1 TAP_15147 (  );
sky130_fd_sc_hd__tap_1 TAP_15148 (  );
sky130_fd_sc_hd__tap_1 TAP_15149 (  );
sky130_fd_sc_hd__tap_1 TAP_1515 (  );
sky130_fd_sc_hd__tap_1 TAP_15150 (  );
sky130_fd_sc_hd__tap_1 TAP_15151 (  );
sky130_fd_sc_hd__tap_1 TAP_15152 (  );
sky130_fd_sc_hd__tap_1 TAP_15153 (  );
sky130_fd_sc_hd__tap_1 TAP_15154 (  );
sky130_fd_sc_hd__tap_1 TAP_15155 (  );
sky130_fd_sc_hd__tap_1 TAP_15156 (  );
sky130_fd_sc_hd__tap_1 TAP_15157 (  );
sky130_fd_sc_hd__tap_1 TAP_15158 (  );
sky130_fd_sc_hd__tap_1 TAP_15159 (  );
sky130_fd_sc_hd__tap_1 TAP_1516 (  );
sky130_fd_sc_hd__tap_1 TAP_15160 (  );
sky130_fd_sc_hd__tap_1 TAP_15161 (  );
sky130_fd_sc_hd__tap_1 TAP_15162 (  );
sky130_fd_sc_hd__tap_1 TAP_15163 (  );
sky130_fd_sc_hd__tap_1 TAP_15164 (  );
sky130_fd_sc_hd__tap_1 TAP_15165 (  );
sky130_fd_sc_hd__tap_1 TAP_15166 (  );
sky130_fd_sc_hd__tap_1 TAP_15167 (  );
sky130_fd_sc_hd__tap_1 TAP_15168 (  );
sky130_fd_sc_hd__tap_1 TAP_15169 (  );
sky130_fd_sc_hd__tap_1 TAP_1517 (  );
sky130_fd_sc_hd__tap_1 TAP_15170 (  );
sky130_fd_sc_hd__tap_1 TAP_15171 (  );
sky130_fd_sc_hd__tap_1 TAP_15172 (  );
sky130_fd_sc_hd__tap_1 TAP_15173 (  );
sky130_fd_sc_hd__tap_1 TAP_15174 (  );
sky130_fd_sc_hd__tap_1 TAP_15175 (  );
sky130_fd_sc_hd__tap_1 TAP_15176 (  );
sky130_fd_sc_hd__tap_1 TAP_15177 (  );
sky130_fd_sc_hd__tap_1 TAP_15178 (  );
sky130_fd_sc_hd__tap_1 TAP_15179 (  );
sky130_fd_sc_hd__tap_1 TAP_1518 (  );
sky130_fd_sc_hd__tap_1 TAP_15180 (  );
sky130_fd_sc_hd__tap_1 TAP_15181 (  );
sky130_fd_sc_hd__tap_1 TAP_15182 (  );
sky130_fd_sc_hd__tap_1 TAP_15183 (  );
sky130_fd_sc_hd__tap_1 TAP_15184 (  );
sky130_fd_sc_hd__tap_1 TAP_15185 (  );
sky130_fd_sc_hd__tap_1 TAP_15186 (  );
sky130_fd_sc_hd__tap_1 TAP_15187 (  );
sky130_fd_sc_hd__tap_1 TAP_15188 (  );
sky130_fd_sc_hd__tap_1 TAP_15189 (  );
sky130_fd_sc_hd__tap_1 TAP_1519 (  );
sky130_fd_sc_hd__tap_1 TAP_15190 (  );
sky130_fd_sc_hd__tap_1 TAP_15191 (  );
sky130_fd_sc_hd__tap_1 TAP_15192 (  );
sky130_fd_sc_hd__tap_1 TAP_15193 (  );
sky130_fd_sc_hd__tap_1 TAP_15194 (  );
sky130_fd_sc_hd__tap_1 TAP_15195 (  );
sky130_fd_sc_hd__tap_1 TAP_15196 (  );
sky130_fd_sc_hd__tap_1 TAP_15197 (  );
sky130_fd_sc_hd__tap_1 TAP_15198 (  );
sky130_fd_sc_hd__tap_1 TAP_15199 (  );
sky130_fd_sc_hd__tap_1 TAP_1520 (  );
sky130_fd_sc_hd__tap_1 TAP_15200 (  );
sky130_fd_sc_hd__tap_1 TAP_15201 (  );
sky130_fd_sc_hd__tap_1 TAP_15202 (  );
sky130_fd_sc_hd__tap_1 TAP_15203 (  );
sky130_fd_sc_hd__tap_1 TAP_15204 (  );
sky130_fd_sc_hd__tap_1 TAP_15205 (  );
sky130_fd_sc_hd__tap_1 TAP_15206 (  );
sky130_fd_sc_hd__tap_1 TAP_15207 (  );
sky130_fd_sc_hd__tap_1 TAP_15208 (  );
sky130_fd_sc_hd__tap_1 TAP_15209 (  );
sky130_fd_sc_hd__tap_1 TAP_1521 (  );
sky130_fd_sc_hd__tap_1 TAP_15210 (  );
sky130_fd_sc_hd__tap_1 TAP_15211 (  );
sky130_fd_sc_hd__tap_1 TAP_15212 (  );
sky130_fd_sc_hd__tap_1 TAP_15213 (  );
sky130_fd_sc_hd__tap_1 TAP_15214 (  );
sky130_fd_sc_hd__tap_1 TAP_15215 (  );
sky130_fd_sc_hd__tap_1 TAP_15216 (  );
sky130_fd_sc_hd__tap_1 TAP_15217 (  );
sky130_fd_sc_hd__tap_1 TAP_15218 (  );
sky130_fd_sc_hd__tap_1 TAP_15219 (  );
sky130_fd_sc_hd__tap_1 TAP_1522 (  );
sky130_fd_sc_hd__tap_1 TAP_15220 (  );
sky130_fd_sc_hd__tap_1 TAP_15221 (  );
sky130_fd_sc_hd__tap_1 TAP_15222 (  );
sky130_fd_sc_hd__tap_1 TAP_15223 (  );
sky130_fd_sc_hd__tap_1 TAP_15224 (  );
sky130_fd_sc_hd__tap_1 TAP_15225 (  );
sky130_fd_sc_hd__tap_1 TAP_15226 (  );
sky130_fd_sc_hd__tap_1 TAP_15227 (  );
sky130_fd_sc_hd__tap_1 TAP_15228 (  );
sky130_fd_sc_hd__tap_1 TAP_15229 (  );
sky130_fd_sc_hd__tap_1 TAP_1523 (  );
sky130_fd_sc_hd__tap_1 TAP_15230 (  );
sky130_fd_sc_hd__tap_1 TAP_15231 (  );
sky130_fd_sc_hd__tap_1 TAP_15232 (  );
sky130_fd_sc_hd__tap_1 TAP_15233 (  );
sky130_fd_sc_hd__tap_1 TAP_15234 (  );
sky130_fd_sc_hd__tap_1 TAP_15235 (  );
sky130_fd_sc_hd__tap_1 TAP_15236 (  );
sky130_fd_sc_hd__tap_1 TAP_15237 (  );
sky130_fd_sc_hd__tap_1 TAP_15238 (  );
sky130_fd_sc_hd__tap_1 TAP_15239 (  );
sky130_fd_sc_hd__tap_1 TAP_1524 (  );
sky130_fd_sc_hd__tap_1 TAP_15240 (  );
sky130_fd_sc_hd__tap_1 TAP_15241 (  );
sky130_fd_sc_hd__tap_1 TAP_15242 (  );
sky130_fd_sc_hd__tap_1 TAP_15243 (  );
sky130_fd_sc_hd__tap_1 TAP_15244 (  );
sky130_fd_sc_hd__tap_1 TAP_15245 (  );
sky130_fd_sc_hd__tap_1 TAP_15246 (  );
sky130_fd_sc_hd__tap_1 TAP_15247 (  );
sky130_fd_sc_hd__tap_1 TAP_15248 (  );
sky130_fd_sc_hd__tap_1 TAP_15249 (  );
sky130_fd_sc_hd__tap_1 TAP_1525 (  );
sky130_fd_sc_hd__tap_1 TAP_15250 (  );
sky130_fd_sc_hd__tap_1 TAP_15251 (  );
sky130_fd_sc_hd__tap_1 TAP_15252 (  );
sky130_fd_sc_hd__tap_1 TAP_15253 (  );
sky130_fd_sc_hd__tap_1 TAP_15254 (  );
sky130_fd_sc_hd__tap_1 TAP_15255 (  );
sky130_fd_sc_hd__tap_1 TAP_15256 (  );
sky130_fd_sc_hd__tap_1 TAP_15257 (  );
sky130_fd_sc_hd__tap_1 TAP_15258 (  );
sky130_fd_sc_hd__tap_1 TAP_15259 (  );
sky130_fd_sc_hd__tap_1 TAP_1526 (  );
sky130_fd_sc_hd__tap_1 TAP_15260 (  );
sky130_fd_sc_hd__tap_1 TAP_15261 (  );
sky130_fd_sc_hd__tap_1 TAP_15262 (  );
sky130_fd_sc_hd__tap_1 TAP_15263 (  );
sky130_fd_sc_hd__tap_1 TAP_15264 (  );
sky130_fd_sc_hd__tap_1 TAP_15265 (  );
sky130_fd_sc_hd__tap_1 TAP_15266 (  );
sky130_fd_sc_hd__tap_1 TAP_15267 (  );
sky130_fd_sc_hd__tap_1 TAP_15268 (  );
sky130_fd_sc_hd__tap_1 TAP_15269 (  );
sky130_fd_sc_hd__tap_1 TAP_1527 (  );
sky130_fd_sc_hd__tap_1 TAP_15270 (  );
sky130_fd_sc_hd__tap_1 TAP_15271 (  );
sky130_fd_sc_hd__tap_1 TAP_15272 (  );
sky130_fd_sc_hd__tap_1 TAP_15273 (  );
sky130_fd_sc_hd__tap_1 TAP_15274 (  );
sky130_fd_sc_hd__tap_1 TAP_15275 (  );
sky130_fd_sc_hd__tap_1 TAP_15276 (  );
sky130_fd_sc_hd__tap_1 TAP_15277 (  );
sky130_fd_sc_hd__tap_1 TAP_15278 (  );
sky130_fd_sc_hd__tap_1 TAP_15279 (  );
sky130_fd_sc_hd__tap_1 TAP_1528 (  );
sky130_fd_sc_hd__tap_1 TAP_15280 (  );
sky130_fd_sc_hd__tap_1 TAP_15281 (  );
sky130_fd_sc_hd__tap_1 TAP_15282 (  );
sky130_fd_sc_hd__tap_1 TAP_15283 (  );
sky130_fd_sc_hd__tap_1 TAP_15284 (  );
sky130_fd_sc_hd__tap_1 TAP_15285 (  );
sky130_fd_sc_hd__tap_1 TAP_15286 (  );
sky130_fd_sc_hd__tap_1 TAP_15287 (  );
sky130_fd_sc_hd__tap_1 TAP_15288 (  );
sky130_fd_sc_hd__tap_1 TAP_15289 (  );
sky130_fd_sc_hd__tap_1 TAP_1529 (  );
sky130_fd_sc_hd__tap_1 TAP_15290 (  );
sky130_fd_sc_hd__tap_1 TAP_15291 (  );
sky130_fd_sc_hd__tap_1 TAP_15292 (  );
sky130_fd_sc_hd__tap_1 TAP_15293 (  );
sky130_fd_sc_hd__tap_1 TAP_15294 (  );
sky130_fd_sc_hd__tap_1 TAP_15295 (  );
sky130_fd_sc_hd__tap_1 TAP_15296 (  );
sky130_fd_sc_hd__tap_1 TAP_15297 (  );
sky130_fd_sc_hd__tap_1 TAP_15298 (  );
sky130_fd_sc_hd__tap_1 TAP_15299 (  );
sky130_fd_sc_hd__tap_1 TAP_1530 (  );
sky130_fd_sc_hd__tap_1 TAP_15300 (  );
sky130_fd_sc_hd__tap_1 TAP_15301 (  );
sky130_fd_sc_hd__tap_1 TAP_15302 (  );
sky130_fd_sc_hd__tap_1 TAP_15303 (  );
sky130_fd_sc_hd__tap_1 TAP_15304 (  );
sky130_fd_sc_hd__tap_1 TAP_15305 (  );
sky130_fd_sc_hd__tap_1 TAP_15306 (  );
sky130_fd_sc_hd__tap_1 TAP_15307 (  );
sky130_fd_sc_hd__tap_1 TAP_15308 (  );
sky130_fd_sc_hd__tap_1 TAP_1531 (  );
sky130_fd_sc_hd__tap_1 TAP_1532 (  );
sky130_fd_sc_hd__tap_1 TAP_1533 (  );
sky130_fd_sc_hd__tap_1 TAP_1534 (  );
sky130_fd_sc_hd__tap_1 TAP_1535 (  );
sky130_fd_sc_hd__tap_1 TAP_1536 (  );
sky130_fd_sc_hd__tap_1 TAP_1537 (  );
sky130_fd_sc_hd__tap_1 TAP_1538 (  );
sky130_fd_sc_hd__tap_1 TAP_1539 (  );
sky130_fd_sc_hd__tap_1 TAP_1540 (  );
sky130_fd_sc_hd__tap_1 TAP_1541 (  );
sky130_fd_sc_hd__tap_1 TAP_1542 (  );
sky130_fd_sc_hd__tap_1 TAP_1543 (  );
sky130_fd_sc_hd__tap_1 TAP_1544 (  );
sky130_fd_sc_hd__tap_1 TAP_1545 (  );
sky130_fd_sc_hd__tap_1 TAP_1546 (  );
sky130_fd_sc_hd__tap_1 TAP_1547 (  );
sky130_fd_sc_hd__tap_1 TAP_1548 (  );
sky130_fd_sc_hd__tap_1 TAP_1549 (  );
sky130_fd_sc_hd__tap_1 TAP_1550 (  );
sky130_fd_sc_hd__tap_1 TAP_1551 (  );
sky130_fd_sc_hd__tap_1 TAP_1552 (  );
sky130_fd_sc_hd__tap_1 TAP_1553 (  );
sky130_fd_sc_hd__tap_1 TAP_1554 (  );
sky130_fd_sc_hd__tap_1 TAP_1555 (  );
sky130_fd_sc_hd__tap_1 TAP_1556 (  );
sky130_fd_sc_hd__tap_1 TAP_1557 (  );
sky130_fd_sc_hd__tap_1 TAP_1558 (  );
sky130_fd_sc_hd__tap_1 TAP_1559 (  );
sky130_fd_sc_hd__tap_1 TAP_1560 (  );
sky130_fd_sc_hd__tap_1 TAP_1561 (  );
sky130_fd_sc_hd__tap_1 TAP_1562 (  );
sky130_fd_sc_hd__tap_1 TAP_1563 (  );
sky130_fd_sc_hd__tap_1 TAP_1564 (  );
sky130_fd_sc_hd__tap_1 TAP_1565 (  );
sky130_fd_sc_hd__tap_1 TAP_1566 (  );
sky130_fd_sc_hd__tap_1 TAP_1567 (  );
sky130_fd_sc_hd__tap_1 TAP_1568 (  );
sky130_fd_sc_hd__tap_1 TAP_1569 (  );
sky130_fd_sc_hd__tap_1 TAP_1570 (  );
sky130_fd_sc_hd__tap_1 TAP_1571 (  );
sky130_fd_sc_hd__tap_1 TAP_1572 (  );
sky130_fd_sc_hd__tap_1 TAP_1573 (  );
sky130_fd_sc_hd__tap_1 TAP_1574 (  );
sky130_fd_sc_hd__tap_1 TAP_1575 (  );
sky130_fd_sc_hd__tap_1 TAP_1576 (  );
sky130_fd_sc_hd__tap_1 TAP_1577 (  );
sky130_fd_sc_hd__tap_1 TAP_1578 (  );
sky130_fd_sc_hd__tap_1 TAP_1579 (  );
sky130_fd_sc_hd__tap_1 TAP_1580 (  );
sky130_fd_sc_hd__tap_1 TAP_1581 (  );
sky130_fd_sc_hd__tap_1 TAP_1582 (  );
sky130_fd_sc_hd__tap_1 TAP_1583 (  );
sky130_fd_sc_hd__tap_1 TAP_1584 (  );
sky130_fd_sc_hd__tap_1 TAP_1585 (  );
sky130_fd_sc_hd__tap_1 TAP_1586 (  );
sky130_fd_sc_hd__tap_1 TAP_1587 (  );
sky130_fd_sc_hd__tap_1 TAP_1588 (  );
sky130_fd_sc_hd__tap_1 TAP_1589 (  );
sky130_fd_sc_hd__tap_1 TAP_1590 (  );
sky130_fd_sc_hd__tap_1 TAP_1591 (  );
sky130_fd_sc_hd__tap_1 TAP_1592 (  );
sky130_fd_sc_hd__tap_1 TAP_1593 (  );
sky130_fd_sc_hd__tap_1 TAP_1594 (  );
sky130_fd_sc_hd__tap_1 TAP_1595 (  );
sky130_fd_sc_hd__tap_1 TAP_1596 (  );
sky130_fd_sc_hd__tap_1 TAP_1597 (  );
sky130_fd_sc_hd__tap_1 TAP_1598 (  );
sky130_fd_sc_hd__tap_1 TAP_1599 (  );
sky130_fd_sc_hd__tap_1 TAP_1600 (  );
sky130_fd_sc_hd__tap_1 TAP_1601 (  );
sky130_fd_sc_hd__tap_1 TAP_1602 (  );
sky130_fd_sc_hd__tap_1 TAP_1603 (  );
sky130_fd_sc_hd__tap_1 TAP_1604 (  );
sky130_fd_sc_hd__tap_1 TAP_1605 (  );
sky130_fd_sc_hd__tap_1 TAP_1606 (  );
sky130_fd_sc_hd__tap_1 TAP_1607 (  );
sky130_fd_sc_hd__tap_1 TAP_1608 (  );
sky130_fd_sc_hd__tap_1 TAP_1609 (  );
sky130_fd_sc_hd__tap_1 TAP_1610 (  );
sky130_fd_sc_hd__tap_1 TAP_1611 (  );
sky130_fd_sc_hd__tap_1 TAP_1612 (  );
sky130_fd_sc_hd__tap_1 TAP_1613 (  );
sky130_fd_sc_hd__tap_1 TAP_1614 (  );
sky130_fd_sc_hd__tap_1 TAP_1615 (  );
sky130_fd_sc_hd__tap_1 TAP_1616 (  );
sky130_fd_sc_hd__tap_1 TAP_1617 (  );
sky130_fd_sc_hd__tap_1 TAP_1618 (  );
sky130_fd_sc_hd__tap_1 TAP_1619 (  );
sky130_fd_sc_hd__tap_1 TAP_1620 (  );
sky130_fd_sc_hd__tap_1 TAP_1621 (  );
sky130_fd_sc_hd__tap_1 TAP_1622 (  );
sky130_fd_sc_hd__tap_1 TAP_1623 (  );
sky130_fd_sc_hd__tap_1 TAP_1624 (  );
sky130_fd_sc_hd__tap_1 TAP_1625 (  );
sky130_fd_sc_hd__tap_1 TAP_1626 (  );
sky130_fd_sc_hd__tap_1 TAP_1627 (  );
sky130_fd_sc_hd__tap_1 TAP_1628 (  );
sky130_fd_sc_hd__tap_1 TAP_1629 (  );
sky130_fd_sc_hd__tap_1 TAP_1630 (  );
sky130_fd_sc_hd__tap_1 TAP_1631 (  );
sky130_fd_sc_hd__tap_1 TAP_1632 (  );
sky130_fd_sc_hd__tap_1 TAP_1633 (  );
sky130_fd_sc_hd__tap_1 TAP_1634 (  );
sky130_fd_sc_hd__tap_1 TAP_1635 (  );
sky130_fd_sc_hd__tap_1 TAP_1636 (  );
sky130_fd_sc_hd__tap_1 TAP_1637 (  );
sky130_fd_sc_hd__tap_1 TAP_1638 (  );
sky130_fd_sc_hd__tap_1 TAP_1639 (  );
sky130_fd_sc_hd__tap_1 TAP_1640 (  );
sky130_fd_sc_hd__tap_1 TAP_1641 (  );
sky130_fd_sc_hd__tap_1 TAP_1642 (  );
sky130_fd_sc_hd__tap_1 TAP_1643 (  );
sky130_fd_sc_hd__tap_1 TAP_1644 (  );
sky130_fd_sc_hd__tap_1 TAP_1645 (  );
sky130_fd_sc_hd__tap_1 TAP_1646 (  );
sky130_fd_sc_hd__tap_1 TAP_1647 (  );
sky130_fd_sc_hd__tap_1 TAP_1648 (  );
sky130_fd_sc_hd__tap_1 TAP_1649 (  );
sky130_fd_sc_hd__tap_1 TAP_1650 (  );
sky130_fd_sc_hd__tap_1 TAP_1651 (  );
sky130_fd_sc_hd__tap_1 TAP_1652 (  );
sky130_fd_sc_hd__tap_1 TAP_1653 (  );
sky130_fd_sc_hd__tap_1 TAP_1654 (  );
sky130_fd_sc_hd__tap_1 TAP_1655 (  );
sky130_fd_sc_hd__tap_1 TAP_1656 (  );
sky130_fd_sc_hd__tap_1 TAP_1657 (  );
sky130_fd_sc_hd__tap_1 TAP_1658 (  );
sky130_fd_sc_hd__tap_1 TAP_1659 (  );
sky130_fd_sc_hd__tap_1 TAP_1660 (  );
sky130_fd_sc_hd__tap_1 TAP_1661 (  );
sky130_fd_sc_hd__tap_1 TAP_1662 (  );
sky130_fd_sc_hd__tap_1 TAP_1663 (  );
sky130_fd_sc_hd__tap_1 TAP_1664 (  );
sky130_fd_sc_hd__tap_1 TAP_1665 (  );
sky130_fd_sc_hd__tap_1 TAP_1666 (  );
sky130_fd_sc_hd__tap_1 TAP_1667 (  );
sky130_fd_sc_hd__tap_1 TAP_1668 (  );
sky130_fd_sc_hd__tap_1 TAP_1669 (  );
sky130_fd_sc_hd__tap_1 TAP_1670 (  );
sky130_fd_sc_hd__tap_1 TAP_1671 (  );
sky130_fd_sc_hd__tap_1 TAP_1672 (  );
sky130_fd_sc_hd__tap_1 TAP_1673 (  );
sky130_fd_sc_hd__tap_1 TAP_1674 (  );
sky130_fd_sc_hd__tap_1 TAP_1675 (  );
sky130_fd_sc_hd__tap_1 TAP_1676 (  );
sky130_fd_sc_hd__tap_1 TAP_1677 (  );
sky130_fd_sc_hd__tap_1 TAP_1678 (  );
sky130_fd_sc_hd__tap_1 TAP_1679 (  );
sky130_fd_sc_hd__tap_1 TAP_1680 (  );
sky130_fd_sc_hd__tap_1 TAP_1681 (  );
sky130_fd_sc_hd__tap_1 TAP_1682 (  );
sky130_fd_sc_hd__tap_1 TAP_1683 (  );
sky130_fd_sc_hd__tap_1 TAP_1684 (  );
sky130_fd_sc_hd__tap_1 TAP_1685 (  );
sky130_fd_sc_hd__tap_1 TAP_1686 (  );
sky130_fd_sc_hd__tap_1 TAP_1687 (  );
sky130_fd_sc_hd__tap_1 TAP_1688 (  );
sky130_fd_sc_hd__tap_1 TAP_1689 (  );
sky130_fd_sc_hd__tap_1 TAP_1690 (  );
sky130_fd_sc_hd__tap_1 TAP_1691 (  );
sky130_fd_sc_hd__tap_1 TAP_1692 (  );
sky130_fd_sc_hd__tap_1 TAP_1693 (  );
sky130_fd_sc_hd__tap_1 TAP_1694 (  );
sky130_fd_sc_hd__tap_1 TAP_1695 (  );
sky130_fd_sc_hd__tap_1 TAP_1696 (  );
sky130_fd_sc_hd__tap_1 TAP_1697 (  );
sky130_fd_sc_hd__tap_1 TAP_1698 (  );
sky130_fd_sc_hd__tap_1 TAP_1699 (  );
sky130_fd_sc_hd__tap_1 TAP_1700 (  );
sky130_fd_sc_hd__tap_1 TAP_1701 (  );
sky130_fd_sc_hd__tap_1 TAP_1702 (  );
sky130_fd_sc_hd__tap_1 TAP_1703 (  );
sky130_fd_sc_hd__tap_1 TAP_1704 (  );
sky130_fd_sc_hd__tap_1 TAP_1705 (  );
sky130_fd_sc_hd__tap_1 TAP_1706 (  );
sky130_fd_sc_hd__tap_1 TAP_1707 (  );
sky130_fd_sc_hd__tap_1 TAP_1708 (  );
sky130_fd_sc_hd__tap_1 TAP_1709 (  );
sky130_fd_sc_hd__tap_1 TAP_1710 (  );
sky130_fd_sc_hd__tap_1 TAP_1711 (  );
sky130_fd_sc_hd__tap_1 TAP_1712 (  );
sky130_fd_sc_hd__tap_1 TAP_1713 (  );
sky130_fd_sc_hd__tap_1 TAP_1714 (  );
sky130_fd_sc_hd__tap_1 TAP_1715 (  );
sky130_fd_sc_hd__tap_1 TAP_1716 (  );
sky130_fd_sc_hd__tap_1 TAP_1717 (  );
sky130_fd_sc_hd__tap_1 TAP_1718 (  );
sky130_fd_sc_hd__tap_1 TAP_1719 (  );
sky130_fd_sc_hd__tap_1 TAP_1720 (  );
sky130_fd_sc_hd__tap_1 TAP_1721 (  );
sky130_fd_sc_hd__tap_1 TAP_1722 (  );
sky130_fd_sc_hd__tap_1 TAP_1723 (  );
sky130_fd_sc_hd__tap_1 TAP_1724 (  );
sky130_fd_sc_hd__tap_1 TAP_1725 (  );
sky130_fd_sc_hd__tap_1 TAP_1726 (  );
sky130_fd_sc_hd__tap_1 TAP_1727 (  );
sky130_fd_sc_hd__tap_1 TAP_1728 (  );
sky130_fd_sc_hd__tap_1 TAP_1729 (  );
sky130_fd_sc_hd__tap_1 TAP_1730 (  );
sky130_fd_sc_hd__tap_1 TAP_1731 (  );
sky130_fd_sc_hd__tap_1 TAP_1732 (  );
sky130_fd_sc_hd__tap_1 TAP_1733 (  );
sky130_fd_sc_hd__tap_1 TAP_1734 (  );
sky130_fd_sc_hd__tap_1 TAP_1735 (  );
sky130_fd_sc_hd__tap_1 TAP_1736 (  );
sky130_fd_sc_hd__tap_1 TAP_1737 (  );
sky130_fd_sc_hd__tap_1 TAP_1738 (  );
sky130_fd_sc_hd__tap_1 TAP_1739 (  );
sky130_fd_sc_hd__tap_1 TAP_1740 (  );
sky130_fd_sc_hd__tap_1 TAP_1741 (  );
sky130_fd_sc_hd__tap_1 TAP_1742 (  );
sky130_fd_sc_hd__tap_1 TAP_1743 (  );
sky130_fd_sc_hd__tap_1 TAP_1744 (  );
sky130_fd_sc_hd__tap_1 TAP_1745 (  );
sky130_fd_sc_hd__tap_1 TAP_1746 (  );
sky130_fd_sc_hd__tap_1 TAP_1747 (  );
sky130_fd_sc_hd__tap_1 TAP_1748 (  );
sky130_fd_sc_hd__tap_1 TAP_1749 (  );
sky130_fd_sc_hd__tap_1 TAP_1750 (  );
sky130_fd_sc_hd__tap_1 TAP_1751 (  );
sky130_fd_sc_hd__tap_1 TAP_1752 (  );
sky130_fd_sc_hd__tap_1 TAP_1753 (  );
sky130_fd_sc_hd__tap_1 TAP_1754 (  );
sky130_fd_sc_hd__tap_1 TAP_1755 (  );
sky130_fd_sc_hd__tap_1 TAP_1756 (  );
sky130_fd_sc_hd__tap_1 TAP_1757 (  );
sky130_fd_sc_hd__tap_1 TAP_1758 (  );
sky130_fd_sc_hd__tap_1 TAP_1759 (  );
sky130_fd_sc_hd__tap_1 TAP_1760 (  );
sky130_fd_sc_hd__tap_1 TAP_1761 (  );
sky130_fd_sc_hd__tap_1 TAP_1762 (  );
sky130_fd_sc_hd__tap_1 TAP_1763 (  );
sky130_fd_sc_hd__tap_1 TAP_1764 (  );
sky130_fd_sc_hd__tap_1 TAP_1765 (  );
sky130_fd_sc_hd__tap_1 TAP_1766 (  );
sky130_fd_sc_hd__tap_1 TAP_1767 (  );
sky130_fd_sc_hd__tap_1 TAP_1768 (  );
sky130_fd_sc_hd__tap_1 TAP_1769 (  );
sky130_fd_sc_hd__tap_1 TAP_1770 (  );
sky130_fd_sc_hd__tap_1 TAP_1771 (  );
sky130_fd_sc_hd__tap_1 TAP_1772 (  );
sky130_fd_sc_hd__tap_1 TAP_1773 (  );
sky130_fd_sc_hd__tap_1 TAP_1774 (  );
sky130_fd_sc_hd__tap_1 TAP_1775 (  );
sky130_fd_sc_hd__tap_1 TAP_1776 (  );
sky130_fd_sc_hd__tap_1 TAP_1777 (  );
sky130_fd_sc_hd__tap_1 TAP_1778 (  );
sky130_fd_sc_hd__tap_1 TAP_1779 (  );
sky130_fd_sc_hd__tap_1 TAP_1780 (  );
sky130_fd_sc_hd__tap_1 TAP_1781 (  );
sky130_fd_sc_hd__tap_1 TAP_1782 (  );
sky130_fd_sc_hd__tap_1 TAP_1783 (  );
sky130_fd_sc_hd__tap_1 TAP_1784 (  );
sky130_fd_sc_hd__tap_1 TAP_1785 (  );
sky130_fd_sc_hd__tap_1 TAP_1786 (  );
sky130_fd_sc_hd__tap_1 TAP_1787 (  );
sky130_fd_sc_hd__tap_1 TAP_1788 (  );
sky130_fd_sc_hd__tap_1 TAP_1789 (  );
sky130_fd_sc_hd__tap_1 TAP_1790 (  );
sky130_fd_sc_hd__tap_1 TAP_1791 (  );
sky130_fd_sc_hd__tap_1 TAP_1792 (  );
sky130_fd_sc_hd__tap_1 TAP_1793 (  );
sky130_fd_sc_hd__tap_1 TAP_1794 (  );
sky130_fd_sc_hd__tap_1 TAP_1795 (  );
sky130_fd_sc_hd__tap_1 TAP_1796 (  );
sky130_fd_sc_hd__tap_1 TAP_1797 (  );
sky130_fd_sc_hd__tap_1 TAP_1798 (  );
sky130_fd_sc_hd__tap_1 TAP_1799 (  );
sky130_fd_sc_hd__tap_1 TAP_1800 (  );
sky130_fd_sc_hd__tap_1 TAP_1801 (  );
sky130_fd_sc_hd__tap_1 TAP_1802 (  );
sky130_fd_sc_hd__tap_1 TAP_1803 (  );
sky130_fd_sc_hd__tap_1 TAP_1804 (  );
sky130_fd_sc_hd__tap_1 TAP_1805 (  );
sky130_fd_sc_hd__tap_1 TAP_1806 (  );
sky130_fd_sc_hd__tap_1 TAP_1807 (  );
sky130_fd_sc_hd__tap_1 TAP_1808 (  );
sky130_fd_sc_hd__tap_1 TAP_1809 (  );
sky130_fd_sc_hd__tap_1 TAP_1810 (  );
sky130_fd_sc_hd__tap_1 TAP_1811 (  );
sky130_fd_sc_hd__tap_1 TAP_1812 (  );
sky130_fd_sc_hd__tap_1 TAP_1813 (  );
sky130_fd_sc_hd__tap_1 TAP_1814 (  );
sky130_fd_sc_hd__tap_1 TAP_1815 (  );
sky130_fd_sc_hd__tap_1 TAP_1816 (  );
sky130_fd_sc_hd__tap_1 TAP_1817 (  );
sky130_fd_sc_hd__tap_1 TAP_1818 (  );
sky130_fd_sc_hd__tap_1 TAP_1819 (  );
sky130_fd_sc_hd__tap_1 TAP_1820 (  );
sky130_fd_sc_hd__tap_1 TAP_1821 (  );
sky130_fd_sc_hd__tap_1 TAP_1822 (  );
sky130_fd_sc_hd__tap_1 TAP_1823 (  );
sky130_fd_sc_hd__tap_1 TAP_1824 (  );
sky130_fd_sc_hd__tap_1 TAP_1825 (  );
sky130_fd_sc_hd__tap_1 TAP_1826 (  );
sky130_fd_sc_hd__tap_1 TAP_1827 (  );
sky130_fd_sc_hd__tap_1 TAP_1828 (  );
sky130_fd_sc_hd__tap_1 TAP_1829 (  );
sky130_fd_sc_hd__tap_1 TAP_1830 (  );
sky130_fd_sc_hd__tap_1 TAP_1831 (  );
sky130_fd_sc_hd__tap_1 TAP_1832 (  );
sky130_fd_sc_hd__tap_1 TAP_1833 (  );
sky130_fd_sc_hd__tap_1 TAP_1834 (  );
sky130_fd_sc_hd__tap_1 TAP_1835 (  );
sky130_fd_sc_hd__tap_1 TAP_1836 (  );
sky130_fd_sc_hd__tap_1 TAP_1837 (  );
sky130_fd_sc_hd__tap_1 TAP_1838 (  );
sky130_fd_sc_hd__tap_1 TAP_1839 (  );
sky130_fd_sc_hd__tap_1 TAP_1840 (  );
sky130_fd_sc_hd__tap_1 TAP_1841 (  );
sky130_fd_sc_hd__tap_1 TAP_1842 (  );
sky130_fd_sc_hd__tap_1 TAP_1843 (  );
sky130_fd_sc_hd__tap_1 TAP_1844 (  );
sky130_fd_sc_hd__tap_1 TAP_1845 (  );
sky130_fd_sc_hd__tap_1 TAP_1846 (  );
sky130_fd_sc_hd__tap_1 TAP_1847 (  );
sky130_fd_sc_hd__tap_1 TAP_1848 (  );
sky130_fd_sc_hd__tap_1 TAP_1849 (  );
sky130_fd_sc_hd__tap_1 TAP_1850 (  );
sky130_fd_sc_hd__tap_1 TAP_1851 (  );
sky130_fd_sc_hd__tap_1 TAP_1852 (  );
sky130_fd_sc_hd__tap_1 TAP_1853 (  );
sky130_fd_sc_hd__tap_1 TAP_1854 (  );
sky130_fd_sc_hd__tap_1 TAP_1855 (  );
sky130_fd_sc_hd__tap_1 TAP_1856 (  );
sky130_fd_sc_hd__tap_1 TAP_1857 (  );
sky130_fd_sc_hd__tap_1 TAP_1858 (  );
sky130_fd_sc_hd__tap_1 TAP_1859 (  );
sky130_fd_sc_hd__tap_1 TAP_1860 (  );
sky130_fd_sc_hd__tap_1 TAP_1861 (  );
sky130_fd_sc_hd__tap_1 TAP_1862 (  );
sky130_fd_sc_hd__tap_1 TAP_1863 (  );
sky130_fd_sc_hd__tap_1 TAP_1864 (  );
sky130_fd_sc_hd__tap_1 TAP_1865 (  );
sky130_fd_sc_hd__tap_1 TAP_1866 (  );
sky130_fd_sc_hd__tap_1 TAP_1867 (  );
sky130_fd_sc_hd__tap_1 TAP_1868 (  );
sky130_fd_sc_hd__tap_1 TAP_1869 (  );
sky130_fd_sc_hd__tap_1 TAP_1870 (  );
sky130_fd_sc_hd__tap_1 TAP_1871 (  );
sky130_fd_sc_hd__tap_1 TAP_1872 (  );
sky130_fd_sc_hd__tap_1 TAP_1873 (  );
sky130_fd_sc_hd__tap_1 TAP_1874 (  );
sky130_fd_sc_hd__tap_1 TAP_1875 (  );
sky130_fd_sc_hd__tap_1 TAP_1876 (  );
sky130_fd_sc_hd__tap_1 TAP_1877 (  );
sky130_fd_sc_hd__tap_1 TAP_1878 (  );
sky130_fd_sc_hd__tap_1 TAP_1879 (  );
sky130_fd_sc_hd__tap_1 TAP_1880 (  );
sky130_fd_sc_hd__tap_1 TAP_1881 (  );
sky130_fd_sc_hd__tap_1 TAP_1882 (  );
sky130_fd_sc_hd__tap_1 TAP_1883 (  );
sky130_fd_sc_hd__tap_1 TAP_1884 (  );
sky130_fd_sc_hd__tap_1 TAP_1885 (  );
sky130_fd_sc_hd__tap_1 TAP_1886 (  );
sky130_fd_sc_hd__tap_1 TAP_1887 (  );
sky130_fd_sc_hd__tap_1 TAP_1888 (  );
sky130_fd_sc_hd__tap_1 TAP_1889 (  );
sky130_fd_sc_hd__tap_1 TAP_1890 (  );
sky130_fd_sc_hd__tap_1 TAP_1891 (  );
sky130_fd_sc_hd__tap_1 TAP_1892 (  );
sky130_fd_sc_hd__tap_1 TAP_1893 (  );
sky130_fd_sc_hd__tap_1 TAP_1894 (  );
sky130_fd_sc_hd__tap_1 TAP_1895 (  );
sky130_fd_sc_hd__tap_1 TAP_1896 (  );
sky130_fd_sc_hd__tap_1 TAP_1897 (  );
sky130_fd_sc_hd__tap_1 TAP_1898 (  );
sky130_fd_sc_hd__tap_1 TAP_1899 (  );
sky130_fd_sc_hd__tap_1 TAP_1900 (  );
sky130_fd_sc_hd__tap_1 TAP_1901 (  );
sky130_fd_sc_hd__tap_1 TAP_1902 (  );
sky130_fd_sc_hd__tap_1 TAP_1903 (  );
sky130_fd_sc_hd__tap_1 TAP_1904 (  );
sky130_fd_sc_hd__tap_1 TAP_1905 (  );
sky130_fd_sc_hd__tap_1 TAP_1906 (  );
sky130_fd_sc_hd__tap_1 TAP_1907 (  );
sky130_fd_sc_hd__tap_1 TAP_1908 (  );
sky130_fd_sc_hd__tap_1 TAP_1909 (  );
sky130_fd_sc_hd__tap_1 TAP_1910 (  );
sky130_fd_sc_hd__tap_1 TAP_1911 (  );
sky130_fd_sc_hd__tap_1 TAP_1912 (  );
sky130_fd_sc_hd__tap_1 TAP_1913 (  );
sky130_fd_sc_hd__tap_1 TAP_1914 (  );
sky130_fd_sc_hd__tap_1 TAP_1915 (  );
sky130_fd_sc_hd__tap_1 TAP_1916 (  );
sky130_fd_sc_hd__tap_1 TAP_1917 (  );
sky130_fd_sc_hd__tap_1 TAP_1918 (  );
sky130_fd_sc_hd__tap_1 TAP_1919 (  );
sky130_fd_sc_hd__tap_1 TAP_1920 (  );
sky130_fd_sc_hd__tap_1 TAP_1921 (  );
sky130_fd_sc_hd__tap_1 TAP_1922 (  );
sky130_fd_sc_hd__tap_1 TAP_1923 (  );
sky130_fd_sc_hd__tap_1 TAP_1924 (  );
sky130_fd_sc_hd__tap_1 TAP_1925 (  );
sky130_fd_sc_hd__tap_1 TAP_1926 (  );
sky130_fd_sc_hd__tap_1 TAP_1927 (  );
sky130_fd_sc_hd__tap_1 TAP_1928 (  );
sky130_fd_sc_hd__tap_1 TAP_1929 (  );
sky130_fd_sc_hd__tap_1 TAP_1930 (  );
sky130_fd_sc_hd__tap_1 TAP_1931 (  );
sky130_fd_sc_hd__tap_1 TAP_1932 (  );
sky130_fd_sc_hd__tap_1 TAP_1933 (  );
sky130_fd_sc_hd__tap_1 TAP_1934 (  );
sky130_fd_sc_hd__tap_1 TAP_1935 (  );
sky130_fd_sc_hd__tap_1 TAP_1936 (  );
sky130_fd_sc_hd__tap_1 TAP_1937 (  );
sky130_fd_sc_hd__tap_1 TAP_1938 (  );
sky130_fd_sc_hd__tap_1 TAP_1939 (  );
sky130_fd_sc_hd__tap_1 TAP_1940 (  );
sky130_fd_sc_hd__tap_1 TAP_1941 (  );
sky130_fd_sc_hd__tap_1 TAP_1942 (  );
sky130_fd_sc_hd__tap_1 TAP_1943 (  );
sky130_fd_sc_hd__tap_1 TAP_1944 (  );
sky130_fd_sc_hd__tap_1 TAP_1945 (  );
sky130_fd_sc_hd__tap_1 TAP_1946 (  );
sky130_fd_sc_hd__tap_1 TAP_1947 (  );
sky130_fd_sc_hd__tap_1 TAP_1948 (  );
sky130_fd_sc_hd__tap_1 TAP_1949 (  );
sky130_fd_sc_hd__tap_1 TAP_1950 (  );
sky130_fd_sc_hd__tap_1 TAP_1951 (  );
sky130_fd_sc_hd__tap_1 TAP_1952 (  );
sky130_fd_sc_hd__tap_1 TAP_1953 (  );
sky130_fd_sc_hd__tap_1 TAP_1954 (  );
sky130_fd_sc_hd__tap_1 TAP_1955 (  );
sky130_fd_sc_hd__tap_1 TAP_1956 (  );
sky130_fd_sc_hd__tap_1 TAP_1957 (  );
sky130_fd_sc_hd__tap_1 TAP_1958 (  );
sky130_fd_sc_hd__tap_1 TAP_1959 (  );
sky130_fd_sc_hd__tap_1 TAP_1960 (  );
sky130_fd_sc_hd__tap_1 TAP_1961 (  );
sky130_fd_sc_hd__tap_1 TAP_1962 (  );
sky130_fd_sc_hd__tap_1 TAP_1963 (  );
sky130_fd_sc_hd__tap_1 TAP_1964 (  );
sky130_fd_sc_hd__tap_1 TAP_1965 (  );
sky130_fd_sc_hd__tap_1 TAP_1966 (  );
sky130_fd_sc_hd__tap_1 TAP_1967 (  );
sky130_fd_sc_hd__tap_1 TAP_1968 (  );
sky130_fd_sc_hd__tap_1 TAP_1969 (  );
sky130_fd_sc_hd__tap_1 TAP_1970 (  );
sky130_fd_sc_hd__tap_1 TAP_1971 (  );
sky130_fd_sc_hd__tap_1 TAP_1972 (  );
sky130_fd_sc_hd__tap_1 TAP_1973 (  );
sky130_fd_sc_hd__tap_1 TAP_1974 (  );
sky130_fd_sc_hd__tap_1 TAP_1975 (  );
sky130_fd_sc_hd__tap_1 TAP_1976 (  );
sky130_fd_sc_hd__tap_1 TAP_1977 (  );
sky130_fd_sc_hd__tap_1 TAP_1978 (  );
sky130_fd_sc_hd__tap_1 TAP_1979 (  );
sky130_fd_sc_hd__tap_1 TAP_1980 (  );
sky130_fd_sc_hd__tap_1 TAP_1981 (  );
sky130_fd_sc_hd__tap_1 TAP_1982 (  );
sky130_fd_sc_hd__tap_1 TAP_1983 (  );
sky130_fd_sc_hd__tap_1 TAP_1984 (  );
sky130_fd_sc_hd__tap_1 TAP_1985 (  );
sky130_fd_sc_hd__tap_1 TAP_1986 (  );
sky130_fd_sc_hd__tap_1 TAP_1987 (  );
sky130_fd_sc_hd__tap_1 TAP_1988 (  );
sky130_fd_sc_hd__tap_1 TAP_1989 (  );
sky130_fd_sc_hd__tap_1 TAP_1990 (  );
sky130_fd_sc_hd__tap_1 TAP_1991 (  );
sky130_fd_sc_hd__tap_1 TAP_1992 (  );
sky130_fd_sc_hd__tap_1 TAP_1993 (  );
sky130_fd_sc_hd__tap_1 TAP_1994 (  );
sky130_fd_sc_hd__tap_1 TAP_1995 (  );
sky130_fd_sc_hd__tap_1 TAP_1996 (  );
sky130_fd_sc_hd__tap_1 TAP_1997 (  );
sky130_fd_sc_hd__tap_1 TAP_1998 (  );
sky130_fd_sc_hd__tap_1 TAP_1999 (  );
sky130_fd_sc_hd__tap_1 TAP_2000 (  );
sky130_fd_sc_hd__tap_1 TAP_2001 (  );
sky130_fd_sc_hd__tap_1 TAP_2002 (  );
sky130_fd_sc_hd__tap_1 TAP_2003 (  );
sky130_fd_sc_hd__tap_1 TAP_2004 (  );
sky130_fd_sc_hd__tap_1 TAP_2005 (  );
sky130_fd_sc_hd__tap_1 TAP_2006 (  );
sky130_fd_sc_hd__tap_1 TAP_2007 (  );
sky130_fd_sc_hd__tap_1 TAP_2008 (  );
sky130_fd_sc_hd__tap_1 TAP_2009 (  );
sky130_fd_sc_hd__tap_1 TAP_2010 (  );
sky130_fd_sc_hd__tap_1 TAP_2011 (  );
sky130_fd_sc_hd__tap_1 TAP_2012 (  );
sky130_fd_sc_hd__tap_1 TAP_2013 (  );
sky130_fd_sc_hd__tap_1 TAP_2014 (  );
sky130_fd_sc_hd__tap_1 TAP_2015 (  );
sky130_fd_sc_hd__tap_1 TAP_2016 (  );
sky130_fd_sc_hd__tap_1 TAP_2017 (  );
sky130_fd_sc_hd__tap_1 TAP_2018 (  );
sky130_fd_sc_hd__tap_1 TAP_2019 (  );
sky130_fd_sc_hd__tap_1 TAP_2020 (  );
sky130_fd_sc_hd__tap_1 TAP_2021 (  );
sky130_fd_sc_hd__tap_1 TAP_2022 (  );
sky130_fd_sc_hd__tap_1 TAP_2023 (  );
sky130_fd_sc_hd__tap_1 TAP_2024 (  );
sky130_fd_sc_hd__tap_1 TAP_2025 (  );
sky130_fd_sc_hd__tap_1 TAP_2026 (  );
sky130_fd_sc_hd__tap_1 TAP_2027 (  );
sky130_fd_sc_hd__tap_1 TAP_2028 (  );
sky130_fd_sc_hd__tap_1 TAP_2029 (  );
sky130_fd_sc_hd__tap_1 TAP_2030 (  );
sky130_fd_sc_hd__tap_1 TAP_2031 (  );
sky130_fd_sc_hd__tap_1 TAP_2032 (  );
sky130_fd_sc_hd__tap_1 TAP_2033 (  );
sky130_fd_sc_hd__tap_1 TAP_2034 (  );
sky130_fd_sc_hd__tap_1 TAP_2035 (  );
sky130_fd_sc_hd__tap_1 TAP_2036 (  );
sky130_fd_sc_hd__tap_1 TAP_2037 (  );
sky130_fd_sc_hd__tap_1 TAP_2038 (  );
sky130_fd_sc_hd__tap_1 TAP_2039 (  );
sky130_fd_sc_hd__tap_1 TAP_2040 (  );
sky130_fd_sc_hd__tap_1 TAP_2041 (  );
sky130_fd_sc_hd__tap_1 TAP_2042 (  );
sky130_fd_sc_hd__tap_1 TAP_2043 (  );
sky130_fd_sc_hd__tap_1 TAP_2044 (  );
sky130_fd_sc_hd__tap_1 TAP_2045 (  );
sky130_fd_sc_hd__tap_1 TAP_2046 (  );
sky130_fd_sc_hd__tap_1 TAP_2047 (  );
sky130_fd_sc_hd__tap_1 TAP_2048 (  );
sky130_fd_sc_hd__tap_1 TAP_2049 (  );
sky130_fd_sc_hd__tap_1 TAP_2050 (  );
sky130_fd_sc_hd__tap_1 TAP_2051 (  );
sky130_fd_sc_hd__tap_1 TAP_2052 (  );
sky130_fd_sc_hd__tap_1 TAP_2053 (  );
sky130_fd_sc_hd__tap_1 TAP_2054 (  );
sky130_fd_sc_hd__tap_1 TAP_2055 (  );
sky130_fd_sc_hd__tap_1 TAP_2056 (  );
sky130_fd_sc_hd__tap_1 TAP_2057 (  );
sky130_fd_sc_hd__tap_1 TAP_2058 (  );
sky130_fd_sc_hd__tap_1 TAP_2059 (  );
sky130_fd_sc_hd__tap_1 TAP_2060 (  );
sky130_fd_sc_hd__tap_1 TAP_2061 (  );
sky130_fd_sc_hd__tap_1 TAP_2062 (  );
sky130_fd_sc_hd__tap_1 TAP_2063 (  );
sky130_fd_sc_hd__tap_1 TAP_2064 (  );
sky130_fd_sc_hd__tap_1 TAP_2065 (  );
sky130_fd_sc_hd__tap_1 TAP_2066 (  );
sky130_fd_sc_hd__tap_1 TAP_2067 (  );
sky130_fd_sc_hd__tap_1 TAP_2068 (  );
sky130_fd_sc_hd__tap_1 TAP_2069 (  );
sky130_fd_sc_hd__tap_1 TAP_2070 (  );
sky130_fd_sc_hd__tap_1 TAP_2071 (  );
sky130_fd_sc_hd__tap_1 TAP_2072 (  );
sky130_fd_sc_hd__tap_1 TAP_2073 (  );
sky130_fd_sc_hd__tap_1 TAP_2074 (  );
sky130_fd_sc_hd__tap_1 TAP_2075 (  );
sky130_fd_sc_hd__tap_1 TAP_2076 (  );
sky130_fd_sc_hd__tap_1 TAP_2077 (  );
sky130_fd_sc_hd__tap_1 TAP_2078 (  );
sky130_fd_sc_hd__tap_1 TAP_2079 (  );
sky130_fd_sc_hd__tap_1 TAP_2080 (  );
sky130_fd_sc_hd__tap_1 TAP_2081 (  );
sky130_fd_sc_hd__tap_1 TAP_2082 (  );
sky130_fd_sc_hd__tap_1 TAP_2083 (  );
sky130_fd_sc_hd__tap_1 TAP_2084 (  );
sky130_fd_sc_hd__tap_1 TAP_2085 (  );
sky130_fd_sc_hd__tap_1 TAP_2086 (  );
sky130_fd_sc_hd__tap_1 TAP_2087 (  );
sky130_fd_sc_hd__tap_1 TAP_2088 (  );
sky130_fd_sc_hd__tap_1 TAP_2089 (  );
sky130_fd_sc_hd__tap_1 TAP_2090 (  );
sky130_fd_sc_hd__tap_1 TAP_2091 (  );
sky130_fd_sc_hd__tap_1 TAP_2092 (  );
sky130_fd_sc_hd__tap_1 TAP_2093 (  );
sky130_fd_sc_hd__tap_1 TAP_2094 (  );
sky130_fd_sc_hd__tap_1 TAP_2095 (  );
sky130_fd_sc_hd__tap_1 TAP_2096 (  );
sky130_fd_sc_hd__tap_1 TAP_2097 (  );
sky130_fd_sc_hd__tap_1 TAP_2098 (  );
sky130_fd_sc_hd__tap_1 TAP_2099 (  );
sky130_fd_sc_hd__tap_1 TAP_2100 (  );
sky130_fd_sc_hd__tap_1 TAP_2101 (  );
sky130_fd_sc_hd__tap_1 TAP_2102 (  );
sky130_fd_sc_hd__tap_1 TAP_2103 (  );
sky130_fd_sc_hd__tap_1 TAP_2104 (  );
sky130_fd_sc_hd__tap_1 TAP_2105 (  );
sky130_fd_sc_hd__tap_1 TAP_2106 (  );
sky130_fd_sc_hd__tap_1 TAP_2107 (  );
sky130_fd_sc_hd__tap_1 TAP_2108 (  );
sky130_fd_sc_hd__tap_1 TAP_2109 (  );
sky130_fd_sc_hd__tap_1 TAP_2110 (  );
sky130_fd_sc_hd__tap_1 TAP_2111 (  );
sky130_fd_sc_hd__tap_1 TAP_2112 (  );
sky130_fd_sc_hd__tap_1 TAP_2113 (  );
sky130_fd_sc_hd__tap_1 TAP_2114 (  );
sky130_fd_sc_hd__tap_1 TAP_2115 (  );
sky130_fd_sc_hd__tap_1 TAP_2116 (  );
sky130_fd_sc_hd__tap_1 TAP_2117 (  );
sky130_fd_sc_hd__tap_1 TAP_2118 (  );
sky130_fd_sc_hd__tap_1 TAP_2119 (  );
sky130_fd_sc_hd__tap_1 TAP_2120 (  );
sky130_fd_sc_hd__tap_1 TAP_2121 (  );
sky130_fd_sc_hd__tap_1 TAP_2122 (  );
sky130_fd_sc_hd__tap_1 TAP_2123 (  );
sky130_fd_sc_hd__tap_1 TAP_2124 (  );
sky130_fd_sc_hd__tap_1 TAP_2125 (  );
sky130_fd_sc_hd__tap_1 TAP_2126 (  );
sky130_fd_sc_hd__tap_1 TAP_2127 (  );
sky130_fd_sc_hd__tap_1 TAP_2128 (  );
sky130_fd_sc_hd__tap_1 TAP_2129 (  );
sky130_fd_sc_hd__tap_1 TAP_2130 (  );
sky130_fd_sc_hd__tap_1 TAP_2131 (  );
sky130_fd_sc_hd__tap_1 TAP_2132 (  );
sky130_fd_sc_hd__tap_1 TAP_2133 (  );
sky130_fd_sc_hd__tap_1 TAP_2134 (  );
sky130_fd_sc_hd__tap_1 TAP_2135 (  );
sky130_fd_sc_hd__tap_1 TAP_2136 (  );
sky130_fd_sc_hd__tap_1 TAP_2137 (  );
sky130_fd_sc_hd__tap_1 TAP_2138 (  );
sky130_fd_sc_hd__tap_1 TAP_2139 (  );
sky130_fd_sc_hd__tap_1 TAP_2140 (  );
sky130_fd_sc_hd__tap_1 TAP_2141 (  );
sky130_fd_sc_hd__tap_1 TAP_2142 (  );
sky130_fd_sc_hd__tap_1 TAP_2143 (  );
sky130_fd_sc_hd__tap_1 TAP_2144 (  );
sky130_fd_sc_hd__tap_1 TAP_2145 (  );
sky130_fd_sc_hd__tap_1 TAP_2146 (  );
sky130_fd_sc_hd__tap_1 TAP_2147 (  );
sky130_fd_sc_hd__tap_1 TAP_2148 (  );
sky130_fd_sc_hd__tap_1 TAP_2149 (  );
sky130_fd_sc_hd__tap_1 TAP_2150 (  );
sky130_fd_sc_hd__tap_1 TAP_2151 (  );
sky130_fd_sc_hd__tap_1 TAP_2152 (  );
sky130_fd_sc_hd__tap_1 TAP_2153 (  );
sky130_fd_sc_hd__tap_1 TAP_2154 (  );
sky130_fd_sc_hd__tap_1 TAP_2155 (  );
sky130_fd_sc_hd__tap_1 TAP_2156 (  );
sky130_fd_sc_hd__tap_1 TAP_2157 (  );
sky130_fd_sc_hd__tap_1 TAP_2158 (  );
sky130_fd_sc_hd__tap_1 TAP_2159 (  );
sky130_fd_sc_hd__tap_1 TAP_2160 (  );
sky130_fd_sc_hd__tap_1 TAP_2161 (  );
sky130_fd_sc_hd__tap_1 TAP_2162 (  );
sky130_fd_sc_hd__tap_1 TAP_2163 (  );
sky130_fd_sc_hd__tap_1 TAP_2164 (  );
sky130_fd_sc_hd__tap_1 TAP_2165 (  );
sky130_fd_sc_hd__tap_1 TAP_2166 (  );
sky130_fd_sc_hd__tap_1 TAP_2167 (  );
sky130_fd_sc_hd__tap_1 TAP_2168 (  );
sky130_fd_sc_hd__tap_1 TAP_2169 (  );
sky130_fd_sc_hd__tap_1 TAP_2170 (  );
sky130_fd_sc_hd__tap_1 TAP_2171 (  );
sky130_fd_sc_hd__tap_1 TAP_2172 (  );
sky130_fd_sc_hd__tap_1 TAP_2173 (  );
sky130_fd_sc_hd__tap_1 TAP_2174 (  );
sky130_fd_sc_hd__tap_1 TAP_2175 (  );
sky130_fd_sc_hd__tap_1 TAP_2176 (  );
sky130_fd_sc_hd__tap_1 TAP_2177 (  );
sky130_fd_sc_hd__tap_1 TAP_2178 (  );
sky130_fd_sc_hd__tap_1 TAP_2179 (  );
sky130_fd_sc_hd__tap_1 TAP_2180 (  );
sky130_fd_sc_hd__tap_1 TAP_2181 (  );
sky130_fd_sc_hd__tap_1 TAP_2182 (  );
sky130_fd_sc_hd__tap_1 TAP_2183 (  );
sky130_fd_sc_hd__tap_1 TAP_2184 (  );
sky130_fd_sc_hd__tap_1 TAP_2185 (  );
sky130_fd_sc_hd__tap_1 TAP_2186 (  );
sky130_fd_sc_hd__tap_1 TAP_2187 (  );
sky130_fd_sc_hd__tap_1 TAP_2188 (  );
sky130_fd_sc_hd__tap_1 TAP_2189 (  );
sky130_fd_sc_hd__tap_1 TAP_2190 (  );
sky130_fd_sc_hd__tap_1 TAP_2191 (  );
sky130_fd_sc_hd__tap_1 TAP_2192 (  );
sky130_fd_sc_hd__tap_1 TAP_2193 (  );
sky130_fd_sc_hd__tap_1 TAP_2194 (  );
sky130_fd_sc_hd__tap_1 TAP_2195 (  );
sky130_fd_sc_hd__tap_1 TAP_2196 (  );
sky130_fd_sc_hd__tap_1 TAP_2197 (  );
sky130_fd_sc_hd__tap_1 TAP_2198 (  );
sky130_fd_sc_hd__tap_1 TAP_2199 (  );
sky130_fd_sc_hd__tap_1 TAP_2200 (  );
sky130_fd_sc_hd__tap_1 TAP_2201 (  );
sky130_fd_sc_hd__tap_1 TAP_2202 (  );
sky130_fd_sc_hd__tap_1 TAP_2203 (  );
sky130_fd_sc_hd__tap_1 TAP_2204 (  );
sky130_fd_sc_hd__tap_1 TAP_2205 (  );
sky130_fd_sc_hd__tap_1 TAP_2206 (  );
sky130_fd_sc_hd__tap_1 TAP_2207 (  );
sky130_fd_sc_hd__tap_1 TAP_2208 (  );
sky130_fd_sc_hd__tap_1 TAP_2209 (  );
sky130_fd_sc_hd__tap_1 TAP_2210 (  );
sky130_fd_sc_hd__tap_1 TAP_2211 (  );
sky130_fd_sc_hd__tap_1 TAP_2212 (  );
sky130_fd_sc_hd__tap_1 TAP_2213 (  );
sky130_fd_sc_hd__tap_1 TAP_2214 (  );
sky130_fd_sc_hd__tap_1 TAP_2215 (  );
sky130_fd_sc_hd__tap_1 TAP_2216 (  );
sky130_fd_sc_hd__tap_1 TAP_2217 (  );
sky130_fd_sc_hd__tap_1 TAP_2218 (  );
sky130_fd_sc_hd__tap_1 TAP_2219 (  );
sky130_fd_sc_hd__tap_1 TAP_2220 (  );
sky130_fd_sc_hd__tap_1 TAP_2221 (  );
sky130_fd_sc_hd__tap_1 TAP_2222 (  );
sky130_fd_sc_hd__tap_1 TAP_2223 (  );
sky130_fd_sc_hd__tap_1 TAP_2224 (  );
sky130_fd_sc_hd__tap_1 TAP_2225 (  );
sky130_fd_sc_hd__tap_1 TAP_2226 (  );
sky130_fd_sc_hd__tap_1 TAP_2227 (  );
sky130_fd_sc_hd__tap_1 TAP_2228 (  );
sky130_fd_sc_hd__tap_1 TAP_2229 (  );
sky130_fd_sc_hd__tap_1 TAP_2230 (  );
sky130_fd_sc_hd__tap_1 TAP_2231 (  );
sky130_fd_sc_hd__tap_1 TAP_2232 (  );
sky130_fd_sc_hd__tap_1 TAP_2233 (  );
sky130_fd_sc_hd__tap_1 TAP_2234 (  );
sky130_fd_sc_hd__tap_1 TAP_2235 (  );
sky130_fd_sc_hd__tap_1 TAP_2236 (  );
sky130_fd_sc_hd__tap_1 TAP_2237 (  );
sky130_fd_sc_hd__tap_1 TAP_2238 (  );
sky130_fd_sc_hd__tap_1 TAP_2239 (  );
sky130_fd_sc_hd__tap_1 TAP_2240 (  );
sky130_fd_sc_hd__tap_1 TAP_2241 (  );
sky130_fd_sc_hd__tap_1 TAP_2242 (  );
sky130_fd_sc_hd__tap_1 TAP_2243 (  );
sky130_fd_sc_hd__tap_1 TAP_2244 (  );
sky130_fd_sc_hd__tap_1 TAP_2245 (  );
sky130_fd_sc_hd__tap_1 TAP_2246 (  );
sky130_fd_sc_hd__tap_1 TAP_2247 (  );
sky130_fd_sc_hd__tap_1 TAP_2248 (  );
sky130_fd_sc_hd__tap_1 TAP_2249 (  );
sky130_fd_sc_hd__tap_1 TAP_2250 (  );
sky130_fd_sc_hd__tap_1 TAP_2251 (  );
sky130_fd_sc_hd__tap_1 TAP_2252 (  );
sky130_fd_sc_hd__tap_1 TAP_2253 (  );
sky130_fd_sc_hd__tap_1 TAP_2254 (  );
sky130_fd_sc_hd__tap_1 TAP_2255 (  );
sky130_fd_sc_hd__tap_1 TAP_2256 (  );
sky130_fd_sc_hd__tap_1 TAP_2257 (  );
sky130_fd_sc_hd__tap_1 TAP_2258 (  );
sky130_fd_sc_hd__tap_1 TAP_2259 (  );
sky130_fd_sc_hd__tap_1 TAP_2260 (  );
sky130_fd_sc_hd__tap_1 TAP_2261 (  );
sky130_fd_sc_hd__tap_1 TAP_2262 (  );
sky130_fd_sc_hd__tap_1 TAP_2263 (  );
sky130_fd_sc_hd__tap_1 TAP_2264 (  );
sky130_fd_sc_hd__tap_1 TAP_2265 (  );
sky130_fd_sc_hd__tap_1 TAP_2266 (  );
sky130_fd_sc_hd__tap_1 TAP_2267 (  );
sky130_fd_sc_hd__tap_1 TAP_2268 (  );
sky130_fd_sc_hd__tap_1 TAP_2269 (  );
sky130_fd_sc_hd__tap_1 TAP_2270 (  );
sky130_fd_sc_hd__tap_1 TAP_2271 (  );
sky130_fd_sc_hd__tap_1 TAP_2272 (  );
sky130_fd_sc_hd__tap_1 TAP_2273 (  );
sky130_fd_sc_hd__tap_1 TAP_2274 (  );
sky130_fd_sc_hd__tap_1 TAP_2275 (  );
sky130_fd_sc_hd__tap_1 TAP_2276 (  );
sky130_fd_sc_hd__tap_1 TAP_2277 (  );
sky130_fd_sc_hd__tap_1 TAP_2278 (  );
sky130_fd_sc_hd__tap_1 TAP_2279 (  );
sky130_fd_sc_hd__tap_1 TAP_2280 (  );
sky130_fd_sc_hd__tap_1 TAP_2281 (  );
sky130_fd_sc_hd__tap_1 TAP_2282 (  );
sky130_fd_sc_hd__tap_1 TAP_2283 (  );
sky130_fd_sc_hd__tap_1 TAP_2284 (  );
sky130_fd_sc_hd__tap_1 TAP_2285 (  );
sky130_fd_sc_hd__tap_1 TAP_2286 (  );
sky130_fd_sc_hd__tap_1 TAP_2287 (  );
sky130_fd_sc_hd__tap_1 TAP_2288 (  );
sky130_fd_sc_hd__tap_1 TAP_2289 (  );
sky130_fd_sc_hd__tap_1 TAP_2290 (  );
sky130_fd_sc_hd__tap_1 TAP_2291 (  );
sky130_fd_sc_hd__tap_1 TAP_2292 (  );
sky130_fd_sc_hd__tap_1 TAP_2293 (  );
sky130_fd_sc_hd__tap_1 TAP_2294 (  );
sky130_fd_sc_hd__tap_1 TAP_2295 (  );
sky130_fd_sc_hd__tap_1 TAP_2296 (  );
sky130_fd_sc_hd__tap_1 TAP_2297 (  );
sky130_fd_sc_hd__tap_1 TAP_2298 (  );
sky130_fd_sc_hd__tap_1 TAP_2299 (  );
sky130_fd_sc_hd__tap_1 TAP_2300 (  );
sky130_fd_sc_hd__tap_1 TAP_2301 (  );
sky130_fd_sc_hd__tap_1 TAP_2302 (  );
sky130_fd_sc_hd__tap_1 TAP_2303 (  );
sky130_fd_sc_hd__tap_1 TAP_2304 (  );
sky130_fd_sc_hd__tap_1 TAP_2305 (  );
sky130_fd_sc_hd__tap_1 TAP_2306 (  );
sky130_fd_sc_hd__tap_1 TAP_2307 (  );
sky130_fd_sc_hd__tap_1 TAP_2308 (  );
sky130_fd_sc_hd__tap_1 TAP_2309 (  );
sky130_fd_sc_hd__tap_1 TAP_2310 (  );
sky130_fd_sc_hd__tap_1 TAP_2311 (  );
sky130_fd_sc_hd__tap_1 TAP_2312 (  );
sky130_fd_sc_hd__tap_1 TAP_2313 (  );
sky130_fd_sc_hd__tap_1 TAP_2314 (  );
sky130_fd_sc_hd__tap_1 TAP_2315 (  );
sky130_fd_sc_hd__tap_1 TAP_2316 (  );
sky130_fd_sc_hd__tap_1 TAP_2317 (  );
sky130_fd_sc_hd__tap_1 TAP_2318 (  );
sky130_fd_sc_hd__tap_1 TAP_2319 (  );
sky130_fd_sc_hd__tap_1 TAP_2320 (  );
sky130_fd_sc_hd__tap_1 TAP_2321 (  );
sky130_fd_sc_hd__tap_1 TAP_2322 (  );
sky130_fd_sc_hd__tap_1 TAP_2323 (  );
sky130_fd_sc_hd__tap_1 TAP_2324 (  );
sky130_fd_sc_hd__tap_1 TAP_2325 (  );
sky130_fd_sc_hd__tap_1 TAP_2326 (  );
sky130_fd_sc_hd__tap_1 TAP_2327 (  );
sky130_fd_sc_hd__tap_1 TAP_2328 (  );
sky130_fd_sc_hd__tap_1 TAP_2329 (  );
sky130_fd_sc_hd__tap_1 TAP_2330 (  );
sky130_fd_sc_hd__tap_1 TAP_2331 (  );
sky130_fd_sc_hd__tap_1 TAP_2332 (  );
sky130_fd_sc_hd__tap_1 TAP_2333 (  );
sky130_fd_sc_hd__tap_1 TAP_2334 (  );
sky130_fd_sc_hd__tap_1 TAP_2335 (  );
sky130_fd_sc_hd__tap_1 TAP_2336 (  );
sky130_fd_sc_hd__tap_1 TAP_2337 (  );
sky130_fd_sc_hd__tap_1 TAP_2338 (  );
sky130_fd_sc_hd__tap_1 TAP_2339 (  );
sky130_fd_sc_hd__tap_1 TAP_2340 (  );
sky130_fd_sc_hd__tap_1 TAP_2341 (  );
sky130_fd_sc_hd__tap_1 TAP_2342 (  );
sky130_fd_sc_hd__tap_1 TAP_2343 (  );
sky130_fd_sc_hd__tap_1 TAP_2344 (  );
sky130_fd_sc_hd__tap_1 TAP_2345 (  );
sky130_fd_sc_hd__tap_1 TAP_2346 (  );
sky130_fd_sc_hd__tap_1 TAP_2347 (  );
sky130_fd_sc_hd__tap_1 TAP_2348 (  );
sky130_fd_sc_hd__tap_1 TAP_2349 (  );
sky130_fd_sc_hd__tap_1 TAP_2350 (  );
sky130_fd_sc_hd__tap_1 TAP_2351 (  );
sky130_fd_sc_hd__tap_1 TAP_2352 (  );
sky130_fd_sc_hd__tap_1 TAP_2353 (  );
sky130_fd_sc_hd__tap_1 TAP_2354 (  );
sky130_fd_sc_hd__tap_1 TAP_2355 (  );
sky130_fd_sc_hd__tap_1 TAP_2356 (  );
sky130_fd_sc_hd__tap_1 TAP_2357 (  );
sky130_fd_sc_hd__tap_1 TAP_2358 (  );
sky130_fd_sc_hd__tap_1 TAP_2359 (  );
sky130_fd_sc_hd__tap_1 TAP_2360 (  );
sky130_fd_sc_hd__tap_1 TAP_2361 (  );
sky130_fd_sc_hd__tap_1 TAP_2362 (  );
sky130_fd_sc_hd__tap_1 TAP_2363 (  );
sky130_fd_sc_hd__tap_1 TAP_2364 (  );
sky130_fd_sc_hd__tap_1 TAP_2365 (  );
sky130_fd_sc_hd__tap_1 TAP_2366 (  );
sky130_fd_sc_hd__tap_1 TAP_2367 (  );
sky130_fd_sc_hd__tap_1 TAP_2368 (  );
sky130_fd_sc_hd__tap_1 TAP_2369 (  );
sky130_fd_sc_hd__tap_1 TAP_2370 (  );
sky130_fd_sc_hd__tap_1 TAP_2371 (  );
sky130_fd_sc_hd__tap_1 TAP_2372 (  );
sky130_fd_sc_hd__tap_1 TAP_2373 (  );
sky130_fd_sc_hd__tap_1 TAP_2374 (  );
sky130_fd_sc_hd__tap_1 TAP_2375 (  );
sky130_fd_sc_hd__tap_1 TAP_2376 (  );
sky130_fd_sc_hd__tap_1 TAP_2377 (  );
sky130_fd_sc_hd__tap_1 TAP_2378 (  );
sky130_fd_sc_hd__tap_1 TAP_2379 (  );
sky130_fd_sc_hd__tap_1 TAP_2380 (  );
sky130_fd_sc_hd__tap_1 TAP_2381 (  );
sky130_fd_sc_hd__tap_1 TAP_2382 (  );
sky130_fd_sc_hd__tap_1 TAP_2383 (  );
sky130_fd_sc_hd__tap_1 TAP_2384 (  );
sky130_fd_sc_hd__tap_1 TAP_2385 (  );
sky130_fd_sc_hd__tap_1 TAP_2386 (  );
sky130_fd_sc_hd__tap_1 TAP_2387 (  );
sky130_fd_sc_hd__tap_1 TAP_2388 (  );
sky130_fd_sc_hd__tap_1 TAP_2389 (  );
sky130_fd_sc_hd__tap_1 TAP_2390 (  );
sky130_fd_sc_hd__tap_1 TAP_2391 (  );
sky130_fd_sc_hd__tap_1 TAP_2392 (  );
sky130_fd_sc_hd__tap_1 TAP_2393 (  );
sky130_fd_sc_hd__tap_1 TAP_2394 (  );
sky130_fd_sc_hd__tap_1 TAP_2395 (  );
sky130_fd_sc_hd__tap_1 TAP_2396 (  );
sky130_fd_sc_hd__tap_1 TAP_2397 (  );
sky130_fd_sc_hd__tap_1 TAP_2398 (  );
sky130_fd_sc_hd__tap_1 TAP_2399 (  );
sky130_fd_sc_hd__tap_1 TAP_2400 (  );
sky130_fd_sc_hd__tap_1 TAP_2401 (  );
sky130_fd_sc_hd__tap_1 TAP_2402 (  );
sky130_fd_sc_hd__tap_1 TAP_2403 (  );
sky130_fd_sc_hd__tap_1 TAP_2404 (  );
sky130_fd_sc_hd__tap_1 TAP_2405 (  );
sky130_fd_sc_hd__tap_1 TAP_2406 (  );
sky130_fd_sc_hd__tap_1 TAP_2407 (  );
sky130_fd_sc_hd__tap_1 TAP_2408 (  );
sky130_fd_sc_hd__tap_1 TAP_2409 (  );
sky130_fd_sc_hd__tap_1 TAP_2410 (  );
sky130_fd_sc_hd__tap_1 TAP_2411 (  );
sky130_fd_sc_hd__tap_1 TAP_2412 (  );
sky130_fd_sc_hd__tap_1 TAP_2413 (  );
sky130_fd_sc_hd__tap_1 TAP_2414 (  );
sky130_fd_sc_hd__tap_1 TAP_2415 (  );
sky130_fd_sc_hd__tap_1 TAP_2416 (  );
sky130_fd_sc_hd__tap_1 TAP_2417 (  );
sky130_fd_sc_hd__tap_1 TAP_2418 (  );
sky130_fd_sc_hd__tap_1 TAP_2419 (  );
sky130_fd_sc_hd__tap_1 TAP_2420 (  );
sky130_fd_sc_hd__tap_1 TAP_2421 (  );
sky130_fd_sc_hd__tap_1 TAP_2422 (  );
sky130_fd_sc_hd__tap_1 TAP_2423 (  );
sky130_fd_sc_hd__tap_1 TAP_2424 (  );
sky130_fd_sc_hd__tap_1 TAP_2425 (  );
sky130_fd_sc_hd__tap_1 TAP_2426 (  );
sky130_fd_sc_hd__tap_1 TAP_2427 (  );
sky130_fd_sc_hd__tap_1 TAP_2428 (  );
sky130_fd_sc_hd__tap_1 TAP_2429 (  );
sky130_fd_sc_hd__tap_1 TAP_2430 (  );
sky130_fd_sc_hd__tap_1 TAP_2431 (  );
sky130_fd_sc_hd__tap_1 TAP_2432 (  );
sky130_fd_sc_hd__tap_1 TAP_2433 (  );
sky130_fd_sc_hd__tap_1 TAP_2434 (  );
sky130_fd_sc_hd__tap_1 TAP_2435 (  );
sky130_fd_sc_hd__tap_1 TAP_2436 (  );
sky130_fd_sc_hd__tap_1 TAP_2437 (  );
sky130_fd_sc_hd__tap_1 TAP_2438 (  );
sky130_fd_sc_hd__tap_1 TAP_2439 (  );
sky130_fd_sc_hd__tap_1 TAP_2440 (  );
sky130_fd_sc_hd__tap_1 TAP_2441 (  );
sky130_fd_sc_hd__tap_1 TAP_2442 (  );
sky130_fd_sc_hd__tap_1 TAP_2443 (  );
sky130_fd_sc_hd__tap_1 TAP_2444 (  );
sky130_fd_sc_hd__tap_1 TAP_2445 (  );
sky130_fd_sc_hd__tap_1 TAP_2446 (  );
sky130_fd_sc_hd__tap_1 TAP_2447 (  );
sky130_fd_sc_hd__tap_1 TAP_2448 (  );
sky130_fd_sc_hd__tap_1 TAP_2449 (  );
sky130_fd_sc_hd__tap_1 TAP_2450 (  );
sky130_fd_sc_hd__tap_1 TAP_2451 (  );
sky130_fd_sc_hd__tap_1 TAP_2452 (  );
sky130_fd_sc_hd__tap_1 TAP_2453 (  );
sky130_fd_sc_hd__tap_1 TAP_2454 (  );
sky130_fd_sc_hd__tap_1 TAP_2455 (  );
sky130_fd_sc_hd__tap_1 TAP_2456 (  );
sky130_fd_sc_hd__tap_1 TAP_2457 (  );
sky130_fd_sc_hd__tap_1 TAP_2458 (  );
sky130_fd_sc_hd__tap_1 TAP_2459 (  );
sky130_fd_sc_hd__tap_1 TAP_2460 (  );
sky130_fd_sc_hd__tap_1 TAP_2461 (  );
sky130_fd_sc_hd__tap_1 TAP_2462 (  );
sky130_fd_sc_hd__tap_1 TAP_2463 (  );
sky130_fd_sc_hd__tap_1 TAP_2464 (  );
sky130_fd_sc_hd__tap_1 TAP_2465 (  );
sky130_fd_sc_hd__tap_1 TAP_2466 (  );
sky130_fd_sc_hd__tap_1 TAP_2467 (  );
sky130_fd_sc_hd__tap_1 TAP_2468 (  );
sky130_fd_sc_hd__tap_1 TAP_2469 (  );
sky130_fd_sc_hd__tap_1 TAP_2470 (  );
sky130_fd_sc_hd__tap_1 TAP_2471 (  );
sky130_fd_sc_hd__tap_1 TAP_2472 (  );
sky130_fd_sc_hd__tap_1 TAP_2473 (  );
sky130_fd_sc_hd__tap_1 TAP_2474 (  );
sky130_fd_sc_hd__tap_1 TAP_2475 (  );
sky130_fd_sc_hd__tap_1 TAP_2476 (  );
sky130_fd_sc_hd__tap_1 TAP_2477 (  );
sky130_fd_sc_hd__tap_1 TAP_2478 (  );
sky130_fd_sc_hd__tap_1 TAP_2479 (  );
sky130_fd_sc_hd__tap_1 TAP_2480 (  );
sky130_fd_sc_hd__tap_1 TAP_2481 (  );
sky130_fd_sc_hd__tap_1 TAP_2482 (  );
sky130_fd_sc_hd__tap_1 TAP_2483 (  );
sky130_fd_sc_hd__tap_1 TAP_2484 (  );
sky130_fd_sc_hd__tap_1 TAP_2485 (  );
sky130_fd_sc_hd__tap_1 TAP_2486 (  );
sky130_fd_sc_hd__tap_1 TAP_2487 (  );
sky130_fd_sc_hd__tap_1 TAP_2488 (  );
sky130_fd_sc_hd__tap_1 TAP_2489 (  );
sky130_fd_sc_hd__tap_1 TAP_2490 (  );
sky130_fd_sc_hd__tap_1 TAP_2491 (  );
sky130_fd_sc_hd__tap_1 TAP_2492 (  );
sky130_fd_sc_hd__tap_1 TAP_2493 (  );
sky130_fd_sc_hd__tap_1 TAP_2494 (  );
sky130_fd_sc_hd__tap_1 TAP_2495 (  );
sky130_fd_sc_hd__tap_1 TAP_2496 (  );
sky130_fd_sc_hd__tap_1 TAP_2497 (  );
sky130_fd_sc_hd__tap_1 TAP_2498 (  );
sky130_fd_sc_hd__tap_1 TAP_2499 (  );
sky130_fd_sc_hd__tap_1 TAP_2500 (  );
sky130_fd_sc_hd__tap_1 TAP_2501 (  );
sky130_fd_sc_hd__tap_1 TAP_2502 (  );
sky130_fd_sc_hd__tap_1 TAP_2503 (  );
sky130_fd_sc_hd__tap_1 TAP_2504 (  );
sky130_fd_sc_hd__tap_1 TAP_2505 (  );
sky130_fd_sc_hd__tap_1 TAP_2506 (  );
sky130_fd_sc_hd__tap_1 TAP_2507 (  );
sky130_fd_sc_hd__tap_1 TAP_2508 (  );
sky130_fd_sc_hd__tap_1 TAP_2509 (  );
sky130_fd_sc_hd__tap_1 TAP_2510 (  );
sky130_fd_sc_hd__tap_1 TAP_2511 (  );
sky130_fd_sc_hd__tap_1 TAP_2512 (  );
sky130_fd_sc_hd__tap_1 TAP_2513 (  );
sky130_fd_sc_hd__tap_1 TAP_2514 (  );
sky130_fd_sc_hd__tap_1 TAP_2515 (  );
sky130_fd_sc_hd__tap_1 TAP_2516 (  );
sky130_fd_sc_hd__tap_1 TAP_2517 (  );
sky130_fd_sc_hd__tap_1 TAP_2518 (  );
sky130_fd_sc_hd__tap_1 TAP_2519 (  );
sky130_fd_sc_hd__tap_1 TAP_2520 (  );
sky130_fd_sc_hd__tap_1 TAP_2521 (  );
sky130_fd_sc_hd__tap_1 TAP_2522 (  );
sky130_fd_sc_hd__tap_1 TAP_2523 (  );
sky130_fd_sc_hd__tap_1 TAP_2524 (  );
sky130_fd_sc_hd__tap_1 TAP_2525 (  );
sky130_fd_sc_hd__tap_1 TAP_2526 (  );
sky130_fd_sc_hd__tap_1 TAP_2527 (  );
sky130_fd_sc_hd__tap_1 TAP_2528 (  );
sky130_fd_sc_hd__tap_1 TAP_2529 (  );
sky130_fd_sc_hd__tap_1 TAP_2530 (  );
sky130_fd_sc_hd__tap_1 TAP_2531 (  );
sky130_fd_sc_hd__tap_1 TAP_2532 (  );
sky130_fd_sc_hd__tap_1 TAP_2533 (  );
sky130_fd_sc_hd__tap_1 TAP_2534 (  );
sky130_fd_sc_hd__tap_1 TAP_2535 (  );
sky130_fd_sc_hd__tap_1 TAP_2536 (  );
sky130_fd_sc_hd__tap_1 TAP_2537 (  );
sky130_fd_sc_hd__tap_1 TAP_2538 (  );
sky130_fd_sc_hd__tap_1 TAP_2539 (  );
sky130_fd_sc_hd__tap_1 TAP_2540 (  );
sky130_fd_sc_hd__tap_1 TAP_2541 (  );
sky130_fd_sc_hd__tap_1 TAP_2542 (  );
sky130_fd_sc_hd__tap_1 TAP_2543 (  );
sky130_fd_sc_hd__tap_1 TAP_2544 (  );
sky130_fd_sc_hd__tap_1 TAP_2545 (  );
sky130_fd_sc_hd__tap_1 TAP_2546 (  );
sky130_fd_sc_hd__tap_1 TAP_2547 (  );
sky130_fd_sc_hd__tap_1 TAP_2548 (  );
sky130_fd_sc_hd__tap_1 TAP_2549 (  );
sky130_fd_sc_hd__tap_1 TAP_2550 (  );
sky130_fd_sc_hd__tap_1 TAP_2551 (  );
sky130_fd_sc_hd__tap_1 TAP_2552 (  );
sky130_fd_sc_hd__tap_1 TAP_2553 (  );
sky130_fd_sc_hd__tap_1 TAP_2554 (  );
sky130_fd_sc_hd__tap_1 TAP_2555 (  );
sky130_fd_sc_hd__tap_1 TAP_2556 (  );
sky130_fd_sc_hd__tap_1 TAP_2557 (  );
sky130_fd_sc_hd__tap_1 TAP_2558 (  );
sky130_fd_sc_hd__tap_1 TAP_2559 (  );
sky130_fd_sc_hd__tap_1 TAP_2560 (  );
sky130_fd_sc_hd__tap_1 TAP_2561 (  );
sky130_fd_sc_hd__tap_1 TAP_2562 (  );
sky130_fd_sc_hd__tap_1 TAP_2563 (  );
sky130_fd_sc_hd__tap_1 TAP_2564 (  );
sky130_fd_sc_hd__tap_1 TAP_2565 (  );
sky130_fd_sc_hd__tap_1 TAP_2566 (  );
sky130_fd_sc_hd__tap_1 TAP_2567 (  );
sky130_fd_sc_hd__tap_1 TAP_2568 (  );
sky130_fd_sc_hd__tap_1 TAP_2569 (  );
sky130_fd_sc_hd__tap_1 TAP_2570 (  );
sky130_fd_sc_hd__tap_1 TAP_2571 (  );
sky130_fd_sc_hd__tap_1 TAP_2572 (  );
sky130_fd_sc_hd__tap_1 TAP_2573 (  );
sky130_fd_sc_hd__tap_1 TAP_2574 (  );
sky130_fd_sc_hd__tap_1 TAP_2575 (  );
sky130_fd_sc_hd__tap_1 TAP_2576 (  );
sky130_fd_sc_hd__tap_1 TAP_2577 (  );
sky130_fd_sc_hd__tap_1 TAP_2578 (  );
sky130_fd_sc_hd__tap_1 TAP_2579 (  );
sky130_fd_sc_hd__tap_1 TAP_2580 (  );
sky130_fd_sc_hd__tap_1 TAP_2581 (  );
sky130_fd_sc_hd__tap_1 TAP_2582 (  );
sky130_fd_sc_hd__tap_1 TAP_2583 (  );
sky130_fd_sc_hd__tap_1 TAP_2584 (  );
sky130_fd_sc_hd__tap_1 TAP_2585 (  );
sky130_fd_sc_hd__tap_1 TAP_2586 (  );
sky130_fd_sc_hd__tap_1 TAP_2587 (  );
sky130_fd_sc_hd__tap_1 TAP_2588 (  );
sky130_fd_sc_hd__tap_1 TAP_2589 (  );
sky130_fd_sc_hd__tap_1 TAP_2590 (  );
sky130_fd_sc_hd__tap_1 TAP_2591 (  );
sky130_fd_sc_hd__tap_1 TAP_2592 (  );
sky130_fd_sc_hd__tap_1 TAP_2593 (  );
sky130_fd_sc_hd__tap_1 TAP_2594 (  );
sky130_fd_sc_hd__tap_1 TAP_2595 (  );
sky130_fd_sc_hd__tap_1 TAP_2596 (  );
sky130_fd_sc_hd__tap_1 TAP_2597 (  );
sky130_fd_sc_hd__tap_1 TAP_2598 (  );
sky130_fd_sc_hd__tap_1 TAP_2599 (  );
sky130_fd_sc_hd__tap_1 TAP_2600 (  );
sky130_fd_sc_hd__tap_1 TAP_2601 (  );
sky130_fd_sc_hd__tap_1 TAP_2602 (  );
sky130_fd_sc_hd__tap_1 TAP_2603 (  );
sky130_fd_sc_hd__tap_1 TAP_2604 (  );
sky130_fd_sc_hd__tap_1 TAP_2605 (  );
sky130_fd_sc_hd__tap_1 TAP_2606 (  );
sky130_fd_sc_hd__tap_1 TAP_2607 (  );
sky130_fd_sc_hd__tap_1 TAP_2608 (  );
sky130_fd_sc_hd__tap_1 TAP_2609 (  );
sky130_fd_sc_hd__tap_1 TAP_2610 (  );
sky130_fd_sc_hd__tap_1 TAP_2611 (  );
sky130_fd_sc_hd__tap_1 TAP_2612 (  );
sky130_fd_sc_hd__tap_1 TAP_2613 (  );
sky130_fd_sc_hd__tap_1 TAP_2614 (  );
sky130_fd_sc_hd__tap_1 TAP_2615 (  );
sky130_fd_sc_hd__tap_1 TAP_2616 (  );
sky130_fd_sc_hd__tap_1 TAP_2617 (  );
sky130_fd_sc_hd__tap_1 TAP_2618 (  );
sky130_fd_sc_hd__tap_1 TAP_2619 (  );
sky130_fd_sc_hd__tap_1 TAP_2620 (  );
sky130_fd_sc_hd__tap_1 TAP_2621 (  );
sky130_fd_sc_hd__tap_1 TAP_2622 (  );
sky130_fd_sc_hd__tap_1 TAP_2623 (  );
sky130_fd_sc_hd__tap_1 TAP_2624 (  );
sky130_fd_sc_hd__tap_1 TAP_2625 (  );
sky130_fd_sc_hd__tap_1 TAP_2626 (  );
sky130_fd_sc_hd__tap_1 TAP_2627 (  );
sky130_fd_sc_hd__tap_1 TAP_2628 (  );
sky130_fd_sc_hd__tap_1 TAP_2629 (  );
sky130_fd_sc_hd__tap_1 TAP_2630 (  );
sky130_fd_sc_hd__tap_1 TAP_2631 (  );
sky130_fd_sc_hd__tap_1 TAP_2632 (  );
sky130_fd_sc_hd__tap_1 TAP_2633 (  );
sky130_fd_sc_hd__tap_1 TAP_2634 (  );
sky130_fd_sc_hd__tap_1 TAP_2635 (  );
sky130_fd_sc_hd__tap_1 TAP_2636 (  );
sky130_fd_sc_hd__tap_1 TAP_2637 (  );
sky130_fd_sc_hd__tap_1 TAP_2638 (  );
sky130_fd_sc_hd__tap_1 TAP_2639 (  );
sky130_fd_sc_hd__tap_1 TAP_2640 (  );
sky130_fd_sc_hd__tap_1 TAP_2641 (  );
sky130_fd_sc_hd__tap_1 TAP_2642 (  );
sky130_fd_sc_hd__tap_1 TAP_2643 (  );
sky130_fd_sc_hd__tap_1 TAP_2644 (  );
sky130_fd_sc_hd__tap_1 TAP_2645 (  );
sky130_fd_sc_hd__tap_1 TAP_2646 (  );
sky130_fd_sc_hd__tap_1 TAP_2647 (  );
sky130_fd_sc_hd__tap_1 TAP_2648 (  );
sky130_fd_sc_hd__tap_1 TAP_2649 (  );
sky130_fd_sc_hd__tap_1 TAP_2650 (  );
sky130_fd_sc_hd__tap_1 TAP_2651 (  );
sky130_fd_sc_hd__tap_1 TAP_2652 (  );
sky130_fd_sc_hd__tap_1 TAP_2653 (  );
sky130_fd_sc_hd__tap_1 TAP_2654 (  );
sky130_fd_sc_hd__tap_1 TAP_2655 (  );
sky130_fd_sc_hd__tap_1 TAP_2656 (  );
sky130_fd_sc_hd__tap_1 TAP_2657 (  );
sky130_fd_sc_hd__tap_1 TAP_2658 (  );
sky130_fd_sc_hd__tap_1 TAP_2659 (  );
sky130_fd_sc_hd__tap_1 TAP_2660 (  );
sky130_fd_sc_hd__tap_1 TAP_2661 (  );
sky130_fd_sc_hd__tap_1 TAP_2662 (  );
sky130_fd_sc_hd__tap_1 TAP_2663 (  );
sky130_fd_sc_hd__tap_1 TAP_2664 (  );
sky130_fd_sc_hd__tap_1 TAP_2665 (  );
sky130_fd_sc_hd__tap_1 TAP_2666 (  );
sky130_fd_sc_hd__tap_1 TAP_2667 (  );
sky130_fd_sc_hd__tap_1 TAP_2668 (  );
sky130_fd_sc_hd__tap_1 TAP_2669 (  );
sky130_fd_sc_hd__tap_1 TAP_2670 (  );
sky130_fd_sc_hd__tap_1 TAP_2671 (  );
sky130_fd_sc_hd__tap_1 TAP_2672 (  );
sky130_fd_sc_hd__tap_1 TAP_2673 (  );
sky130_fd_sc_hd__tap_1 TAP_2674 (  );
sky130_fd_sc_hd__tap_1 TAP_2675 (  );
sky130_fd_sc_hd__tap_1 TAP_2676 (  );
sky130_fd_sc_hd__tap_1 TAP_2677 (  );
sky130_fd_sc_hd__tap_1 TAP_2678 (  );
sky130_fd_sc_hd__tap_1 TAP_2679 (  );
sky130_fd_sc_hd__tap_1 TAP_2680 (  );
sky130_fd_sc_hd__tap_1 TAP_2681 (  );
sky130_fd_sc_hd__tap_1 TAP_2682 (  );
sky130_fd_sc_hd__tap_1 TAP_2683 (  );
sky130_fd_sc_hd__tap_1 TAP_2684 (  );
sky130_fd_sc_hd__tap_1 TAP_2685 (  );
sky130_fd_sc_hd__tap_1 TAP_2686 (  );
sky130_fd_sc_hd__tap_1 TAP_2687 (  );
sky130_fd_sc_hd__tap_1 TAP_2688 (  );
sky130_fd_sc_hd__tap_1 TAP_2689 (  );
sky130_fd_sc_hd__tap_1 TAP_2690 (  );
sky130_fd_sc_hd__tap_1 TAP_2691 (  );
sky130_fd_sc_hd__tap_1 TAP_2692 (  );
sky130_fd_sc_hd__tap_1 TAP_2693 (  );
sky130_fd_sc_hd__tap_1 TAP_2694 (  );
sky130_fd_sc_hd__tap_1 TAP_2695 (  );
sky130_fd_sc_hd__tap_1 TAP_2696 (  );
sky130_fd_sc_hd__tap_1 TAP_2697 (  );
sky130_fd_sc_hd__tap_1 TAP_2698 (  );
sky130_fd_sc_hd__tap_1 TAP_2699 (  );
sky130_fd_sc_hd__tap_1 TAP_2700 (  );
sky130_fd_sc_hd__tap_1 TAP_2701 (  );
sky130_fd_sc_hd__tap_1 TAP_2702 (  );
sky130_fd_sc_hd__tap_1 TAP_2703 (  );
sky130_fd_sc_hd__tap_1 TAP_2704 (  );
sky130_fd_sc_hd__tap_1 TAP_2705 (  );
sky130_fd_sc_hd__tap_1 TAP_2706 (  );
sky130_fd_sc_hd__tap_1 TAP_2707 (  );
sky130_fd_sc_hd__tap_1 TAP_2708 (  );
sky130_fd_sc_hd__tap_1 TAP_2709 (  );
sky130_fd_sc_hd__tap_1 TAP_2710 (  );
sky130_fd_sc_hd__tap_1 TAP_2711 (  );
sky130_fd_sc_hd__tap_1 TAP_2712 (  );
sky130_fd_sc_hd__tap_1 TAP_2713 (  );
sky130_fd_sc_hd__tap_1 TAP_2714 (  );
sky130_fd_sc_hd__tap_1 TAP_2715 (  );
sky130_fd_sc_hd__tap_1 TAP_2716 (  );
sky130_fd_sc_hd__tap_1 TAP_2717 (  );
sky130_fd_sc_hd__tap_1 TAP_2718 (  );
sky130_fd_sc_hd__tap_1 TAP_2719 (  );
sky130_fd_sc_hd__tap_1 TAP_2720 (  );
sky130_fd_sc_hd__tap_1 TAP_2721 (  );
sky130_fd_sc_hd__tap_1 TAP_2722 (  );
sky130_fd_sc_hd__tap_1 TAP_2723 (  );
sky130_fd_sc_hd__tap_1 TAP_2724 (  );
sky130_fd_sc_hd__tap_1 TAP_2725 (  );
sky130_fd_sc_hd__tap_1 TAP_2726 (  );
sky130_fd_sc_hd__tap_1 TAP_2727 (  );
sky130_fd_sc_hd__tap_1 TAP_2728 (  );
sky130_fd_sc_hd__tap_1 TAP_2729 (  );
sky130_fd_sc_hd__tap_1 TAP_2730 (  );
sky130_fd_sc_hd__tap_1 TAP_2731 (  );
sky130_fd_sc_hd__tap_1 TAP_2732 (  );
sky130_fd_sc_hd__tap_1 TAP_2733 (  );
sky130_fd_sc_hd__tap_1 TAP_2734 (  );
sky130_fd_sc_hd__tap_1 TAP_2735 (  );
sky130_fd_sc_hd__tap_1 TAP_2736 (  );
sky130_fd_sc_hd__tap_1 TAP_2737 (  );
sky130_fd_sc_hd__tap_1 TAP_2738 (  );
sky130_fd_sc_hd__tap_1 TAP_2739 (  );
sky130_fd_sc_hd__tap_1 TAP_2740 (  );
sky130_fd_sc_hd__tap_1 TAP_2741 (  );
sky130_fd_sc_hd__tap_1 TAP_2742 (  );
sky130_fd_sc_hd__tap_1 TAP_2743 (  );
sky130_fd_sc_hd__tap_1 TAP_2744 (  );
sky130_fd_sc_hd__tap_1 TAP_2745 (  );
sky130_fd_sc_hd__tap_1 TAP_2746 (  );
sky130_fd_sc_hd__tap_1 TAP_2747 (  );
sky130_fd_sc_hd__tap_1 TAP_2748 (  );
sky130_fd_sc_hd__tap_1 TAP_2749 (  );
sky130_fd_sc_hd__tap_1 TAP_2750 (  );
sky130_fd_sc_hd__tap_1 TAP_2751 (  );
sky130_fd_sc_hd__tap_1 TAP_2752 (  );
sky130_fd_sc_hd__tap_1 TAP_2753 (  );
sky130_fd_sc_hd__tap_1 TAP_2754 (  );
sky130_fd_sc_hd__tap_1 TAP_2755 (  );
sky130_fd_sc_hd__tap_1 TAP_2756 (  );
sky130_fd_sc_hd__tap_1 TAP_2757 (  );
sky130_fd_sc_hd__tap_1 TAP_2758 (  );
sky130_fd_sc_hd__tap_1 TAP_2759 (  );
sky130_fd_sc_hd__tap_1 TAP_2760 (  );
sky130_fd_sc_hd__tap_1 TAP_2761 (  );
sky130_fd_sc_hd__tap_1 TAP_2762 (  );
sky130_fd_sc_hd__tap_1 TAP_2763 (  );
sky130_fd_sc_hd__tap_1 TAP_2764 (  );
sky130_fd_sc_hd__tap_1 TAP_2765 (  );
sky130_fd_sc_hd__tap_1 TAP_2766 (  );
sky130_fd_sc_hd__tap_1 TAP_2767 (  );
sky130_fd_sc_hd__tap_1 TAP_2768 (  );
sky130_fd_sc_hd__tap_1 TAP_2769 (  );
sky130_fd_sc_hd__tap_1 TAP_2770 (  );
sky130_fd_sc_hd__tap_1 TAP_2771 (  );
sky130_fd_sc_hd__tap_1 TAP_2772 (  );
sky130_fd_sc_hd__tap_1 TAP_2773 (  );
sky130_fd_sc_hd__tap_1 TAP_2774 (  );
sky130_fd_sc_hd__tap_1 TAP_2775 (  );
sky130_fd_sc_hd__tap_1 TAP_2776 (  );
sky130_fd_sc_hd__tap_1 TAP_2777 (  );
sky130_fd_sc_hd__tap_1 TAP_2778 (  );
sky130_fd_sc_hd__tap_1 TAP_2779 (  );
sky130_fd_sc_hd__tap_1 TAP_2780 (  );
sky130_fd_sc_hd__tap_1 TAP_2781 (  );
sky130_fd_sc_hd__tap_1 TAP_2782 (  );
sky130_fd_sc_hd__tap_1 TAP_2783 (  );
sky130_fd_sc_hd__tap_1 TAP_2784 (  );
sky130_fd_sc_hd__tap_1 TAP_2785 (  );
sky130_fd_sc_hd__tap_1 TAP_2786 (  );
sky130_fd_sc_hd__tap_1 TAP_2787 (  );
sky130_fd_sc_hd__tap_1 TAP_2788 (  );
sky130_fd_sc_hd__tap_1 TAP_2789 (  );
sky130_fd_sc_hd__tap_1 TAP_2790 (  );
sky130_fd_sc_hd__tap_1 TAP_2791 (  );
sky130_fd_sc_hd__tap_1 TAP_2792 (  );
sky130_fd_sc_hd__tap_1 TAP_2793 (  );
sky130_fd_sc_hd__tap_1 TAP_2794 (  );
sky130_fd_sc_hd__tap_1 TAP_2795 (  );
sky130_fd_sc_hd__tap_1 TAP_2796 (  );
sky130_fd_sc_hd__tap_1 TAP_2797 (  );
sky130_fd_sc_hd__tap_1 TAP_2798 (  );
sky130_fd_sc_hd__tap_1 TAP_2799 (  );
sky130_fd_sc_hd__tap_1 TAP_2800 (  );
sky130_fd_sc_hd__tap_1 TAP_2801 (  );
sky130_fd_sc_hd__tap_1 TAP_2802 (  );
sky130_fd_sc_hd__tap_1 TAP_2803 (  );
sky130_fd_sc_hd__tap_1 TAP_2804 (  );
sky130_fd_sc_hd__tap_1 TAP_2805 (  );
sky130_fd_sc_hd__tap_1 TAP_2806 (  );
sky130_fd_sc_hd__tap_1 TAP_2807 (  );
sky130_fd_sc_hd__tap_1 TAP_2808 (  );
sky130_fd_sc_hd__tap_1 TAP_2809 (  );
sky130_fd_sc_hd__tap_1 TAP_2810 (  );
sky130_fd_sc_hd__tap_1 TAP_2811 (  );
sky130_fd_sc_hd__tap_1 TAP_2812 (  );
sky130_fd_sc_hd__tap_1 TAP_2813 (  );
sky130_fd_sc_hd__tap_1 TAP_2814 (  );
sky130_fd_sc_hd__tap_1 TAP_2815 (  );
sky130_fd_sc_hd__tap_1 TAP_2816 (  );
sky130_fd_sc_hd__tap_1 TAP_2817 (  );
sky130_fd_sc_hd__tap_1 TAP_2818 (  );
sky130_fd_sc_hd__tap_1 TAP_2819 (  );
sky130_fd_sc_hd__tap_1 TAP_2820 (  );
sky130_fd_sc_hd__tap_1 TAP_2821 (  );
sky130_fd_sc_hd__tap_1 TAP_2822 (  );
sky130_fd_sc_hd__tap_1 TAP_2823 (  );
sky130_fd_sc_hd__tap_1 TAP_2824 (  );
sky130_fd_sc_hd__tap_1 TAP_2825 (  );
sky130_fd_sc_hd__tap_1 TAP_2826 (  );
sky130_fd_sc_hd__tap_1 TAP_2827 (  );
sky130_fd_sc_hd__tap_1 TAP_2828 (  );
sky130_fd_sc_hd__tap_1 TAP_2829 (  );
sky130_fd_sc_hd__tap_1 TAP_2830 (  );
sky130_fd_sc_hd__tap_1 TAP_2831 (  );
sky130_fd_sc_hd__tap_1 TAP_2832 (  );
sky130_fd_sc_hd__tap_1 TAP_2833 (  );
sky130_fd_sc_hd__tap_1 TAP_2834 (  );
sky130_fd_sc_hd__tap_1 TAP_2835 (  );
sky130_fd_sc_hd__tap_1 TAP_2836 (  );
sky130_fd_sc_hd__tap_1 TAP_2837 (  );
sky130_fd_sc_hd__tap_1 TAP_2838 (  );
sky130_fd_sc_hd__tap_1 TAP_2839 (  );
sky130_fd_sc_hd__tap_1 TAP_2840 (  );
sky130_fd_sc_hd__tap_1 TAP_2841 (  );
sky130_fd_sc_hd__tap_1 TAP_2842 (  );
sky130_fd_sc_hd__tap_1 TAP_2843 (  );
sky130_fd_sc_hd__tap_1 TAP_2844 (  );
sky130_fd_sc_hd__tap_1 TAP_2845 (  );
sky130_fd_sc_hd__tap_1 TAP_2846 (  );
sky130_fd_sc_hd__tap_1 TAP_2847 (  );
sky130_fd_sc_hd__tap_1 TAP_2848 (  );
sky130_fd_sc_hd__tap_1 TAP_2849 (  );
sky130_fd_sc_hd__tap_1 TAP_2850 (  );
sky130_fd_sc_hd__tap_1 TAP_2851 (  );
sky130_fd_sc_hd__tap_1 TAP_2852 (  );
sky130_fd_sc_hd__tap_1 TAP_2853 (  );
sky130_fd_sc_hd__tap_1 TAP_2854 (  );
sky130_fd_sc_hd__tap_1 TAP_2855 (  );
sky130_fd_sc_hd__tap_1 TAP_2856 (  );
sky130_fd_sc_hd__tap_1 TAP_2857 (  );
sky130_fd_sc_hd__tap_1 TAP_2858 (  );
sky130_fd_sc_hd__tap_1 TAP_2859 (  );
sky130_fd_sc_hd__tap_1 TAP_2860 (  );
sky130_fd_sc_hd__tap_1 TAP_2861 (  );
sky130_fd_sc_hd__tap_1 TAP_2862 (  );
sky130_fd_sc_hd__tap_1 TAP_2863 (  );
sky130_fd_sc_hd__tap_1 TAP_2864 (  );
sky130_fd_sc_hd__tap_1 TAP_2865 (  );
sky130_fd_sc_hd__tap_1 TAP_2866 (  );
sky130_fd_sc_hd__tap_1 TAP_2867 (  );
sky130_fd_sc_hd__tap_1 TAP_2868 (  );
sky130_fd_sc_hd__tap_1 TAP_2869 (  );
sky130_fd_sc_hd__tap_1 TAP_2870 (  );
sky130_fd_sc_hd__tap_1 TAP_2871 (  );
sky130_fd_sc_hd__tap_1 TAP_2872 (  );
sky130_fd_sc_hd__tap_1 TAP_2873 (  );
sky130_fd_sc_hd__tap_1 TAP_2874 (  );
sky130_fd_sc_hd__tap_1 TAP_2875 (  );
sky130_fd_sc_hd__tap_1 TAP_2876 (  );
sky130_fd_sc_hd__tap_1 TAP_2877 (  );
sky130_fd_sc_hd__tap_1 TAP_2878 (  );
sky130_fd_sc_hd__tap_1 TAP_2879 (  );
sky130_fd_sc_hd__tap_1 TAP_2880 (  );
sky130_fd_sc_hd__tap_1 TAP_2881 (  );
sky130_fd_sc_hd__tap_1 TAP_2882 (  );
sky130_fd_sc_hd__tap_1 TAP_2883 (  );
sky130_fd_sc_hd__tap_1 TAP_2884 (  );
sky130_fd_sc_hd__tap_1 TAP_2885 (  );
sky130_fd_sc_hd__tap_1 TAP_2886 (  );
sky130_fd_sc_hd__tap_1 TAP_2887 (  );
sky130_fd_sc_hd__tap_1 TAP_2888 (  );
sky130_fd_sc_hd__tap_1 TAP_2889 (  );
sky130_fd_sc_hd__tap_1 TAP_2890 (  );
sky130_fd_sc_hd__tap_1 TAP_2891 (  );
sky130_fd_sc_hd__tap_1 TAP_2892 (  );
sky130_fd_sc_hd__tap_1 TAP_2893 (  );
sky130_fd_sc_hd__tap_1 TAP_2894 (  );
sky130_fd_sc_hd__tap_1 TAP_2895 (  );
sky130_fd_sc_hd__tap_1 TAP_2896 (  );
sky130_fd_sc_hd__tap_1 TAP_2897 (  );
sky130_fd_sc_hd__tap_1 TAP_2898 (  );
sky130_fd_sc_hd__tap_1 TAP_2899 (  );
sky130_fd_sc_hd__tap_1 TAP_2900 (  );
sky130_fd_sc_hd__tap_1 TAP_2901 (  );
sky130_fd_sc_hd__tap_1 TAP_2902 (  );
sky130_fd_sc_hd__tap_1 TAP_2903 (  );
sky130_fd_sc_hd__tap_1 TAP_2904 (  );
sky130_fd_sc_hd__tap_1 TAP_2905 (  );
sky130_fd_sc_hd__tap_1 TAP_2906 (  );
sky130_fd_sc_hd__tap_1 TAP_2907 (  );
sky130_fd_sc_hd__tap_1 TAP_2908 (  );
sky130_fd_sc_hd__tap_1 TAP_2909 (  );
sky130_fd_sc_hd__tap_1 TAP_2910 (  );
sky130_fd_sc_hd__tap_1 TAP_2911 (  );
sky130_fd_sc_hd__tap_1 TAP_2912 (  );
sky130_fd_sc_hd__tap_1 TAP_2913 (  );
sky130_fd_sc_hd__tap_1 TAP_2914 (  );
sky130_fd_sc_hd__tap_1 TAP_2915 (  );
sky130_fd_sc_hd__tap_1 TAP_2916 (  );
sky130_fd_sc_hd__tap_1 TAP_2917 (  );
sky130_fd_sc_hd__tap_1 TAP_2918 (  );
sky130_fd_sc_hd__tap_1 TAP_2919 (  );
sky130_fd_sc_hd__tap_1 TAP_2920 (  );
sky130_fd_sc_hd__tap_1 TAP_2921 (  );
sky130_fd_sc_hd__tap_1 TAP_2922 (  );
sky130_fd_sc_hd__tap_1 TAP_2923 (  );
sky130_fd_sc_hd__tap_1 TAP_2924 (  );
sky130_fd_sc_hd__tap_1 TAP_2925 (  );
sky130_fd_sc_hd__tap_1 TAP_2926 (  );
sky130_fd_sc_hd__tap_1 TAP_2927 (  );
sky130_fd_sc_hd__tap_1 TAP_2928 (  );
sky130_fd_sc_hd__tap_1 TAP_2929 (  );
sky130_fd_sc_hd__tap_1 TAP_2930 (  );
sky130_fd_sc_hd__tap_1 TAP_2931 (  );
sky130_fd_sc_hd__tap_1 TAP_2932 (  );
sky130_fd_sc_hd__tap_1 TAP_2933 (  );
sky130_fd_sc_hd__tap_1 TAP_2934 (  );
sky130_fd_sc_hd__tap_1 TAP_2935 (  );
sky130_fd_sc_hd__tap_1 TAP_2936 (  );
sky130_fd_sc_hd__tap_1 TAP_2937 (  );
sky130_fd_sc_hd__tap_1 TAP_2938 (  );
sky130_fd_sc_hd__tap_1 TAP_2939 (  );
sky130_fd_sc_hd__tap_1 TAP_2940 (  );
sky130_fd_sc_hd__tap_1 TAP_2941 (  );
sky130_fd_sc_hd__tap_1 TAP_2942 (  );
sky130_fd_sc_hd__tap_1 TAP_2943 (  );
sky130_fd_sc_hd__tap_1 TAP_2944 (  );
sky130_fd_sc_hd__tap_1 TAP_2945 (  );
sky130_fd_sc_hd__tap_1 TAP_2946 (  );
sky130_fd_sc_hd__tap_1 TAP_2947 (  );
sky130_fd_sc_hd__tap_1 TAP_2948 (  );
sky130_fd_sc_hd__tap_1 TAP_2949 (  );
sky130_fd_sc_hd__tap_1 TAP_2950 (  );
sky130_fd_sc_hd__tap_1 TAP_2951 (  );
sky130_fd_sc_hd__tap_1 TAP_2952 (  );
sky130_fd_sc_hd__tap_1 TAP_2953 (  );
sky130_fd_sc_hd__tap_1 TAP_2954 (  );
sky130_fd_sc_hd__tap_1 TAP_2955 (  );
sky130_fd_sc_hd__tap_1 TAP_2956 (  );
sky130_fd_sc_hd__tap_1 TAP_2957 (  );
sky130_fd_sc_hd__tap_1 TAP_2958 (  );
sky130_fd_sc_hd__tap_1 TAP_2959 (  );
sky130_fd_sc_hd__tap_1 TAP_2960 (  );
sky130_fd_sc_hd__tap_1 TAP_2961 (  );
sky130_fd_sc_hd__tap_1 TAP_2962 (  );
sky130_fd_sc_hd__tap_1 TAP_2963 (  );
sky130_fd_sc_hd__tap_1 TAP_2964 (  );
sky130_fd_sc_hd__tap_1 TAP_2965 (  );
sky130_fd_sc_hd__tap_1 TAP_2966 (  );
sky130_fd_sc_hd__tap_1 TAP_2967 (  );
sky130_fd_sc_hd__tap_1 TAP_2968 (  );
sky130_fd_sc_hd__tap_1 TAP_2969 (  );
sky130_fd_sc_hd__tap_1 TAP_2970 (  );
sky130_fd_sc_hd__tap_1 TAP_2971 (  );
sky130_fd_sc_hd__tap_1 TAP_2972 (  );
sky130_fd_sc_hd__tap_1 TAP_2973 (  );
sky130_fd_sc_hd__tap_1 TAP_2974 (  );
sky130_fd_sc_hd__tap_1 TAP_2975 (  );
sky130_fd_sc_hd__tap_1 TAP_2976 (  );
sky130_fd_sc_hd__tap_1 TAP_2977 (  );
sky130_fd_sc_hd__tap_1 TAP_2978 (  );
sky130_fd_sc_hd__tap_1 TAP_2979 (  );
sky130_fd_sc_hd__tap_1 TAP_2980 (  );
sky130_fd_sc_hd__tap_1 TAP_2981 (  );
sky130_fd_sc_hd__tap_1 TAP_2982 (  );
sky130_fd_sc_hd__tap_1 TAP_2983 (  );
sky130_fd_sc_hd__tap_1 TAP_2984 (  );
sky130_fd_sc_hd__tap_1 TAP_2985 (  );
sky130_fd_sc_hd__tap_1 TAP_2986 (  );
sky130_fd_sc_hd__tap_1 TAP_2987 (  );
sky130_fd_sc_hd__tap_1 TAP_2988 (  );
sky130_fd_sc_hd__tap_1 TAP_2989 (  );
sky130_fd_sc_hd__tap_1 TAP_2990 (  );
sky130_fd_sc_hd__tap_1 TAP_2991 (  );
sky130_fd_sc_hd__tap_1 TAP_2992 (  );
sky130_fd_sc_hd__tap_1 TAP_2993 (  );
sky130_fd_sc_hd__tap_1 TAP_2994 (  );
sky130_fd_sc_hd__tap_1 TAP_2995 (  );
sky130_fd_sc_hd__tap_1 TAP_2996 (  );
sky130_fd_sc_hd__tap_1 TAP_2997 (  );
sky130_fd_sc_hd__tap_1 TAP_2998 (  );
sky130_fd_sc_hd__tap_1 TAP_2999 (  );
sky130_fd_sc_hd__tap_1 TAP_3000 (  );
sky130_fd_sc_hd__tap_1 TAP_3001 (  );
sky130_fd_sc_hd__tap_1 TAP_3002 (  );
sky130_fd_sc_hd__tap_1 TAP_3003 (  );
sky130_fd_sc_hd__tap_1 TAP_3004 (  );
sky130_fd_sc_hd__tap_1 TAP_3005 (  );
sky130_fd_sc_hd__tap_1 TAP_3006 (  );
sky130_fd_sc_hd__tap_1 TAP_3007 (  );
sky130_fd_sc_hd__tap_1 TAP_3008 (  );
sky130_fd_sc_hd__tap_1 TAP_3009 (  );
sky130_fd_sc_hd__tap_1 TAP_3010 (  );
sky130_fd_sc_hd__tap_1 TAP_3011 (  );
sky130_fd_sc_hd__tap_1 TAP_3012 (  );
sky130_fd_sc_hd__tap_1 TAP_3013 (  );
sky130_fd_sc_hd__tap_1 TAP_3014 (  );
sky130_fd_sc_hd__tap_1 TAP_3015 (  );
sky130_fd_sc_hd__tap_1 TAP_3016 (  );
sky130_fd_sc_hd__tap_1 TAP_3017 (  );
sky130_fd_sc_hd__tap_1 TAP_3018 (  );
sky130_fd_sc_hd__tap_1 TAP_3019 (  );
sky130_fd_sc_hd__tap_1 TAP_3020 (  );
sky130_fd_sc_hd__tap_1 TAP_3021 (  );
sky130_fd_sc_hd__tap_1 TAP_3022 (  );
sky130_fd_sc_hd__tap_1 TAP_3023 (  );
sky130_fd_sc_hd__tap_1 TAP_3024 (  );
sky130_fd_sc_hd__tap_1 TAP_3025 (  );
sky130_fd_sc_hd__tap_1 TAP_3026 (  );
sky130_fd_sc_hd__tap_1 TAP_3027 (  );
sky130_fd_sc_hd__tap_1 TAP_3028 (  );
sky130_fd_sc_hd__tap_1 TAP_3029 (  );
sky130_fd_sc_hd__tap_1 TAP_3030 (  );
sky130_fd_sc_hd__tap_1 TAP_3031 (  );
sky130_fd_sc_hd__tap_1 TAP_3032 (  );
sky130_fd_sc_hd__tap_1 TAP_3033 (  );
sky130_fd_sc_hd__tap_1 TAP_3034 (  );
sky130_fd_sc_hd__tap_1 TAP_3035 (  );
sky130_fd_sc_hd__tap_1 TAP_3036 (  );
sky130_fd_sc_hd__tap_1 TAP_3037 (  );
sky130_fd_sc_hd__tap_1 TAP_3038 (  );
sky130_fd_sc_hd__tap_1 TAP_3039 (  );
sky130_fd_sc_hd__tap_1 TAP_3040 (  );
sky130_fd_sc_hd__tap_1 TAP_3041 (  );
sky130_fd_sc_hd__tap_1 TAP_3042 (  );
sky130_fd_sc_hd__tap_1 TAP_3043 (  );
sky130_fd_sc_hd__tap_1 TAP_3044 (  );
sky130_fd_sc_hd__tap_1 TAP_3045 (  );
sky130_fd_sc_hd__tap_1 TAP_3046 (  );
sky130_fd_sc_hd__tap_1 TAP_3047 (  );
sky130_fd_sc_hd__tap_1 TAP_3048 (  );
sky130_fd_sc_hd__tap_1 TAP_3049 (  );
sky130_fd_sc_hd__tap_1 TAP_3050 (  );
sky130_fd_sc_hd__tap_1 TAP_3051 (  );
sky130_fd_sc_hd__tap_1 TAP_3052 (  );
sky130_fd_sc_hd__tap_1 TAP_3053 (  );
sky130_fd_sc_hd__tap_1 TAP_3054 (  );
sky130_fd_sc_hd__tap_1 TAP_3055 (  );
sky130_fd_sc_hd__tap_1 TAP_3056 (  );
sky130_fd_sc_hd__tap_1 TAP_3057 (  );
sky130_fd_sc_hd__tap_1 TAP_3058 (  );
sky130_fd_sc_hd__tap_1 TAP_3059 (  );
sky130_fd_sc_hd__tap_1 TAP_3060 (  );
sky130_fd_sc_hd__tap_1 TAP_3061 (  );
sky130_fd_sc_hd__tap_1 TAP_3062 (  );
sky130_fd_sc_hd__tap_1 TAP_3063 (  );
sky130_fd_sc_hd__tap_1 TAP_3064 (  );
sky130_fd_sc_hd__tap_1 TAP_3065 (  );
sky130_fd_sc_hd__tap_1 TAP_3066 (  );
sky130_fd_sc_hd__tap_1 TAP_3067 (  );
sky130_fd_sc_hd__tap_1 TAP_3068 (  );
sky130_fd_sc_hd__tap_1 TAP_3069 (  );
sky130_fd_sc_hd__tap_1 TAP_3070 (  );
sky130_fd_sc_hd__tap_1 TAP_3071 (  );
sky130_fd_sc_hd__tap_1 TAP_3072 (  );
sky130_fd_sc_hd__tap_1 TAP_3073 (  );
sky130_fd_sc_hd__tap_1 TAP_3074 (  );
sky130_fd_sc_hd__tap_1 TAP_3075 (  );
sky130_fd_sc_hd__tap_1 TAP_3076 (  );
sky130_fd_sc_hd__tap_1 TAP_3077 (  );
sky130_fd_sc_hd__tap_1 TAP_3078 (  );
sky130_fd_sc_hd__tap_1 TAP_3079 (  );
sky130_fd_sc_hd__tap_1 TAP_3080 (  );
sky130_fd_sc_hd__tap_1 TAP_3081 (  );
sky130_fd_sc_hd__tap_1 TAP_3082 (  );
sky130_fd_sc_hd__tap_1 TAP_3083 (  );
sky130_fd_sc_hd__tap_1 TAP_3084 (  );
sky130_fd_sc_hd__tap_1 TAP_3085 (  );
sky130_fd_sc_hd__tap_1 TAP_3086 (  );
sky130_fd_sc_hd__tap_1 TAP_3087 (  );
sky130_fd_sc_hd__tap_1 TAP_3088 (  );
sky130_fd_sc_hd__tap_1 TAP_3089 (  );
sky130_fd_sc_hd__tap_1 TAP_3090 (  );
sky130_fd_sc_hd__tap_1 TAP_3091 (  );
sky130_fd_sc_hd__tap_1 TAP_3092 (  );
sky130_fd_sc_hd__tap_1 TAP_3093 (  );
sky130_fd_sc_hd__tap_1 TAP_3094 (  );
sky130_fd_sc_hd__tap_1 TAP_3095 (  );
sky130_fd_sc_hd__tap_1 TAP_3096 (  );
sky130_fd_sc_hd__tap_1 TAP_3097 (  );
sky130_fd_sc_hd__tap_1 TAP_3098 (  );
sky130_fd_sc_hd__tap_1 TAP_3099 (  );
sky130_fd_sc_hd__tap_1 TAP_3100 (  );
sky130_fd_sc_hd__tap_1 TAP_3101 (  );
sky130_fd_sc_hd__tap_1 TAP_3102 (  );
sky130_fd_sc_hd__tap_1 TAP_3103 (  );
sky130_fd_sc_hd__tap_1 TAP_3104 (  );
sky130_fd_sc_hd__tap_1 TAP_3105 (  );
sky130_fd_sc_hd__tap_1 TAP_3106 (  );
sky130_fd_sc_hd__tap_1 TAP_3107 (  );
sky130_fd_sc_hd__tap_1 TAP_3108 (  );
sky130_fd_sc_hd__tap_1 TAP_3109 (  );
sky130_fd_sc_hd__tap_1 TAP_3110 (  );
sky130_fd_sc_hd__tap_1 TAP_3111 (  );
sky130_fd_sc_hd__tap_1 TAP_3112 (  );
sky130_fd_sc_hd__tap_1 TAP_3113 (  );
sky130_fd_sc_hd__tap_1 TAP_3114 (  );
sky130_fd_sc_hd__tap_1 TAP_3115 (  );
sky130_fd_sc_hd__tap_1 TAP_3116 (  );
sky130_fd_sc_hd__tap_1 TAP_3117 (  );
sky130_fd_sc_hd__tap_1 TAP_3118 (  );
sky130_fd_sc_hd__tap_1 TAP_3119 (  );
sky130_fd_sc_hd__tap_1 TAP_3120 (  );
sky130_fd_sc_hd__tap_1 TAP_3121 (  );
sky130_fd_sc_hd__tap_1 TAP_3122 (  );
sky130_fd_sc_hd__tap_1 TAP_3123 (  );
sky130_fd_sc_hd__tap_1 TAP_3124 (  );
sky130_fd_sc_hd__tap_1 TAP_3125 (  );
sky130_fd_sc_hd__tap_1 TAP_3126 (  );
sky130_fd_sc_hd__tap_1 TAP_3127 (  );
sky130_fd_sc_hd__tap_1 TAP_3128 (  );
sky130_fd_sc_hd__tap_1 TAP_3129 (  );
sky130_fd_sc_hd__tap_1 TAP_3130 (  );
sky130_fd_sc_hd__tap_1 TAP_3131 (  );
sky130_fd_sc_hd__tap_1 TAP_3132 (  );
sky130_fd_sc_hd__tap_1 TAP_3133 (  );
sky130_fd_sc_hd__tap_1 TAP_3134 (  );
sky130_fd_sc_hd__tap_1 TAP_3135 (  );
sky130_fd_sc_hd__tap_1 TAP_3136 (  );
sky130_fd_sc_hd__tap_1 TAP_3137 (  );
sky130_fd_sc_hd__tap_1 TAP_3138 (  );
sky130_fd_sc_hd__tap_1 TAP_3139 (  );
sky130_fd_sc_hd__tap_1 TAP_3140 (  );
sky130_fd_sc_hd__tap_1 TAP_3141 (  );
sky130_fd_sc_hd__tap_1 TAP_3142 (  );
sky130_fd_sc_hd__tap_1 TAP_3143 (  );
sky130_fd_sc_hd__tap_1 TAP_3144 (  );
sky130_fd_sc_hd__tap_1 TAP_3145 (  );
sky130_fd_sc_hd__tap_1 TAP_3146 (  );
sky130_fd_sc_hd__tap_1 TAP_3147 (  );
sky130_fd_sc_hd__tap_1 TAP_3148 (  );
sky130_fd_sc_hd__tap_1 TAP_3149 (  );
sky130_fd_sc_hd__tap_1 TAP_3150 (  );
sky130_fd_sc_hd__tap_1 TAP_3151 (  );
sky130_fd_sc_hd__tap_1 TAP_3152 (  );
sky130_fd_sc_hd__tap_1 TAP_3153 (  );
sky130_fd_sc_hd__tap_1 TAP_3154 (  );
sky130_fd_sc_hd__tap_1 TAP_3155 (  );
sky130_fd_sc_hd__tap_1 TAP_3156 (  );
sky130_fd_sc_hd__tap_1 TAP_3157 (  );
sky130_fd_sc_hd__tap_1 TAP_3158 (  );
sky130_fd_sc_hd__tap_1 TAP_3159 (  );
sky130_fd_sc_hd__tap_1 TAP_3160 (  );
sky130_fd_sc_hd__tap_1 TAP_3161 (  );
sky130_fd_sc_hd__tap_1 TAP_3162 (  );
sky130_fd_sc_hd__tap_1 TAP_3163 (  );
sky130_fd_sc_hd__tap_1 TAP_3164 (  );
sky130_fd_sc_hd__tap_1 TAP_3165 (  );
sky130_fd_sc_hd__tap_1 TAP_3166 (  );
sky130_fd_sc_hd__tap_1 TAP_3167 (  );
sky130_fd_sc_hd__tap_1 TAP_3168 (  );
sky130_fd_sc_hd__tap_1 TAP_3169 (  );
sky130_fd_sc_hd__tap_1 TAP_3170 (  );
sky130_fd_sc_hd__tap_1 TAP_3171 (  );
sky130_fd_sc_hd__tap_1 TAP_3172 (  );
sky130_fd_sc_hd__tap_1 TAP_3173 (  );
sky130_fd_sc_hd__tap_1 TAP_3174 (  );
sky130_fd_sc_hd__tap_1 TAP_3175 (  );
sky130_fd_sc_hd__tap_1 TAP_3176 (  );
sky130_fd_sc_hd__tap_1 TAP_3177 (  );
sky130_fd_sc_hd__tap_1 TAP_3178 (  );
sky130_fd_sc_hd__tap_1 TAP_3179 (  );
sky130_fd_sc_hd__tap_1 TAP_3180 (  );
sky130_fd_sc_hd__tap_1 TAP_3181 (  );
sky130_fd_sc_hd__tap_1 TAP_3182 (  );
sky130_fd_sc_hd__tap_1 TAP_3183 (  );
sky130_fd_sc_hd__tap_1 TAP_3184 (  );
sky130_fd_sc_hd__tap_1 TAP_3185 (  );
sky130_fd_sc_hd__tap_1 TAP_3186 (  );
sky130_fd_sc_hd__tap_1 TAP_3187 (  );
sky130_fd_sc_hd__tap_1 TAP_3188 (  );
sky130_fd_sc_hd__tap_1 TAP_3189 (  );
sky130_fd_sc_hd__tap_1 TAP_3190 (  );
sky130_fd_sc_hd__tap_1 TAP_3191 (  );
sky130_fd_sc_hd__tap_1 TAP_3192 (  );
sky130_fd_sc_hd__tap_1 TAP_3193 (  );
sky130_fd_sc_hd__tap_1 TAP_3194 (  );
sky130_fd_sc_hd__tap_1 TAP_3195 (  );
sky130_fd_sc_hd__tap_1 TAP_3196 (  );
sky130_fd_sc_hd__tap_1 TAP_3197 (  );
sky130_fd_sc_hd__tap_1 TAP_3198 (  );
sky130_fd_sc_hd__tap_1 TAP_3199 (  );
sky130_fd_sc_hd__tap_1 TAP_3200 (  );
sky130_fd_sc_hd__tap_1 TAP_3201 (  );
sky130_fd_sc_hd__tap_1 TAP_3202 (  );
sky130_fd_sc_hd__tap_1 TAP_3203 (  );
sky130_fd_sc_hd__tap_1 TAP_3204 (  );
sky130_fd_sc_hd__tap_1 TAP_3205 (  );
sky130_fd_sc_hd__tap_1 TAP_3206 (  );
sky130_fd_sc_hd__tap_1 TAP_3207 (  );
sky130_fd_sc_hd__tap_1 TAP_3208 (  );
sky130_fd_sc_hd__tap_1 TAP_3209 (  );
sky130_fd_sc_hd__tap_1 TAP_3210 (  );
sky130_fd_sc_hd__tap_1 TAP_3211 (  );
sky130_fd_sc_hd__tap_1 TAP_3212 (  );
sky130_fd_sc_hd__tap_1 TAP_3213 (  );
sky130_fd_sc_hd__tap_1 TAP_3214 (  );
sky130_fd_sc_hd__tap_1 TAP_3215 (  );
sky130_fd_sc_hd__tap_1 TAP_3216 (  );
sky130_fd_sc_hd__tap_1 TAP_3217 (  );
sky130_fd_sc_hd__tap_1 TAP_3218 (  );
sky130_fd_sc_hd__tap_1 TAP_3219 (  );
sky130_fd_sc_hd__tap_1 TAP_3220 (  );
sky130_fd_sc_hd__tap_1 TAP_3221 (  );
sky130_fd_sc_hd__tap_1 TAP_3222 (  );
sky130_fd_sc_hd__tap_1 TAP_3223 (  );
sky130_fd_sc_hd__tap_1 TAP_3224 (  );
sky130_fd_sc_hd__tap_1 TAP_3225 (  );
sky130_fd_sc_hd__tap_1 TAP_3226 (  );
sky130_fd_sc_hd__tap_1 TAP_3227 (  );
sky130_fd_sc_hd__tap_1 TAP_3228 (  );
sky130_fd_sc_hd__tap_1 TAP_3229 (  );
sky130_fd_sc_hd__tap_1 TAP_3230 (  );
sky130_fd_sc_hd__tap_1 TAP_3231 (  );
sky130_fd_sc_hd__tap_1 TAP_3232 (  );
sky130_fd_sc_hd__tap_1 TAP_3233 (  );
sky130_fd_sc_hd__tap_1 TAP_3234 (  );
sky130_fd_sc_hd__tap_1 TAP_3235 (  );
sky130_fd_sc_hd__tap_1 TAP_3236 (  );
sky130_fd_sc_hd__tap_1 TAP_3237 (  );
sky130_fd_sc_hd__tap_1 TAP_3238 (  );
sky130_fd_sc_hd__tap_1 TAP_3239 (  );
sky130_fd_sc_hd__tap_1 TAP_3240 (  );
sky130_fd_sc_hd__tap_1 TAP_3241 (  );
sky130_fd_sc_hd__tap_1 TAP_3242 (  );
sky130_fd_sc_hd__tap_1 TAP_3243 (  );
sky130_fd_sc_hd__tap_1 TAP_3244 (  );
sky130_fd_sc_hd__tap_1 TAP_3245 (  );
sky130_fd_sc_hd__tap_1 TAP_3246 (  );
sky130_fd_sc_hd__tap_1 TAP_3247 (  );
sky130_fd_sc_hd__tap_1 TAP_3248 (  );
sky130_fd_sc_hd__tap_1 TAP_3249 (  );
sky130_fd_sc_hd__tap_1 TAP_3250 (  );
sky130_fd_sc_hd__tap_1 TAP_3251 (  );
sky130_fd_sc_hd__tap_1 TAP_3252 (  );
sky130_fd_sc_hd__tap_1 TAP_3253 (  );
sky130_fd_sc_hd__tap_1 TAP_3254 (  );
sky130_fd_sc_hd__tap_1 TAP_3255 (  );
sky130_fd_sc_hd__tap_1 TAP_3256 (  );
sky130_fd_sc_hd__tap_1 TAP_3257 (  );
sky130_fd_sc_hd__tap_1 TAP_3258 (  );
sky130_fd_sc_hd__tap_1 TAP_3259 (  );
sky130_fd_sc_hd__tap_1 TAP_3260 (  );
sky130_fd_sc_hd__tap_1 TAP_3261 (  );
sky130_fd_sc_hd__tap_1 TAP_3262 (  );
sky130_fd_sc_hd__tap_1 TAP_3263 (  );
sky130_fd_sc_hd__tap_1 TAP_3264 (  );
sky130_fd_sc_hd__tap_1 TAP_3265 (  );
sky130_fd_sc_hd__tap_1 TAP_3266 (  );
sky130_fd_sc_hd__tap_1 TAP_3267 (  );
sky130_fd_sc_hd__tap_1 TAP_3268 (  );
sky130_fd_sc_hd__tap_1 TAP_3269 (  );
sky130_fd_sc_hd__tap_1 TAP_3270 (  );
sky130_fd_sc_hd__tap_1 TAP_3271 (  );
sky130_fd_sc_hd__tap_1 TAP_3272 (  );
sky130_fd_sc_hd__tap_1 TAP_3273 (  );
sky130_fd_sc_hd__tap_1 TAP_3274 (  );
sky130_fd_sc_hd__tap_1 TAP_3275 (  );
sky130_fd_sc_hd__tap_1 TAP_3276 (  );
sky130_fd_sc_hd__tap_1 TAP_3277 (  );
sky130_fd_sc_hd__tap_1 TAP_3278 (  );
sky130_fd_sc_hd__tap_1 TAP_3279 (  );
sky130_fd_sc_hd__tap_1 TAP_3280 (  );
sky130_fd_sc_hd__tap_1 TAP_3281 (  );
sky130_fd_sc_hd__tap_1 TAP_3282 (  );
sky130_fd_sc_hd__tap_1 TAP_3283 (  );
sky130_fd_sc_hd__tap_1 TAP_3284 (  );
sky130_fd_sc_hd__tap_1 TAP_3285 (  );
sky130_fd_sc_hd__tap_1 TAP_3286 (  );
sky130_fd_sc_hd__tap_1 TAP_3287 (  );
sky130_fd_sc_hd__tap_1 TAP_3288 (  );
sky130_fd_sc_hd__tap_1 TAP_3289 (  );
sky130_fd_sc_hd__tap_1 TAP_3290 (  );
sky130_fd_sc_hd__tap_1 TAP_3291 (  );
sky130_fd_sc_hd__tap_1 TAP_3292 (  );
sky130_fd_sc_hd__tap_1 TAP_3293 (  );
sky130_fd_sc_hd__tap_1 TAP_3294 (  );
sky130_fd_sc_hd__tap_1 TAP_3295 (  );
sky130_fd_sc_hd__tap_1 TAP_3296 (  );
sky130_fd_sc_hd__tap_1 TAP_3297 (  );
sky130_fd_sc_hd__tap_1 TAP_3298 (  );
sky130_fd_sc_hd__tap_1 TAP_3299 (  );
sky130_fd_sc_hd__tap_1 TAP_3300 (  );
sky130_fd_sc_hd__tap_1 TAP_3301 (  );
sky130_fd_sc_hd__tap_1 TAP_3302 (  );
sky130_fd_sc_hd__tap_1 TAP_3303 (  );
sky130_fd_sc_hd__tap_1 TAP_3304 (  );
sky130_fd_sc_hd__tap_1 TAP_3305 (  );
sky130_fd_sc_hd__tap_1 TAP_3306 (  );
sky130_fd_sc_hd__tap_1 TAP_3307 (  );
sky130_fd_sc_hd__tap_1 TAP_3308 (  );
sky130_fd_sc_hd__tap_1 TAP_3309 (  );
sky130_fd_sc_hd__tap_1 TAP_3310 (  );
sky130_fd_sc_hd__tap_1 TAP_3311 (  );
sky130_fd_sc_hd__tap_1 TAP_3312 (  );
sky130_fd_sc_hd__tap_1 TAP_3313 (  );
sky130_fd_sc_hd__tap_1 TAP_3314 (  );
sky130_fd_sc_hd__tap_1 TAP_3315 (  );
sky130_fd_sc_hd__tap_1 TAP_3316 (  );
sky130_fd_sc_hd__tap_1 TAP_3317 (  );
sky130_fd_sc_hd__tap_1 TAP_3318 (  );
sky130_fd_sc_hd__tap_1 TAP_3319 (  );
sky130_fd_sc_hd__tap_1 TAP_3320 (  );
sky130_fd_sc_hd__tap_1 TAP_3321 (  );
sky130_fd_sc_hd__tap_1 TAP_3322 (  );
sky130_fd_sc_hd__tap_1 TAP_3323 (  );
sky130_fd_sc_hd__tap_1 TAP_3324 (  );
sky130_fd_sc_hd__tap_1 TAP_3325 (  );
sky130_fd_sc_hd__tap_1 TAP_3326 (  );
sky130_fd_sc_hd__tap_1 TAP_3327 (  );
sky130_fd_sc_hd__tap_1 TAP_3328 (  );
sky130_fd_sc_hd__tap_1 TAP_3329 (  );
sky130_fd_sc_hd__tap_1 TAP_3330 (  );
sky130_fd_sc_hd__tap_1 TAP_3331 (  );
sky130_fd_sc_hd__tap_1 TAP_3332 (  );
sky130_fd_sc_hd__tap_1 TAP_3333 (  );
sky130_fd_sc_hd__tap_1 TAP_3334 (  );
sky130_fd_sc_hd__tap_1 TAP_3335 (  );
sky130_fd_sc_hd__tap_1 TAP_3336 (  );
sky130_fd_sc_hd__tap_1 TAP_3337 (  );
sky130_fd_sc_hd__tap_1 TAP_3338 (  );
sky130_fd_sc_hd__tap_1 TAP_3339 (  );
sky130_fd_sc_hd__tap_1 TAP_3340 (  );
sky130_fd_sc_hd__tap_1 TAP_3341 (  );
sky130_fd_sc_hd__tap_1 TAP_3342 (  );
sky130_fd_sc_hd__tap_1 TAP_3343 (  );
sky130_fd_sc_hd__tap_1 TAP_3344 (  );
sky130_fd_sc_hd__tap_1 TAP_3345 (  );
sky130_fd_sc_hd__tap_1 TAP_3346 (  );
sky130_fd_sc_hd__tap_1 TAP_3347 (  );
sky130_fd_sc_hd__tap_1 TAP_3348 (  );
sky130_fd_sc_hd__tap_1 TAP_3349 (  );
sky130_fd_sc_hd__tap_1 TAP_3350 (  );
sky130_fd_sc_hd__tap_1 TAP_3351 (  );
sky130_fd_sc_hd__tap_1 TAP_3352 (  );
sky130_fd_sc_hd__tap_1 TAP_3353 (  );
sky130_fd_sc_hd__tap_1 TAP_3354 (  );
sky130_fd_sc_hd__tap_1 TAP_3355 (  );
sky130_fd_sc_hd__tap_1 TAP_3356 (  );
sky130_fd_sc_hd__tap_1 TAP_3357 (  );
sky130_fd_sc_hd__tap_1 TAP_3358 (  );
sky130_fd_sc_hd__tap_1 TAP_3359 (  );
sky130_fd_sc_hd__tap_1 TAP_3360 (  );
sky130_fd_sc_hd__tap_1 TAP_3361 (  );
sky130_fd_sc_hd__tap_1 TAP_3362 (  );
sky130_fd_sc_hd__tap_1 TAP_3363 (  );
sky130_fd_sc_hd__tap_1 TAP_3364 (  );
sky130_fd_sc_hd__tap_1 TAP_3365 (  );
sky130_fd_sc_hd__tap_1 TAP_3366 (  );
sky130_fd_sc_hd__tap_1 TAP_3367 (  );
sky130_fd_sc_hd__tap_1 TAP_3368 (  );
sky130_fd_sc_hd__tap_1 TAP_3369 (  );
sky130_fd_sc_hd__tap_1 TAP_3370 (  );
sky130_fd_sc_hd__tap_1 TAP_3371 (  );
sky130_fd_sc_hd__tap_1 TAP_3372 (  );
sky130_fd_sc_hd__tap_1 TAP_3373 (  );
sky130_fd_sc_hd__tap_1 TAP_3374 (  );
sky130_fd_sc_hd__tap_1 TAP_3375 (  );
sky130_fd_sc_hd__tap_1 TAP_3376 (  );
sky130_fd_sc_hd__tap_1 TAP_3377 (  );
sky130_fd_sc_hd__tap_1 TAP_3378 (  );
sky130_fd_sc_hd__tap_1 TAP_3379 (  );
sky130_fd_sc_hd__tap_1 TAP_3380 (  );
sky130_fd_sc_hd__tap_1 TAP_3381 (  );
sky130_fd_sc_hd__tap_1 TAP_3382 (  );
sky130_fd_sc_hd__tap_1 TAP_3383 (  );
sky130_fd_sc_hd__tap_1 TAP_3384 (  );
sky130_fd_sc_hd__tap_1 TAP_3385 (  );
sky130_fd_sc_hd__tap_1 TAP_3386 (  );
sky130_fd_sc_hd__tap_1 TAP_3387 (  );
sky130_fd_sc_hd__tap_1 TAP_3388 (  );
sky130_fd_sc_hd__tap_1 TAP_3389 (  );
sky130_fd_sc_hd__tap_1 TAP_3390 (  );
sky130_fd_sc_hd__tap_1 TAP_3391 (  );
sky130_fd_sc_hd__tap_1 TAP_3392 (  );
sky130_fd_sc_hd__tap_1 TAP_3393 (  );
sky130_fd_sc_hd__tap_1 TAP_3394 (  );
sky130_fd_sc_hd__tap_1 TAP_3395 (  );
sky130_fd_sc_hd__tap_1 TAP_3396 (  );
sky130_fd_sc_hd__tap_1 TAP_3397 (  );
sky130_fd_sc_hd__tap_1 TAP_3398 (  );
sky130_fd_sc_hd__tap_1 TAP_3399 (  );
sky130_fd_sc_hd__tap_1 TAP_3400 (  );
sky130_fd_sc_hd__tap_1 TAP_3401 (  );
sky130_fd_sc_hd__tap_1 TAP_3402 (  );
sky130_fd_sc_hd__tap_1 TAP_3403 (  );
sky130_fd_sc_hd__tap_1 TAP_3404 (  );
sky130_fd_sc_hd__tap_1 TAP_3405 (  );
sky130_fd_sc_hd__tap_1 TAP_3406 (  );
sky130_fd_sc_hd__tap_1 TAP_3407 (  );
sky130_fd_sc_hd__tap_1 TAP_3408 (  );
sky130_fd_sc_hd__tap_1 TAP_3409 (  );
sky130_fd_sc_hd__tap_1 TAP_3410 (  );
sky130_fd_sc_hd__tap_1 TAP_3411 (  );
sky130_fd_sc_hd__tap_1 TAP_3412 (  );
sky130_fd_sc_hd__tap_1 TAP_3413 (  );
sky130_fd_sc_hd__tap_1 TAP_3414 (  );
sky130_fd_sc_hd__tap_1 TAP_3415 (  );
sky130_fd_sc_hd__tap_1 TAP_3416 (  );
sky130_fd_sc_hd__tap_1 TAP_3417 (  );
sky130_fd_sc_hd__tap_1 TAP_3418 (  );
sky130_fd_sc_hd__tap_1 TAP_3419 (  );
sky130_fd_sc_hd__tap_1 TAP_3420 (  );
sky130_fd_sc_hd__tap_1 TAP_3421 (  );
sky130_fd_sc_hd__tap_1 TAP_3422 (  );
sky130_fd_sc_hd__tap_1 TAP_3423 (  );
sky130_fd_sc_hd__tap_1 TAP_3424 (  );
sky130_fd_sc_hd__tap_1 TAP_3425 (  );
sky130_fd_sc_hd__tap_1 TAP_3426 (  );
sky130_fd_sc_hd__tap_1 TAP_3427 (  );
sky130_fd_sc_hd__tap_1 TAP_3428 (  );
sky130_fd_sc_hd__tap_1 TAP_3429 (  );
sky130_fd_sc_hd__tap_1 TAP_3430 (  );
sky130_fd_sc_hd__tap_1 TAP_3431 (  );
sky130_fd_sc_hd__tap_1 TAP_3432 (  );
sky130_fd_sc_hd__tap_1 TAP_3433 (  );
sky130_fd_sc_hd__tap_1 TAP_3434 (  );
sky130_fd_sc_hd__tap_1 TAP_3435 (  );
sky130_fd_sc_hd__tap_1 TAP_3436 (  );
sky130_fd_sc_hd__tap_1 TAP_3437 (  );
sky130_fd_sc_hd__tap_1 TAP_3438 (  );
sky130_fd_sc_hd__tap_1 TAP_3439 (  );
sky130_fd_sc_hd__tap_1 TAP_3440 (  );
sky130_fd_sc_hd__tap_1 TAP_3441 (  );
sky130_fd_sc_hd__tap_1 TAP_3442 (  );
sky130_fd_sc_hd__tap_1 TAP_3443 (  );
sky130_fd_sc_hd__tap_1 TAP_3444 (  );
sky130_fd_sc_hd__tap_1 TAP_3445 (  );
sky130_fd_sc_hd__tap_1 TAP_3446 (  );
sky130_fd_sc_hd__tap_1 TAP_3447 (  );
sky130_fd_sc_hd__tap_1 TAP_3448 (  );
sky130_fd_sc_hd__tap_1 TAP_3449 (  );
sky130_fd_sc_hd__tap_1 TAP_3450 (  );
sky130_fd_sc_hd__tap_1 TAP_3451 (  );
sky130_fd_sc_hd__tap_1 TAP_3452 (  );
sky130_fd_sc_hd__tap_1 TAP_3453 (  );
sky130_fd_sc_hd__tap_1 TAP_3454 (  );
sky130_fd_sc_hd__tap_1 TAP_3455 (  );
sky130_fd_sc_hd__tap_1 TAP_3456 (  );
sky130_fd_sc_hd__tap_1 TAP_3457 (  );
sky130_fd_sc_hd__tap_1 TAP_3458 (  );
sky130_fd_sc_hd__tap_1 TAP_3459 (  );
sky130_fd_sc_hd__tap_1 TAP_3460 (  );
sky130_fd_sc_hd__tap_1 TAP_3461 (  );
sky130_fd_sc_hd__tap_1 TAP_3462 (  );
sky130_fd_sc_hd__tap_1 TAP_3463 (  );
sky130_fd_sc_hd__tap_1 TAP_3464 (  );
sky130_fd_sc_hd__tap_1 TAP_3465 (  );
sky130_fd_sc_hd__tap_1 TAP_3466 (  );
sky130_fd_sc_hd__tap_1 TAP_3467 (  );
sky130_fd_sc_hd__tap_1 TAP_3468 (  );
sky130_fd_sc_hd__tap_1 TAP_3469 (  );
sky130_fd_sc_hd__tap_1 TAP_3470 (  );
sky130_fd_sc_hd__tap_1 TAP_3471 (  );
sky130_fd_sc_hd__tap_1 TAP_3472 (  );
sky130_fd_sc_hd__tap_1 TAP_3473 (  );
sky130_fd_sc_hd__tap_1 TAP_3474 (  );
sky130_fd_sc_hd__tap_1 TAP_3475 (  );
sky130_fd_sc_hd__tap_1 TAP_3476 (  );
sky130_fd_sc_hd__tap_1 TAP_3477 (  );
sky130_fd_sc_hd__tap_1 TAP_3478 (  );
sky130_fd_sc_hd__tap_1 TAP_3479 (  );
sky130_fd_sc_hd__tap_1 TAP_3480 (  );
sky130_fd_sc_hd__tap_1 TAP_3481 (  );
sky130_fd_sc_hd__tap_1 TAP_3482 (  );
sky130_fd_sc_hd__tap_1 TAP_3483 (  );
sky130_fd_sc_hd__tap_1 TAP_3484 (  );
sky130_fd_sc_hd__tap_1 TAP_3485 (  );
sky130_fd_sc_hd__tap_1 TAP_3486 (  );
sky130_fd_sc_hd__tap_1 TAP_3487 (  );
sky130_fd_sc_hd__tap_1 TAP_3488 (  );
sky130_fd_sc_hd__tap_1 TAP_3489 (  );
sky130_fd_sc_hd__tap_1 TAP_3490 (  );
sky130_fd_sc_hd__tap_1 TAP_3491 (  );
sky130_fd_sc_hd__tap_1 TAP_3492 (  );
sky130_fd_sc_hd__tap_1 TAP_3493 (  );
sky130_fd_sc_hd__tap_1 TAP_3494 (  );
sky130_fd_sc_hd__tap_1 TAP_3495 (  );
sky130_fd_sc_hd__tap_1 TAP_3496 (  );
sky130_fd_sc_hd__tap_1 TAP_3497 (  );
sky130_fd_sc_hd__tap_1 TAP_3498 (  );
sky130_fd_sc_hd__tap_1 TAP_3499 (  );
sky130_fd_sc_hd__tap_1 TAP_3500 (  );
sky130_fd_sc_hd__tap_1 TAP_3501 (  );
sky130_fd_sc_hd__tap_1 TAP_3502 (  );
sky130_fd_sc_hd__tap_1 TAP_3503 (  );
sky130_fd_sc_hd__tap_1 TAP_3504 (  );
sky130_fd_sc_hd__tap_1 TAP_3505 (  );
sky130_fd_sc_hd__tap_1 TAP_3506 (  );
sky130_fd_sc_hd__tap_1 TAP_3507 (  );
sky130_fd_sc_hd__tap_1 TAP_3508 (  );
sky130_fd_sc_hd__tap_1 TAP_3509 (  );
sky130_fd_sc_hd__tap_1 TAP_3510 (  );
sky130_fd_sc_hd__tap_1 TAP_3511 (  );
sky130_fd_sc_hd__tap_1 TAP_3512 (  );
sky130_fd_sc_hd__tap_1 TAP_3513 (  );
sky130_fd_sc_hd__tap_1 TAP_3514 (  );
sky130_fd_sc_hd__tap_1 TAP_3515 (  );
sky130_fd_sc_hd__tap_1 TAP_3516 (  );
sky130_fd_sc_hd__tap_1 TAP_3517 (  );
sky130_fd_sc_hd__tap_1 TAP_3518 (  );
sky130_fd_sc_hd__tap_1 TAP_3519 (  );
sky130_fd_sc_hd__tap_1 TAP_3520 (  );
sky130_fd_sc_hd__tap_1 TAP_3521 (  );
sky130_fd_sc_hd__tap_1 TAP_3522 (  );
sky130_fd_sc_hd__tap_1 TAP_3523 (  );
sky130_fd_sc_hd__tap_1 TAP_3524 (  );
sky130_fd_sc_hd__tap_1 TAP_3525 (  );
sky130_fd_sc_hd__tap_1 TAP_3526 (  );
sky130_fd_sc_hd__tap_1 TAP_3527 (  );
sky130_fd_sc_hd__tap_1 TAP_3528 (  );
sky130_fd_sc_hd__tap_1 TAP_3529 (  );
sky130_fd_sc_hd__tap_1 TAP_3530 (  );
sky130_fd_sc_hd__tap_1 TAP_3531 (  );
sky130_fd_sc_hd__tap_1 TAP_3532 (  );
sky130_fd_sc_hd__tap_1 TAP_3533 (  );
sky130_fd_sc_hd__tap_1 TAP_3534 (  );
sky130_fd_sc_hd__tap_1 TAP_3535 (  );
sky130_fd_sc_hd__tap_1 TAP_3536 (  );
sky130_fd_sc_hd__tap_1 TAP_3537 (  );
sky130_fd_sc_hd__tap_1 TAP_3538 (  );
sky130_fd_sc_hd__tap_1 TAP_3539 (  );
sky130_fd_sc_hd__tap_1 TAP_3540 (  );
sky130_fd_sc_hd__tap_1 TAP_3541 (  );
sky130_fd_sc_hd__tap_1 TAP_3542 (  );
sky130_fd_sc_hd__tap_1 TAP_3543 (  );
sky130_fd_sc_hd__tap_1 TAP_3544 (  );
sky130_fd_sc_hd__tap_1 TAP_3545 (  );
sky130_fd_sc_hd__tap_1 TAP_3546 (  );
sky130_fd_sc_hd__tap_1 TAP_3547 (  );
sky130_fd_sc_hd__tap_1 TAP_3548 (  );
sky130_fd_sc_hd__tap_1 TAP_3549 (  );
sky130_fd_sc_hd__tap_1 TAP_3550 (  );
sky130_fd_sc_hd__tap_1 TAP_3551 (  );
sky130_fd_sc_hd__tap_1 TAP_3552 (  );
sky130_fd_sc_hd__tap_1 TAP_3553 (  );
sky130_fd_sc_hd__tap_1 TAP_3554 (  );
sky130_fd_sc_hd__tap_1 TAP_3555 (  );
sky130_fd_sc_hd__tap_1 TAP_3556 (  );
sky130_fd_sc_hd__tap_1 TAP_3557 (  );
sky130_fd_sc_hd__tap_1 TAP_3558 (  );
sky130_fd_sc_hd__tap_1 TAP_3559 (  );
sky130_fd_sc_hd__tap_1 TAP_3560 (  );
sky130_fd_sc_hd__tap_1 TAP_3561 (  );
sky130_fd_sc_hd__tap_1 TAP_3562 (  );
sky130_fd_sc_hd__tap_1 TAP_3563 (  );
sky130_fd_sc_hd__tap_1 TAP_3564 (  );
sky130_fd_sc_hd__tap_1 TAP_3565 (  );
sky130_fd_sc_hd__tap_1 TAP_3566 (  );
sky130_fd_sc_hd__tap_1 TAP_3567 (  );
sky130_fd_sc_hd__tap_1 TAP_3568 (  );
sky130_fd_sc_hd__tap_1 TAP_3569 (  );
sky130_fd_sc_hd__tap_1 TAP_3570 (  );
sky130_fd_sc_hd__tap_1 TAP_3571 (  );
sky130_fd_sc_hd__tap_1 TAP_3572 (  );
sky130_fd_sc_hd__tap_1 TAP_3573 (  );
sky130_fd_sc_hd__tap_1 TAP_3574 (  );
sky130_fd_sc_hd__tap_1 TAP_3575 (  );
sky130_fd_sc_hd__tap_1 TAP_3576 (  );
sky130_fd_sc_hd__tap_1 TAP_3577 (  );
sky130_fd_sc_hd__tap_1 TAP_3578 (  );
sky130_fd_sc_hd__tap_1 TAP_3579 (  );
sky130_fd_sc_hd__tap_1 TAP_3580 (  );
sky130_fd_sc_hd__tap_1 TAP_3581 (  );
sky130_fd_sc_hd__tap_1 TAP_3582 (  );
sky130_fd_sc_hd__tap_1 TAP_3583 (  );
sky130_fd_sc_hd__tap_1 TAP_3584 (  );
sky130_fd_sc_hd__tap_1 TAP_3585 (  );
sky130_fd_sc_hd__tap_1 TAP_3586 (  );
sky130_fd_sc_hd__tap_1 TAP_3587 (  );
sky130_fd_sc_hd__tap_1 TAP_3588 (  );
sky130_fd_sc_hd__tap_1 TAP_3589 (  );
sky130_fd_sc_hd__tap_1 TAP_3590 (  );
sky130_fd_sc_hd__tap_1 TAP_3591 (  );
sky130_fd_sc_hd__tap_1 TAP_3592 (  );
sky130_fd_sc_hd__tap_1 TAP_3593 (  );
sky130_fd_sc_hd__tap_1 TAP_3594 (  );
sky130_fd_sc_hd__tap_1 TAP_3595 (  );
sky130_fd_sc_hd__tap_1 TAP_3596 (  );
sky130_fd_sc_hd__tap_1 TAP_3597 (  );
sky130_fd_sc_hd__tap_1 TAP_3598 (  );
sky130_fd_sc_hd__tap_1 TAP_3599 (  );
sky130_fd_sc_hd__tap_1 TAP_3600 (  );
sky130_fd_sc_hd__tap_1 TAP_3601 (  );
sky130_fd_sc_hd__tap_1 TAP_3602 (  );
sky130_fd_sc_hd__tap_1 TAP_3603 (  );
sky130_fd_sc_hd__tap_1 TAP_3604 (  );
sky130_fd_sc_hd__tap_1 TAP_3605 (  );
sky130_fd_sc_hd__tap_1 TAP_3606 (  );
sky130_fd_sc_hd__tap_1 TAP_3607 (  );
sky130_fd_sc_hd__tap_1 TAP_3608 (  );
sky130_fd_sc_hd__tap_1 TAP_3609 (  );
sky130_fd_sc_hd__tap_1 TAP_3610 (  );
sky130_fd_sc_hd__tap_1 TAP_3611 (  );
sky130_fd_sc_hd__tap_1 TAP_3612 (  );
sky130_fd_sc_hd__tap_1 TAP_3613 (  );
sky130_fd_sc_hd__tap_1 TAP_3614 (  );
sky130_fd_sc_hd__tap_1 TAP_3615 (  );
sky130_fd_sc_hd__tap_1 TAP_3616 (  );
sky130_fd_sc_hd__tap_1 TAP_3617 (  );
sky130_fd_sc_hd__tap_1 TAP_3618 (  );
sky130_fd_sc_hd__tap_1 TAP_3619 (  );
sky130_fd_sc_hd__tap_1 TAP_3620 (  );
sky130_fd_sc_hd__tap_1 TAP_3621 (  );
sky130_fd_sc_hd__tap_1 TAP_3622 (  );
sky130_fd_sc_hd__tap_1 TAP_3623 (  );
sky130_fd_sc_hd__tap_1 TAP_3624 (  );
sky130_fd_sc_hd__tap_1 TAP_3625 (  );
sky130_fd_sc_hd__tap_1 TAP_3626 (  );
sky130_fd_sc_hd__tap_1 TAP_3627 (  );
sky130_fd_sc_hd__tap_1 TAP_3628 (  );
sky130_fd_sc_hd__tap_1 TAP_3629 (  );
sky130_fd_sc_hd__tap_1 TAP_3630 (  );
sky130_fd_sc_hd__tap_1 TAP_3631 (  );
sky130_fd_sc_hd__tap_1 TAP_3632 (  );
sky130_fd_sc_hd__tap_1 TAP_3633 (  );
sky130_fd_sc_hd__tap_1 TAP_3634 (  );
sky130_fd_sc_hd__tap_1 TAP_3635 (  );
sky130_fd_sc_hd__tap_1 TAP_3636 (  );
sky130_fd_sc_hd__tap_1 TAP_3637 (  );
sky130_fd_sc_hd__tap_1 TAP_3638 (  );
sky130_fd_sc_hd__tap_1 TAP_3639 (  );
sky130_fd_sc_hd__tap_1 TAP_3640 (  );
sky130_fd_sc_hd__tap_1 TAP_3641 (  );
sky130_fd_sc_hd__tap_1 TAP_3642 (  );
sky130_fd_sc_hd__tap_1 TAP_3643 (  );
sky130_fd_sc_hd__tap_1 TAP_3644 (  );
sky130_fd_sc_hd__tap_1 TAP_3645 (  );
sky130_fd_sc_hd__tap_1 TAP_3646 (  );
sky130_fd_sc_hd__tap_1 TAP_3647 (  );
sky130_fd_sc_hd__tap_1 TAP_3648 (  );
sky130_fd_sc_hd__tap_1 TAP_3649 (  );
sky130_fd_sc_hd__tap_1 TAP_3650 (  );
sky130_fd_sc_hd__tap_1 TAP_3651 (  );
sky130_fd_sc_hd__tap_1 TAP_3652 (  );
sky130_fd_sc_hd__tap_1 TAP_3653 (  );
sky130_fd_sc_hd__tap_1 TAP_3654 (  );
sky130_fd_sc_hd__tap_1 TAP_3655 (  );
sky130_fd_sc_hd__tap_1 TAP_3656 (  );
sky130_fd_sc_hd__tap_1 TAP_3657 (  );
sky130_fd_sc_hd__tap_1 TAP_3658 (  );
sky130_fd_sc_hd__tap_1 TAP_3659 (  );
sky130_fd_sc_hd__tap_1 TAP_3660 (  );
sky130_fd_sc_hd__tap_1 TAP_3661 (  );
sky130_fd_sc_hd__tap_1 TAP_3662 (  );
sky130_fd_sc_hd__tap_1 TAP_3663 (  );
sky130_fd_sc_hd__tap_1 TAP_3664 (  );
sky130_fd_sc_hd__tap_1 TAP_3665 (  );
sky130_fd_sc_hd__tap_1 TAP_3666 (  );
sky130_fd_sc_hd__tap_1 TAP_3667 (  );
sky130_fd_sc_hd__tap_1 TAP_3668 (  );
sky130_fd_sc_hd__tap_1 TAP_3669 (  );
sky130_fd_sc_hd__tap_1 TAP_3670 (  );
sky130_fd_sc_hd__tap_1 TAP_3671 (  );
sky130_fd_sc_hd__tap_1 TAP_3672 (  );
sky130_fd_sc_hd__tap_1 TAP_3673 (  );
sky130_fd_sc_hd__tap_1 TAP_3674 (  );
sky130_fd_sc_hd__tap_1 TAP_3675 (  );
sky130_fd_sc_hd__tap_1 TAP_3676 (  );
sky130_fd_sc_hd__tap_1 TAP_3677 (  );
sky130_fd_sc_hd__tap_1 TAP_3678 (  );
sky130_fd_sc_hd__tap_1 TAP_3679 (  );
sky130_fd_sc_hd__tap_1 TAP_3680 (  );
sky130_fd_sc_hd__tap_1 TAP_3681 (  );
sky130_fd_sc_hd__tap_1 TAP_3682 (  );
sky130_fd_sc_hd__tap_1 TAP_3683 (  );
sky130_fd_sc_hd__tap_1 TAP_3684 (  );
sky130_fd_sc_hd__tap_1 TAP_3685 (  );
sky130_fd_sc_hd__tap_1 TAP_3686 (  );
sky130_fd_sc_hd__tap_1 TAP_3687 (  );
sky130_fd_sc_hd__tap_1 TAP_3688 (  );
sky130_fd_sc_hd__tap_1 TAP_3689 (  );
sky130_fd_sc_hd__tap_1 TAP_3690 (  );
sky130_fd_sc_hd__tap_1 TAP_3691 (  );
sky130_fd_sc_hd__tap_1 TAP_3692 (  );
sky130_fd_sc_hd__tap_1 TAP_3693 (  );
sky130_fd_sc_hd__tap_1 TAP_3694 (  );
sky130_fd_sc_hd__tap_1 TAP_3695 (  );
sky130_fd_sc_hd__tap_1 TAP_3696 (  );
sky130_fd_sc_hd__tap_1 TAP_3697 (  );
sky130_fd_sc_hd__tap_1 TAP_3698 (  );
sky130_fd_sc_hd__tap_1 TAP_3699 (  );
sky130_fd_sc_hd__tap_1 TAP_3700 (  );
sky130_fd_sc_hd__tap_1 TAP_3701 (  );
sky130_fd_sc_hd__tap_1 TAP_3702 (  );
sky130_fd_sc_hd__tap_1 TAP_3703 (  );
sky130_fd_sc_hd__tap_1 TAP_3704 (  );
sky130_fd_sc_hd__tap_1 TAP_3705 (  );
sky130_fd_sc_hd__tap_1 TAP_3706 (  );
sky130_fd_sc_hd__tap_1 TAP_3707 (  );
sky130_fd_sc_hd__tap_1 TAP_3708 (  );
sky130_fd_sc_hd__tap_1 TAP_3709 (  );
sky130_fd_sc_hd__tap_1 TAP_3710 (  );
sky130_fd_sc_hd__tap_1 TAP_3711 (  );
sky130_fd_sc_hd__tap_1 TAP_3712 (  );
sky130_fd_sc_hd__tap_1 TAP_3713 (  );
sky130_fd_sc_hd__tap_1 TAP_3714 (  );
sky130_fd_sc_hd__tap_1 TAP_3715 (  );
sky130_fd_sc_hd__tap_1 TAP_3716 (  );
sky130_fd_sc_hd__tap_1 TAP_3717 (  );
sky130_fd_sc_hd__tap_1 TAP_3718 (  );
sky130_fd_sc_hd__tap_1 TAP_3719 (  );
sky130_fd_sc_hd__tap_1 TAP_3720 (  );
sky130_fd_sc_hd__tap_1 TAP_3721 (  );
sky130_fd_sc_hd__tap_1 TAP_3722 (  );
sky130_fd_sc_hd__tap_1 TAP_3723 (  );
sky130_fd_sc_hd__tap_1 TAP_3724 (  );
sky130_fd_sc_hd__tap_1 TAP_3725 (  );
sky130_fd_sc_hd__tap_1 TAP_3726 (  );
sky130_fd_sc_hd__tap_1 TAP_3727 (  );
sky130_fd_sc_hd__tap_1 TAP_3728 (  );
sky130_fd_sc_hd__tap_1 TAP_3729 (  );
sky130_fd_sc_hd__tap_1 TAP_3730 (  );
sky130_fd_sc_hd__tap_1 TAP_3731 (  );
sky130_fd_sc_hd__tap_1 TAP_3732 (  );
sky130_fd_sc_hd__tap_1 TAP_3733 (  );
sky130_fd_sc_hd__tap_1 TAP_3734 (  );
sky130_fd_sc_hd__tap_1 TAP_3735 (  );
sky130_fd_sc_hd__tap_1 TAP_3736 (  );
sky130_fd_sc_hd__tap_1 TAP_3737 (  );
sky130_fd_sc_hd__tap_1 TAP_3738 (  );
sky130_fd_sc_hd__tap_1 TAP_3739 (  );
sky130_fd_sc_hd__tap_1 TAP_3740 (  );
sky130_fd_sc_hd__tap_1 TAP_3741 (  );
sky130_fd_sc_hd__tap_1 TAP_3742 (  );
sky130_fd_sc_hd__tap_1 TAP_3743 (  );
sky130_fd_sc_hd__tap_1 TAP_3744 (  );
sky130_fd_sc_hd__tap_1 TAP_3745 (  );
sky130_fd_sc_hd__tap_1 TAP_3746 (  );
sky130_fd_sc_hd__tap_1 TAP_3747 (  );
sky130_fd_sc_hd__tap_1 TAP_3748 (  );
sky130_fd_sc_hd__tap_1 TAP_3749 (  );
sky130_fd_sc_hd__tap_1 TAP_3750 (  );
sky130_fd_sc_hd__tap_1 TAP_3751 (  );
sky130_fd_sc_hd__tap_1 TAP_3752 (  );
sky130_fd_sc_hd__tap_1 TAP_3753 (  );
sky130_fd_sc_hd__tap_1 TAP_3754 (  );
sky130_fd_sc_hd__tap_1 TAP_3755 (  );
sky130_fd_sc_hd__tap_1 TAP_3756 (  );
sky130_fd_sc_hd__tap_1 TAP_3757 (  );
sky130_fd_sc_hd__tap_1 TAP_3758 (  );
sky130_fd_sc_hd__tap_1 TAP_3759 (  );
sky130_fd_sc_hd__tap_1 TAP_3760 (  );
sky130_fd_sc_hd__tap_1 TAP_3761 (  );
sky130_fd_sc_hd__tap_1 TAP_3762 (  );
sky130_fd_sc_hd__tap_1 TAP_3763 (  );
sky130_fd_sc_hd__tap_1 TAP_3764 (  );
sky130_fd_sc_hd__tap_1 TAP_3765 (  );
sky130_fd_sc_hd__tap_1 TAP_3766 (  );
sky130_fd_sc_hd__tap_1 TAP_3767 (  );
sky130_fd_sc_hd__tap_1 TAP_3768 (  );
sky130_fd_sc_hd__tap_1 TAP_3769 (  );
sky130_fd_sc_hd__tap_1 TAP_3770 (  );
sky130_fd_sc_hd__tap_1 TAP_3771 (  );
sky130_fd_sc_hd__tap_1 TAP_3772 (  );
sky130_fd_sc_hd__tap_1 TAP_3773 (  );
sky130_fd_sc_hd__tap_1 TAP_3774 (  );
sky130_fd_sc_hd__tap_1 TAP_3775 (  );
sky130_fd_sc_hd__tap_1 TAP_3776 (  );
sky130_fd_sc_hd__tap_1 TAP_3777 (  );
sky130_fd_sc_hd__tap_1 TAP_3778 (  );
sky130_fd_sc_hd__tap_1 TAP_3779 (  );
sky130_fd_sc_hd__tap_1 TAP_3780 (  );
sky130_fd_sc_hd__tap_1 TAP_3781 (  );
sky130_fd_sc_hd__tap_1 TAP_3782 (  );
sky130_fd_sc_hd__tap_1 TAP_3783 (  );
sky130_fd_sc_hd__tap_1 TAP_3784 (  );
sky130_fd_sc_hd__tap_1 TAP_3785 (  );
sky130_fd_sc_hd__tap_1 TAP_3786 (  );
sky130_fd_sc_hd__tap_1 TAP_3787 (  );
sky130_fd_sc_hd__tap_1 TAP_3788 (  );
sky130_fd_sc_hd__tap_1 TAP_3789 (  );
sky130_fd_sc_hd__tap_1 TAP_3790 (  );
sky130_fd_sc_hd__tap_1 TAP_3791 (  );
sky130_fd_sc_hd__tap_1 TAP_3792 (  );
sky130_fd_sc_hd__tap_1 TAP_3793 (  );
sky130_fd_sc_hd__tap_1 TAP_3794 (  );
sky130_fd_sc_hd__tap_1 TAP_3795 (  );
sky130_fd_sc_hd__tap_1 TAP_3796 (  );
sky130_fd_sc_hd__tap_1 TAP_3797 (  );
sky130_fd_sc_hd__tap_1 TAP_3798 (  );
sky130_fd_sc_hd__tap_1 TAP_3799 (  );
sky130_fd_sc_hd__tap_1 TAP_3800 (  );
sky130_fd_sc_hd__tap_1 TAP_3801 (  );
sky130_fd_sc_hd__tap_1 TAP_3802 (  );
sky130_fd_sc_hd__tap_1 TAP_3803 (  );
sky130_fd_sc_hd__tap_1 TAP_3804 (  );
sky130_fd_sc_hd__tap_1 TAP_3805 (  );
sky130_fd_sc_hd__tap_1 TAP_3806 (  );
sky130_fd_sc_hd__tap_1 TAP_3807 (  );
sky130_fd_sc_hd__tap_1 TAP_3808 (  );
sky130_fd_sc_hd__tap_1 TAP_3809 (  );
sky130_fd_sc_hd__tap_1 TAP_3810 (  );
sky130_fd_sc_hd__tap_1 TAP_3811 (  );
sky130_fd_sc_hd__tap_1 TAP_3812 (  );
sky130_fd_sc_hd__tap_1 TAP_3813 (  );
sky130_fd_sc_hd__tap_1 TAP_3814 (  );
sky130_fd_sc_hd__tap_1 TAP_3815 (  );
sky130_fd_sc_hd__tap_1 TAP_3816 (  );
sky130_fd_sc_hd__tap_1 TAP_3817 (  );
sky130_fd_sc_hd__tap_1 TAP_3818 (  );
sky130_fd_sc_hd__tap_1 TAP_3819 (  );
sky130_fd_sc_hd__tap_1 TAP_3820 (  );
sky130_fd_sc_hd__tap_1 TAP_3821 (  );
sky130_fd_sc_hd__tap_1 TAP_3822 (  );
sky130_fd_sc_hd__tap_1 TAP_3823 (  );
sky130_fd_sc_hd__tap_1 TAP_3824 (  );
sky130_fd_sc_hd__tap_1 TAP_3825 (  );
sky130_fd_sc_hd__tap_1 TAP_3826 (  );
sky130_fd_sc_hd__tap_1 TAP_3827 (  );
sky130_fd_sc_hd__tap_1 TAP_3828 (  );
sky130_fd_sc_hd__tap_1 TAP_3829 (  );
sky130_fd_sc_hd__tap_1 TAP_3830 (  );
sky130_fd_sc_hd__tap_1 TAP_3831 (  );
sky130_fd_sc_hd__tap_1 TAP_3832 (  );
sky130_fd_sc_hd__tap_1 TAP_3833 (  );
sky130_fd_sc_hd__tap_1 TAP_3834 (  );
sky130_fd_sc_hd__tap_1 TAP_3835 (  );
sky130_fd_sc_hd__tap_1 TAP_3836 (  );
sky130_fd_sc_hd__tap_1 TAP_3837 (  );
sky130_fd_sc_hd__tap_1 TAP_3838 (  );
sky130_fd_sc_hd__tap_1 TAP_3839 (  );
sky130_fd_sc_hd__tap_1 TAP_3840 (  );
sky130_fd_sc_hd__tap_1 TAP_3841 (  );
sky130_fd_sc_hd__tap_1 TAP_3842 (  );
sky130_fd_sc_hd__tap_1 TAP_3843 (  );
sky130_fd_sc_hd__tap_1 TAP_3844 (  );
sky130_fd_sc_hd__tap_1 TAP_3845 (  );
sky130_fd_sc_hd__tap_1 TAP_3846 (  );
sky130_fd_sc_hd__tap_1 TAP_3847 (  );
sky130_fd_sc_hd__tap_1 TAP_3848 (  );
sky130_fd_sc_hd__tap_1 TAP_3849 (  );
sky130_fd_sc_hd__tap_1 TAP_3850 (  );
sky130_fd_sc_hd__tap_1 TAP_3851 (  );
sky130_fd_sc_hd__tap_1 TAP_3852 (  );
sky130_fd_sc_hd__tap_1 TAP_3853 (  );
sky130_fd_sc_hd__tap_1 TAP_3854 (  );
sky130_fd_sc_hd__tap_1 TAP_3855 (  );
sky130_fd_sc_hd__tap_1 TAP_3856 (  );
sky130_fd_sc_hd__tap_1 TAP_3857 (  );
sky130_fd_sc_hd__tap_1 TAP_3858 (  );
sky130_fd_sc_hd__tap_1 TAP_3859 (  );
sky130_fd_sc_hd__tap_1 TAP_3860 (  );
sky130_fd_sc_hd__tap_1 TAP_3861 (  );
sky130_fd_sc_hd__tap_1 TAP_3862 (  );
sky130_fd_sc_hd__tap_1 TAP_3863 (  );
sky130_fd_sc_hd__tap_1 TAP_3864 (  );
sky130_fd_sc_hd__tap_1 TAP_3865 (  );
sky130_fd_sc_hd__tap_1 TAP_3866 (  );
sky130_fd_sc_hd__tap_1 TAP_3867 (  );
sky130_fd_sc_hd__tap_1 TAP_3868 (  );
sky130_fd_sc_hd__tap_1 TAP_3869 (  );
sky130_fd_sc_hd__tap_1 TAP_3870 (  );
sky130_fd_sc_hd__tap_1 TAP_3871 (  );
sky130_fd_sc_hd__tap_1 TAP_3872 (  );
sky130_fd_sc_hd__tap_1 TAP_3873 (  );
sky130_fd_sc_hd__tap_1 TAP_3874 (  );
sky130_fd_sc_hd__tap_1 TAP_3875 (  );
sky130_fd_sc_hd__tap_1 TAP_3876 (  );
sky130_fd_sc_hd__tap_1 TAP_3877 (  );
sky130_fd_sc_hd__tap_1 TAP_3878 (  );
sky130_fd_sc_hd__tap_1 TAP_3879 (  );
sky130_fd_sc_hd__tap_1 TAP_3880 (  );
sky130_fd_sc_hd__tap_1 TAP_3881 (  );
sky130_fd_sc_hd__tap_1 TAP_3882 (  );
sky130_fd_sc_hd__tap_1 TAP_3883 (  );
sky130_fd_sc_hd__tap_1 TAP_3884 (  );
sky130_fd_sc_hd__tap_1 TAP_3885 (  );
sky130_fd_sc_hd__tap_1 TAP_3886 (  );
sky130_fd_sc_hd__tap_1 TAP_3887 (  );
sky130_fd_sc_hd__tap_1 TAP_3888 (  );
sky130_fd_sc_hd__tap_1 TAP_3889 (  );
sky130_fd_sc_hd__tap_1 TAP_3890 (  );
sky130_fd_sc_hd__tap_1 TAP_3891 (  );
sky130_fd_sc_hd__tap_1 TAP_3892 (  );
sky130_fd_sc_hd__tap_1 TAP_3893 (  );
sky130_fd_sc_hd__tap_1 TAP_3894 (  );
sky130_fd_sc_hd__tap_1 TAP_3895 (  );
sky130_fd_sc_hd__tap_1 TAP_3896 (  );
sky130_fd_sc_hd__tap_1 TAP_3897 (  );
sky130_fd_sc_hd__tap_1 TAP_3898 (  );
sky130_fd_sc_hd__tap_1 TAP_3899 (  );
sky130_fd_sc_hd__tap_1 TAP_3900 (  );
sky130_fd_sc_hd__tap_1 TAP_3901 (  );
sky130_fd_sc_hd__tap_1 TAP_3902 (  );
sky130_fd_sc_hd__tap_1 TAP_3903 (  );
sky130_fd_sc_hd__tap_1 TAP_3904 (  );
sky130_fd_sc_hd__tap_1 TAP_3905 (  );
sky130_fd_sc_hd__tap_1 TAP_3906 (  );
sky130_fd_sc_hd__tap_1 TAP_3907 (  );
sky130_fd_sc_hd__tap_1 TAP_3908 (  );
sky130_fd_sc_hd__tap_1 TAP_3909 (  );
sky130_fd_sc_hd__tap_1 TAP_3910 (  );
sky130_fd_sc_hd__tap_1 TAP_3911 (  );
sky130_fd_sc_hd__tap_1 TAP_3912 (  );
sky130_fd_sc_hd__tap_1 TAP_3913 (  );
sky130_fd_sc_hd__tap_1 TAP_3914 (  );
sky130_fd_sc_hd__tap_1 TAP_3915 (  );
sky130_fd_sc_hd__tap_1 TAP_3916 (  );
sky130_fd_sc_hd__tap_1 TAP_3917 (  );
sky130_fd_sc_hd__tap_1 TAP_3918 (  );
sky130_fd_sc_hd__tap_1 TAP_3919 (  );
sky130_fd_sc_hd__tap_1 TAP_3920 (  );
sky130_fd_sc_hd__tap_1 TAP_3921 (  );
sky130_fd_sc_hd__tap_1 TAP_3922 (  );
sky130_fd_sc_hd__tap_1 TAP_3923 (  );
sky130_fd_sc_hd__tap_1 TAP_3924 (  );
sky130_fd_sc_hd__tap_1 TAP_3925 (  );
sky130_fd_sc_hd__tap_1 TAP_3926 (  );
sky130_fd_sc_hd__tap_1 TAP_3927 (  );
sky130_fd_sc_hd__tap_1 TAP_3928 (  );
sky130_fd_sc_hd__tap_1 TAP_3929 (  );
sky130_fd_sc_hd__tap_1 TAP_3930 (  );
sky130_fd_sc_hd__tap_1 TAP_3931 (  );
sky130_fd_sc_hd__tap_1 TAP_3932 (  );
sky130_fd_sc_hd__tap_1 TAP_3933 (  );
sky130_fd_sc_hd__tap_1 TAP_3934 (  );
sky130_fd_sc_hd__tap_1 TAP_3935 (  );
sky130_fd_sc_hd__tap_1 TAP_3936 (  );
sky130_fd_sc_hd__tap_1 TAP_3937 (  );
sky130_fd_sc_hd__tap_1 TAP_3938 (  );
sky130_fd_sc_hd__tap_1 TAP_3939 (  );
sky130_fd_sc_hd__tap_1 TAP_3940 (  );
sky130_fd_sc_hd__tap_1 TAP_3941 (  );
sky130_fd_sc_hd__tap_1 TAP_3942 (  );
sky130_fd_sc_hd__tap_1 TAP_3943 (  );
sky130_fd_sc_hd__tap_1 TAP_3944 (  );
sky130_fd_sc_hd__tap_1 TAP_3945 (  );
sky130_fd_sc_hd__tap_1 TAP_3946 (  );
sky130_fd_sc_hd__tap_1 TAP_3947 (  );
sky130_fd_sc_hd__tap_1 TAP_3948 (  );
sky130_fd_sc_hd__tap_1 TAP_3949 (  );
sky130_fd_sc_hd__tap_1 TAP_3950 (  );
sky130_fd_sc_hd__tap_1 TAP_3951 (  );
sky130_fd_sc_hd__tap_1 TAP_3952 (  );
sky130_fd_sc_hd__tap_1 TAP_3953 (  );
sky130_fd_sc_hd__tap_1 TAP_3954 (  );
sky130_fd_sc_hd__tap_1 TAP_3955 (  );
sky130_fd_sc_hd__tap_1 TAP_3956 (  );
sky130_fd_sc_hd__tap_1 TAP_3957 (  );
sky130_fd_sc_hd__tap_1 TAP_3958 (  );
sky130_fd_sc_hd__tap_1 TAP_3959 (  );
sky130_fd_sc_hd__tap_1 TAP_3960 (  );
sky130_fd_sc_hd__tap_1 TAP_3961 (  );
sky130_fd_sc_hd__tap_1 TAP_3962 (  );
sky130_fd_sc_hd__tap_1 TAP_3963 (  );
sky130_fd_sc_hd__tap_1 TAP_3964 (  );
sky130_fd_sc_hd__tap_1 TAP_3965 (  );
sky130_fd_sc_hd__tap_1 TAP_3966 (  );
sky130_fd_sc_hd__tap_1 TAP_3967 (  );
sky130_fd_sc_hd__tap_1 TAP_3968 (  );
sky130_fd_sc_hd__tap_1 TAP_3969 (  );
sky130_fd_sc_hd__tap_1 TAP_3970 (  );
sky130_fd_sc_hd__tap_1 TAP_3971 (  );
sky130_fd_sc_hd__tap_1 TAP_3972 (  );
sky130_fd_sc_hd__tap_1 TAP_3973 (  );
sky130_fd_sc_hd__tap_1 TAP_3974 (  );
sky130_fd_sc_hd__tap_1 TAP_3975 (  );
sky130_fd_sc_hd__tap_1 TAP_3976 (  );
sky130_fd_sc_hd__tap_1 TAP_3977 (  );
sky130_fd_sc_hd__tap_1 TAP_3978 (  );
sky130_fd_sc_hd__tap_1 TAP_3979 (  );
sky130_fd_sc_hd__tap_1 TAP_3980 (  );
sky130_fd_sc_hd__tap_1 TAP_3981 (  );
sky130_fd_sc_hd__tap_1 TAP_3982 (  );
sky130_fd_sc_hd__tap_1 TAP_3983 (  );
sky130_fd_sc_hd__tap_1 TAP_3984 (  );
sky130_fd_sc_hd__tap_1 TAP_3985 (  );
sky130_fd_sc_hd__tap_1 TAP_3986 (  );
sky130_fd_sc_hd__tap_1 TAP_3987 (  );
sky130_fd_sc_hd__tap_1 TAP_3988 (  );
sky130_fd_sc_hd__tap_1 TAP_3989 (  );
sky130_fd_sc_hd__tap_1 TAP_3990 (  );
sky130_fd_sc_hd__tap_1 TAP_3991 (  );
sky130_fd_sc_hd__tap_1 TAP_3992 (  );
sky130_fd_sc_hd__tap_1 TAP_3993 (  );
sky130_fd_sc_hd__tap_1 TAP_3994 (  );
sky130_fd_sc_hd__tap_1 TAP_3995 (  );
sky130_fd_sc_hd__tap_1 TAP_3996 (  );
sky130_fd_sc_hd__tap_1 TAP_3997 (  );
sky130_fd_sc_hd__tap_1 TAP_3998 (  );
sky130_fd_sc_hd__tap_1 TAP_3999 (  );
sky130_fd_sc_hd__tap_1 TAP_4000 (  );
sky130_fd_sc_hd__tap_1 TAP_4001 (  );
sky130_fd_sc_hd__tap_1 TAP_4002 (  );
sky130_fd_sc_hd__tap_1 TAP_4003 (  );
sky130_fd_sc_hd__tap_1 TAP_4004 (  );
sky130_fd_sc_hd__tap_1 TAP_4005 (  );
sky130_fd_sc_hd__tap_1 TAP_4006 (  );
sky130_fd_sc_hd__tap_1 TAP_4007 (  );
sky130_fd_sc_hd__tap_1 TAP_4008 (  );
sky130_fd_sc_hd__tap_1 TAP_4009 (  );
sky130_fd_sc_hd__tap_1 TAP_4010 (  );
sky130_fd_sc_hd__tap_1 TAP_4011 (  );
sky130_fd_sc_hd__tap_1 TAP_4012 (  );
sky130_fd_sc_hd__tap_1 TAP_4013 (  );
sky130_fd_sc_hd__tap_1 TAP_4014 (  );
sky130_fd_sc_hd__tap_1 TAP_4015 (  );
sky130_fd_sc_hd__tap_1 TAP_4016 (  );
sky130_fd_sc_hd__tap_1 TAP_4017 (  );
sky130_fd_sc_hd__tap_1 TAP_4018 (  );
sky130_fd_sc_hd__tap_1 TAP_4019 (  );
sky130_fd_sc_hd__tap_1 TAP_4020 (  );
sky130_fd_sc_hd__tap_1 TAP_4021 (  );
sky130_fd_sc_hd__tap_1 TAP_4022 (  );
sky130_fd_sc_hd__tap_1 TAP_4023 (  );
sky130_fd_sc_hd__tap_1 TAP_4024 (  );
sky130_fd_sc_hd__tap_1 TAP_4025 (  );
sky130_fd_sc_hd__tap_1 TAP_4026 (  );
sky130_fd_sc_hd__tap_1 TAP_4027 (  );
sky130_fd_sc_hd__tap_1 TAP_4028 (  );
sky130_fd_sc_hd__tap_1 TAP_4029 (  );
sky130_fd_sc_hd__tap_1 TAP_4030 (  );
sky130_fd_sc_hd__tap_1 TAP_4031 (  );
sky130_fd_sc_hd__tap_1 TAP_4032 (  );
sky130_fd_sc_hd__tap_1 TAP_4033 (  );
sky130_fd_sc_hd__tap_1 TAP_4034 (  );
sky130_fd_sc_hd__tap_1 TAP_4035 (  );
sky130_fd_sc_hd__tap_1 TAP_4036 (  );
sky130_fd_sc_hd__tap_1 TAP_4037 (  );
sky130_fd_sc_hd__tap_1 TAP_4038 (  );
sky130_fd_sc_hd__tap_1 TAP_4039 (  );
sky130_fd_sc_hd__tap_1 TAP_4040 (  );
sky130_fd_sc_hd__tap_1 TAP_4041 (  );
sky130_fd_sc_hd__tap_1 TAP_4042 (  );
sky130_fd_sc_hd__tap_1 TAP_4043 (  );
sky130_fd_sc_hd__tap_1 TAP_4044 (  );
sky130_fd_sc_hd__tap_1 TAP_4045 (  );
sky130_fd_sc_hd__tap_1 TAP_4046 (  );
sky130_fd_sc_hd__tap_1 TAP_4047 (  );
sky130_fd_sc_hd__tap_1 TAP_4048 (  );
sky130_fd_sc_hd__tap_1 TAP_4049 (  );
sky130_fd_sc_hd__tap_1 TAP_4050 (  );
sky130_fd_sc_hd__tap_1 TAP_4051 (  );
sky130_fd_sc_hd__tap_1 TAP_4052 (  );
sky130_fd_sc_hd__tap_1 TAP_4053 (  );
sky130_fd_sc_hd__tap_1 TAP_4054 (  );
sky130_fd_sc_hd__tap_1 TAP_4055 (  );
sky130_fd_sc_hd__tap_1 TAP_4056 (  );
sky130_fd_sc_hd__tap_1 TAP_4057 (  );
sky130_fd_sc_hd__tap_1 TAP_4058 (  );
sky130_fd_sc_hd__tap_1 TAP_4059 (  );
sky130_fd_sc_hd__tap_1 TAP_4060 (  );
sky130_fd_sc_hd__tap_1 TAP_4061 (  );
sky130_fd_sc_hd__tap_1 TAP_4062 (  );
sky130_fd_sc_hd__tap_1 TAP_4063 (  );
sky130_fd_sc_hd__tap_1 TAP_4064 (  );
sky130_fd_sc_hd__tap_1 TAP_4065 (  );
sky130_fd_sc_hd__tap_1 TAP_4066 (  );
sky130_fd_sc_hd__tap_1 TAP_4067 (  );
sky130_fd_sc_hd__tap_1 TAP_4068 (  );
sky130_fd_sc_hd__tap_1 TAP_4069 (  );
sky130_fd_sc_hd__tap_1 TAP_4070 (  );
sky130_fd_sc_hd__tap_1 TAP_4071 (  );
sky130_fd_sc_hd__tap_1 TAP_4072 (  );
sky130_fd_sc_hd__tap_1 TAP_4073 (  );
sky130_fd_sc_hd__tap_1 TAP_4074 (  );
sky130_fd_sc_hd__tap_1 TAP_4075 (  );
sky130_fd_sc_hd__tap_1 TAP_4076 (  );
sky130_fd_sc_hd__tap_1 TAP_4077 (  );
sky130_fd_sc_hd__tap_1 TAP_4078 (  );
sky130_fd_sc_hd__tap_1 TAP_4079 (  );
sky130_fd_sc_hd__tap_1 TAP_4080 (  );
sky130_fd_sc_hd__tap_1 TAP_4081 (  );
sky130_fd_sc_hd__tap_1 TAP_4082 (  );
sky130_fd_sc_hd__tap_1 TAP_4083 (  );
sky130_fd_sc_hd__tap_1 TAP_4084 (  );
sky130_fd_sc_hd__tap_1 TAP_4085 (  );
sky130_fd_sc_hd__tap_1 TAP_4086 (  );
sky130_fd_sc_hd__tap_1 TAP_4087 (  );
sky130_fd_sc_hd__tap_1 TAP_4088 (  );
sky130_fd_sc_hd__tap_1 TAP_4089 (  );
sky130_fd_sc_hd__tap_1 TAP_4090 (  );
sky130_fd_sc_hd__tap_1 TAP_4091 (  );
sky130_fd_sc_hd__tap_1 TAP_4092 (  );
sky130_fd_sc_hd__tap_1 TAP_4093 (  );
sky130_fd_sc_hd__tap_1 TAP_4094 (  );
sky130_fd_sc_hd__tap_1 TAP_4095 (  );
sky130_fd_sc_hd__tap_1 TAP_4096 (  );
sky130_fd_sc_hd__tap_1 TAP_4097 (  );
sky130_fd_sc_hd__tap_1 TAP_4098 (  );
sky130_fd_sc_hd__tap_1 TAP_4099 (  );
sky130_fd_sc_hd__tap_1 TAP_4100 (  );
sky130_fd_sc_hd__tap_1 TAP_4101 (  );
sky130_fd_sc_hd__tap_1 TAP_4102 (  );
sky130_fd_sc_hd__tap_1 TAP_4103 (  );
sky130_fd_sc_hd__tap_1 TAP_4104 (  );
sky130_fd_sc_hd__tap_1 TAP_4105 (  );
sky130_fd_sc_hd__tap_1 TAP_4106 (  );
sky130_fd_sc_hd__tap_1 TAP_4107 (  );
sky130_fd_sc_hd__tap_1 TAP_4108 (  );
sky130_fd_sc_hd__tap_1 TAP_4109 (  );
sky130_fd_sc_hd__tap_1 TAP_4110 (  );
sky130_fd_sc_hd__tap_1 TAP_4111 (  );
sky130_fd_sc_hd__tap_1 TAP_4112 (  );
sky130_fd_sc_hd__tap_1 TAP_4113 (  );
sky130_fd_sc_hd__tap_1 TAP_4114 (  );
sky130_fd_sc_hd__tap_1 TAP_4115 (  );
sky130_fd_sc_hd__tap_1 TAP_4116 (  );
sky130_fd_sc_hd__tap_1 TAP_4117 (  );
sky130_fd_sc_hd__tap_1 TAP_4118 (  );
sky130_fd_sc_hd__tap_1 TAP_4119 (  );
sky130_fd_sc_hd__tap_1 TAP_4120 (  );
sky130_fd_sc_hd__tap_1 TAP_4121 (  );
sky130_fd_sc_hd__tap_1 TAP_4122 (  );
sky130_fd_sc_hd__tap_1 TAP_4123 (  );
sky130_fd_sc_hd__tap_1 TAP_4124 (  );
sky130_fd_sc_hd__tap_1 TAP_4125 (  );
sky130_fd_sc_hd__tap_1 TAP_4126 (  );
sky130_fd_sc_hd__tap_1 TAP_4127 (  );
sky130_fd_sc_hd__tap_1 TAP_4128 (  );
sky130_fd_sc_hd__tap_1 TAP_4129 (  );
sky130_fd_sc_hd__tap_1 TAP_4130 (  );
sky130_fd_sc_hd__tap_1 TAP_4131 (  );
sky130_fd_sc_hd__tap_1 TAP_4132 (  );
sky130_fd_sc_hd__tap_1 TAP_4133 (  );
sky130_fd_sc_hd__tap_1 TAP_4134 (  );
sky130_fd_sc_hd__tap_1 TAP_4135 (  );
sky130_fd_sc_hd__tap_1 TAP_4136 (  );
sky130_fd_sc_hd__tap_1 TAP_4137 (  );
sky130_fd_sc_hd__tap_1 TAP_4138 (  );
sky130_fd_sc_hd__tap_1 TAP_4139 (  );
sky130_fd_sc_hd__tap_1 TAP_4140 (  );
sky130_fd_sc_hd__tap_1 TAP_4141 (  );
sky130_fd_sc_hd__tap_1 TAP_4142 (  );
sky130_fd_sc_hd__tap_1 TAP_4143 (  );
sky130_fd_sc_hd__tap_1 TAP_4144 (  );
sky130_fd_sc_hd__tap_1 TAP_4145 (  );
sky130_fd_sc_hd__tap_1 TAP_4146 (  );
sky130_fd_sc_hd__tap_1 TAP_4147 (  );
sky130_fd_sc_hd__tap_1 TAP_4148 (  );
sky130_fd_sc_hd__tap_1 TAP_4149 (  );
sky130_fd_sc_hd__tap_1 TAP_4150 (  );
sky130_fd_sc_hd__tap_1 TAP_4151 (  );
sky130_fd_sc_hd__tap_1 TAP_4152 (  );
sky130_fd_sc_hd__tap_1 TAP_4153 (  );
sky130_fd_sc_hd__tap_1 TAP_4154 (  );
sky130_fd_sc_hd__tap_1 TAP_4155 (  );
sky130_fd_sc_hd__tap_1 TAP_4156 (  );
sky130_fd_sc_hd__tap_1 TAP_4157 (  );
sky130_fd_sc_hd__tap_1 TAP_4158 (  );
sky130_fd_sc_hd__tap_1 TAP_4159 (  );
sky130_fd_sc_hd__tap_1 TAP_4160 (  );
sky130_fd_sc_hd__tap_1 TAP_4161 (  );
sky130_fd_sc_hd__tap_1 TAP_4162 (  );
sky130_fd_sc_hd__tap_1 TAP_4163 (  );
sky130_fd_sc_hd__tap_1 TAP_4164 (  );
sky130_fd_sc_hd__tap_1 TAP_4165 (  );
sky130_fd_sc_hd__tap_1 TAP_4166 (  );
sky130_fd_sc_hd__tap_1 TAP_4167 (  );
sky130_fd_sc_hd__tap_1 TAP_4168 (  );
sky130_fd_sc_hd__tap_1 TAP_4169 (  );
sky130_fd_sc_hd__tap_1 TAP_4170 (  );
sky130_fd_sc_hd__tap_1 TAP_4171 (  );
sky130_fd_sc_hd__tap_1 TAP_4172 (  );
sky130_fd_sc_hd__tap_1 TAP_4173 (  );
sky130_fd_sc_hd__tap_1 TAP_4174 (  );
sky130_fd_sc_hd__tap_1 TAP_4175 (  );
sky130_fd_sc_hd__tap_1 TAP_4176 (  );
sky130_fd_sc_hd__tap_1 TAP_4177 (  );
sky130_fd_sc_hd__tap_1 TAP_4178 (  );
sky130_fd_sc_hd__tap_1 TAP_4179 (  );
sky130_fd_sc_hd__tap_1 TAP_4180 (  );
sky130_fd_sc_hd__tap_1 TAP_4181 (  );
sky130_fd_sc_hd__tap_1 TAP_4182 (  );
sky130_fd_sc_hd__tap_1 TAP_4183 (  );
sky130_fd_sc_hd__tap_1 TAP_4184 (  );
sky130_fd_sc_hd__tap_1 TAP_4185 (  );
sky130_fd_sc_hd__tap_1 TAP_4186 (  );
sky130_fd_sc_hd__tap_1 TAP_4187 (  );
sky130_fd_sc_hd__tap_1 TAP_4188 (  );
sky130_fd_sc_hd__tap_1 TAP_4189 (  );
sky130_fd_sc_hd__tap_1 TAP_4190 (  );
sky130_fd_sc_hd__tap_1 TAP_4191 (  );
sky130_fd_sc_hd__tap_1 TAP_4192 (  );
sky130_fd_sc_hd__tap_1 TAP_4193 (  );
sky130_fd_sc_hd__tap_1 TAP_4194 (  );
sky130_fd_sc_hd__tap_1 TAP_4195 (  );
sky130_fd_sc_hd__tap_1 TAP_4196 (  );
sky130_fd_sc_hd__tap_1 TAP_4197 (  );
sky130_fd_sc_hd__tap_1 TAP_4198 (  );
sky130_fd_sc_hd__tap_1 TAP_4199 (  );
sky130_fd_sc_hd__tap_1 TAP_4200 (  );
sky130_fd_sc_hd__tap_1 TAP_4201 (  );
sky130_fd_sc_hd__tap_1 TAP_4202 (  );
sky130_fd_sc_hd__tap_1 TAP_4203 (  );
sky130_fd_sc_hd__tap_1 TAP_4204 (  );
sky130_fd_sc_hd__tap_1 TAP_4205 (  );
sky130_fd_sc_hd__tap_1 TAP_4206 (  );
sky130_fd_sc_hd__tap_1 TAP_4207 (  );
sky130_fd_sc_hd__tap_1 TAP_4208 (  );
sky130_fd_sc_hd__tap_1 TAP_4209 (  );
sky130_fd_sc_hd__tap_1 TAP_4210 (  );
sky130_fd_sc_hd__tap_1 TAP_4211 (  );
sky130_fd_sc_hd__tap_1 TAP_4212 (  );
sky130_fd_sc_hd__tap_1 TAP_4213 (  );
sky130_fd_sc_hd__tap_1 TAP_4214 (  );
sky130_fd_sc_hd__tap_1 TAP_4215 (  );
sky130_fd_sc_hd__tap_1 TAP_4216 (  );
sky130_fd_sc_hd__tap_1 TAP_4217 (  );
sky130_fd_sc_hd__tap_1 TAP_4218 (  );
sky130_fd_sc_hd__tap_1 TAP_4219 (  );
sky130_fd_sc_hd__tap_1 TAP_4220 (  );
sky130_fd_sc_hd__tap_1 TAP_4221 (  );
sky130_fd_sc_hd__tap_1 TAP_4222 (  );
sky130_fd_sc_hd__tap_1 TAP_4223 (  );
sky130_fd_sc_hd__tap_1 TAP_4224 (  );
sky130_fd_sc_hd__tap_1 TAP_4225 (  );
sky130_fd_sc_hd__tap_1 TAP_4226 (  );
sky130_fd_sc_hd__tap_1 TAP_4227 (  );
sky130_fd_sc_hd__tap_1 TAP_4228 (  );
sky130_fd_sc_hd__tap_1 TAP_4229 (  );
sky130_fd_sc_hd__tap_1 TAP_4230 (  );
sky130_fd_sc_hd__tap_1 TAP_4231 (  );
sky130_fd_sc_hd__tap_1 TAP_4232 (  );
sky130_fd_sc_hd__tap_1 TAP_4233 (  );
sky130_fd_sc_hd__tap_1 TAP_4234 (  );
sky130_fd_sc_hd__tap_1 TAP_4235 (  );
sky130_fd_sc_hd__tap_1 TAP_4236 (  );
sky130_fd_sc_hd__tap_1 TAP_4237 (  );
sky130_fd_sc_hd__tap_1 TAP_4238 (  );
sky130_fd_sc_hd__tap_1 TAP_4239 (  );
sky130_fd_sc_hd__tap_1 TAP_4240 (  );
sky130_fd_sc_hd__tap_1 TAP_4241 (  );
sky130_fd_sc_hd__tap_1 TAP_4242 (  );
sky130_fd_sc_hd__tap_1 TAP_4243 (  );
sky130_fd_sc_hd__tap_1 TAP_4244 (  );
sky130_fd_sc_hd__tap_1 TAP_4245 (  );
sky130_fd_sc_hd__tap_1 TAP_4246 (  );
sky130_fd_sc_hd__tap_1 TAP_4247 (  );
sky130_fd_sc_hd__tap_1 TAP_4248 (  );
sky130_fd_sc_hd__tap_1 TAP_4249 (  );
sky130_fd_sc_hd__tap_1 TAP_4250 (  );
sky130_fd_sc_hd__tap_1 TAP_4251 (  );
sky130_fd_sc_hd__tap_1 TAP_4252 (  );
sky130_fd_sc_hd__tap_1 TAP_4253 (  );
sky130_fd_sc_hd__tap_1 TAP_4254 (  );
sky130_fd_sc_hd__tap_1 TAP_4255 (  );
sky130_fd_sc_hd__tap_1 TAP_4256 (  );
sky130_fd_sc_hd__tap_1 TAP_4257 (  );
sky130_fd_sc_hd__tap_1 TAP_4258 (  );
sky130_fd_sc_hd__tap_1 TAP_4259 (  );
sky130_fd_sc_hd__tap_1 TAP_4260 (  );
sky130_fd_sc_hd__tap_1 TAP_4261 (  );
sky130_fd_sc_hd__tap_1 TAP_4262 (  );
sky130_fd_sc_hd__tap_1 TAP_4263 (  );
sky130_fd_sc_hd__tap_1 TAP_4264 (  );
sky130_fd_sc_hd__tap_1 TAP_4265 (  );
sky130_fd_sc_hd__tap_1 TAP_4266 (  );
sky130_fd_sc_hd__tap_1 TAP_4267 (  );
sky130_fd_sc_hd__tap_1 TAP_4268 (  );
sky130_fd_sc_hd__tap_1 TAP_4269 (  );
sky130_fd_sc_hd__tap_1 TAP_4270 (  );
sky130_fd_sc_hd__tap_1 TAP_4271 (  );
sky130_fd_sc_hd__tap_1 TAP_4272 (  );
sky130_fd_sc_hd__tap_1 TAP_4273 (  );
sky130_fd_sc_hd__tap_1 TAP_4274 (  );
sky130_fd_sc_hd__tap_1 TAP_4275 (  );
sky130_fd_sc_hd__tap_1 TAP_4276 (  );
sky130_fd_sc_hd__tap_1 TAP_4277 (  );
sky130_fd_sc_hd__tap_1 TAP_4278 (  );
sky130_fd_sc_hd__tap_1 TAP_4279 (  );
sky130_fd_sc_hd__tap_1 TAP_4280 (  );
sky130_fd_sc_hd__tap_1 TAP_4281 (  );
sky130_fd_sc_hd__tap_1 TAP_4282 (  );
sky130_fd_sc_hd__tap_1 TAP_4283 (  );
sky130_fd_sc_hd__tap_1 TAP_4284 (  );
sky130_fd_sc_hd__tap_1 TAP_4285 (  );
sky130_fd_sc_hd__tap_1 TAP_4286 (  );
sky130_fd_sc_hd__tap_1 TAP_4287 (  );
sky130_fd_sc_hd__tap_1 TAP_4288 (  );
sky130_fd_sc_hd__tap_1 TAP_4289 (  );
sky130_fd_sc_hd__tap_1 TAP_4290 (  );
sky130_fd_sc_hd__tap_1 TAP_4291 (  );
sky130_fd_sc_hd__tap_1 TAP_4292 (  );
sky130_fd_sc_hd__tap_1 TAP_4293 (  );
sky130_fd_sc_hd__tap_1 TAP_4294 (  );
sky130_fd_sc_hd__tap_1 TAP_4295 (  );
sky130_fd_sc_hd__tap_1 TAP_4296 (  );
sky130_fd_sc_hd__tap_1 TAP_4297 (  );
sky130_fd_sc_hd__tap_1 TAP_4298 (  );
sky130_fd_sc_hd__tap_1 TAP_4299 (  );
sky130_fd_sc_hd__tap_1 TAP_4300 (  );
sky130_fd_sc_hd__tap_1 TAP_4301 (  );
sky130_fd_sc_hd__tap_1 TAP_4302 (  );
sky130_fd_sc_hd__tap_1 TAP_4303 (  );
sky130_fd_sc_hd__tap_1 TAP_4304 (  );
sky130_fd_sc_hd__tap_1 TAP_4305 (  );
sky130_fd_sc_hd__tap_1 TAP_4306 (  );
sky130_fd_sc_hd__tap_1 TAP_4307 (  );
sky130_fd_sc_hd__tap_1 TAP_4308 (  );
sky130_fd_sc_hd__tap_1 TAP_4309 (  );
sky130_fd_sc_hd__tap_1 TAP_4310 (  );
sky130_fd_sc_hd__tap_1 TAP_4311 (  );
sky130_fd_sc_hd__tap_1 TAP_4312 (  );
sky130_fd_sc_hd__tap_1 TAP_4313 (  );
sky130_fd_sc_hd__tap_1 TAP_4314 (  );
sky130_fd_sc_hd__tap_1 TAP_4315 (  );
sky130_fd_sc_hd__tap_1 TAP_4316 (  );
sky130_fd_sc_hd__tap_1 TAP_4317 (  );
sky130_fd_sc_hd__tap_1 TAP_4318 (  );
sky130_fd_sc_hd__tap_1 TAP_4319 (  );
sky130_fd_sc_hd__tap_1 TAP_4320 (  );
sky130_fd_sc_hd__tap_1 TAP_4321 (  );
sky130_fd_sc_hd__tap_1 TAP_4322 (  );
sky130_fd_sc_hd__tap_1 TAP_4323 (  );
sky130_fd_sc_hd__tap_1 TAP_4324 (  );
sky130_fd_sc_hd__tap_1 TAP_4325 (  );
sky130_fd_sc_hd__tap_1 TAP_4326 (  );
sky130_fd_sc_hd__tap_1 TAP_4327 (  );
sky130_fd_sc_hd__tap_1 TAP_4328 (  );
sky130_fd_sc_hd__tap_1 TAP_4329 (  );
sky130_fd_sc_hd__tap_1 TAP_4330 (  );
sky130_fd_sc_hd__tap_1 TAP_4331 (  );
sky130_fd_sc_hd__tap_1 TAP_4332 (  );
sky130_fd_sc_hd__tap_1 TAP_4333 (  );
sky130_fd_sc_hd__tap_1 TAP_4334 (  );
sky130_fd_sc_hd__tap_1 TAP_4335 (  );
sky130_fd_sc_hd__tap_1 TAP_4336 (  );
sky130_fd_sc_hd__tap_1 TAP_4337 (  );
sky130_fd_sc_hd__tap_1 TAP_4338 (  );
sky130_fd_sc_hd__tap_1 TAP_4339 (  );
sky130_fd_sc_hd__tap_1 TAP_4340 (  );
sky130_fd_sc_hd__tap_1 TAP_4341 (  );
sky130_fd_sc_hd__tap_1 TAP_4342 (  );
sky130_fd_sc_hd__tap_1 TAP_4343 (  );
sky130_fd_sc_hd__tap_1 TAP_4344 (  );
sky130_fd_sc_hd__tap_1 TAP_4345 (  );
sky130_fd_sc_hd__tap_1 TAP_4346 (  );
sky130_fd_sc_hd__tap_1 TAP_4347 (  );
sky130_fd_sc_hd__tap_1 TAP_4348 (  );
sky130_fd_sc_hd__tap_1 TAP_4349 (  );
sky130_fd_sc_hd__tap_1 TAP_4350 (  );
sky130_fd_sc_hd__tap_1 TAP_4351 (  );
sky130_fd_sc_hd__tap_1 TAP_4352 (  );
sky130_fd_sc_hd__tap_1 TAP_4353 (  );
sky130_fd_sc_hd__tap_1 TAP_4354 (  );
sky130_fd_sc_hd__tap_1 TAP_4355 (  );
sky130_fd_sc_hd__tap_1 TAP_4356 (  );
sky130_fd_sc_hd__tap_1 TAP_4357 (  );
sky130_fd_sc_hd__tap_1 TAP_4358 (  );
sky130_fd_sc_hd__tap_1 TAP_4359 (  );
sky130_fd_sc_hd__tap_1 TAP_4360 (  );
sky130_fd_sc_hd__tap_1 TAP_4361 (  );
sky130_fd_sc_hd__tap_1 TAP_4362 (  );
sky130_fd_sc_hd__tap_1 TAP_4363 (  );
sky130_fd_sc_hd__tap_1 TAP_4364 (  );
sky130_fd_sc_hd__tap_1 TAP_4365 (  );
sky130_fd_sc_hd__tap_1 TAP_4366 (  );
sky130_fd_sc_hd__tap_1 TAP_4367 (  );
sky130_fd_sc_hd__tap_1 TAP_4368 (  );
sky130_fd_sc_hd__tap_1 TAP_4369 (  );
sky130_fd_sc_hd__tap_1 TAP_4370 (  );
sky130_fd_sc_hd__tap_1 TAP_4371 (  );
sky130_fd_sc_hd__tap_1 TAP_4372 (  );
sky130_fd_sc_hd__tap_1 TAP_4373 (  );
sky130_fd_sc_hd__tap_1 TAP_4374 (  );
sky130_fd_sc_hd__tap_1 TAP_4375 (  );
sky130_fd_sc_hd__tap_1 TAP_4376 (  );
sky130_fd_sc_hd__tap_1 TAP_4377 (  );
sky130_fd_sc_hd__tap_1 TAP_4378 (  );
sky130_fd_sc_hd__tap_1 TAP_4379 (  );
sky130_fd_sc_hd__tap_1 TAP_4380 (  );
sky130_fd_sc_hd__tap_1 TAP_4381 (  );
sky130_fd_sc_hd__tap_1 TAP_4382 (  );
sky130_fd_sc_hd__tap_1 TAP_4383 (  );
sky130_fd_sc_hd__tap_1 TAP_4384 (  );
sky130_fd_sc_hd__tap_1 TAP_4385 (  );
sky130_fd_sc_hd__tap_1 TAP_4386 (  );
sky130_fd_sc_hd__tap_1 TAP_4387 (  );
sky130_fd_sc_hd__tap_1 TAP_4388 (  );
sky130_fd_sc_hd__tap_1 TAP_4389 (  );
sky130_fd_sc_hd__tap_1 TAP_4390 (  );
sky130_fd_sc_hd__tap_1 TAP_4391 (  );
sky130_fd_sc_hd__tap_1 TAP_4392 (  );
sky130_fd_sc_hd__tap_1 TAP_4393 (  );
sky130_fd_sc_hd__tap_1 TAP_4394 (  );
sky130_fd_sc_hd__tap_1 TAP_4395 (  );
sky130_fd_sc_hd__tap_1 TAP_4396 (  );
sky130_fd_sc_hd__tap_1 TAP_4397 (  );
sky130_fd_sc_hd__tap_1 TAP_4398 (  );
sky130_fd_sc_hd__tap_1 TAP_4399 (  );
sky130_fd_sc_hd__tap_1 TAP_4400 (  );
sky130_fd_sc_hd__tap_1 TAP_4401 (  );
sky130_fd_sc_hd__tap_1 TAP_4402 (  );
sky130_fd_sc_hd__tap_1 TAP_4403 (  );
sky130_fd_sc_hd__tap_1 TAP_4404 (  );
sky130_fd_sc_hd__tap_1 TAP_4405 (  );
sky130_fd_sc_hd__tap_1 TAP_4406 (  );
sky130_fd_sc_hd__tap_1 TAP_4407 (  );
sky130_fd_sc_hd__tap_1 TAP_4408 (  );
sky130_fd_sc_hd__tap_1 TAP_4409 (  );
sky130_fd_sc_hd__tap_1 TAP_4410 (  );
sky130_fd_sc_hd__tap_1 TAP_4411 (  );
sky130_fd_sc_hd__tap_1 TAP_4412 (  );
sky130_fd_sc_hd__tap_1 TAP_4413 (  );
sky130_fd_sc_hd__tap_1 TAP_4414 (  );
sky130_fd_sc_hd__tap_1 TAP_4415 (  );
sky130_fd_sc_hd__tap_1 TAP_4416 (  );
sky130_fd_sc_hd__tap_1 TAP_4417 (  );
sky130_fd_sc_hd__tap_1 TAP_4418 (  );
sky130_fd_sc_hd__tap_1 TAP_4419 (  );
sky130_fd_sc_hd__tap_1 TAP_4420 (  );
sky130_fd_sc_hd__tap_1 TAP_4421 (  );
sky130_fd_sc_hd__tap_1 TAP_4422 (  );
sky130_fd_sc_hd__tap_1 TAP_4423 (  );
sky130_fd_sc_hd__tap_1 TAP_4424 (  );
sky130_fd_sc_hd__tap_1 TAP_4425 (  );
sky130_fd_sc_hd__tap_1 TAP_4426 (  );
sky130_fd_sc_hd__tap_1 TAP_4427 (  );
sky130_fd_sc_hd__tap_1 TAP_4428 (  );
sky130_fd_sc_hd__tap_1 TAP_4429 (  );
sky130_fd_sc_hd__tap_1 TAP_4430 (  );
sky130_fd_sc_hd__tap_1 TAP_4431 (  );
sky130_fd_sc_hd__tap_1 TAP_4432 (  );
sky130_fd_sc_hd__tap_1 TAP_4433 (  );
sky130_fd_sc_hd__tap_1 TAP_4434 (  );
sky130_fd_sc_hd__tap_1 TAP_4435 (  );
sky130_fd_sc_hd__tap_1 TAP_4436 (  );
sky130_fd_sc_hd__tap_1 TAP_4437 (  );
sky130_fd_sc_hd__tap_1 TAP_4438 (  );
sky130_fd_sc_hd__tap_1 TAP_4439 (  );
sky130_fd_sc_hd__tap_1 TAP_4440 (  );
sky130_fd_sc_hd__tap_1 TAP_4441 (  );
sky130_fd_sc_hd__tap_1 TAP_4442 (  );
sky130_fd_sc_hd__tap_1 TAP_4443 (  );
sky130_fd_sc_hd__tap_1 TAP_4444 (  );
sky130_fd_sc_hd__tap_1 TAP_4445 (  );
sky130_fd_sc_hd__tap_1 TAP_4446 (  );
sky130_fd_sc_hd__tap_1 TAP_4447 (  );
sky130_fd_sc_hd__tap_1 TAP_4448 (  );
sky130_fd_sc_hd__tap_1 TAP_4449 (  );
sky130_fd_sc_hd__tap_1 TAP_4450 (  );
sky130_fd_sc_hd__tap_1 TAP_4451 (  );
sky130_fd_sc_hd__tap_1 TAP_4452 (  );
sky130_fd_sc_hd__tap_1 TAP_4453 (  );
sky130_fd_sc_hd__tap_1 TAP_4454 (  );
sky130_fd_sc_hd__tap_1 TAP_4455 (  );
sky130_fd_sc_hd__tap_1 TAP_4456 (  );
sky130_fd_sc_hd__tap_1 TAP_4457 (  );
sky130_fd_sc_hd__tap_1 TAP_4458 (  );
sky130_fd_sc_hd__tap_1 TAP_4459 (  );
sky130_fd_sc_hd__tap_1 TAP_4460 (  );
sky130_fd_sc_hd__tap_1 TAP_4461 (  );
sky130_fd_sc_hd__tap_1 TAP_4462 (  );
sky130_fd_sc_hd__tap_1 TAP_4463 (  );
sky130_fd_sc_hd__tap_1 TAP_4464 (  );
sky130_fd_sc_hd__tap_1 TAP_4465 (  );
sky130_fd_sc_hd__tap_1 TAP_4466 (  );
sky130_fd_sc_hd__tap_1 TAP_4467 (  );
sky130_fd_sc_hd__tap_1 TAP_4468 (  );
sky130_fd_sc_hd__tap_1 TAP_4469 (  );
sky130_fd_sc_hd__tap_1 TAP_4470 (  );
sky130_fd_sc_hd__tap_1 TAP_4471 (  );
sky130_fd_sc_hd__tap_1 TAP_4472 (  );
sky130_fd_sc_hd__tap_1 TAP_4473 (  );
sky130_fd_sc_hd__tap_1 TAP_4474 (  );
sky130_fd_sc_hd__tap_1 TAP_4475 (  );
sky130_fd_sc_hd__tap_1 TAP_4476 (  );
sky130_fd_sc_hd__tap_1 TAP_4477 (  );
sky130_fd_sc_hd__tap_1 TAP_4478 (  );
sky130_fd_sc_hd__tap_1 TAP_4479 (  );
sky130_fd_sc_hd__tap_1 TAP_4480 (  );
sky130_fd_sc_hd__tap_1 TAP_4481 (  );
sky130_fd_sc_hd__tap_1 TAP_4482 (  );
sky130_fd_sc_hd__tap_1 TAP_4483 (  );
sky130_fd_sc_hd__tap_1 TAP_4484 (  );
sky130_fd_sc_hd__tap_1 TAP_4485 (  );
sky130_fd_sc_hd__tap_1 TAP_4486 (  );
sky130_fd_sc_hd__tap_1 TAP_4487 (  );
sky130_fd_sc_hd__tap_1 TAP_4488 (  );
sky130_fd_sc_hd__tap_1 TAP_4489 (  );
sky130_fd_sc_hd__tap_1 TAP_4490 (  );
sky130_fd_sc_hd__tap_1 TAP_4491 (  );
sky130_fd_sc_hd__tap_1 TAP_4492 (  );
sky130_fd_sc_hd__tap_1 TAP_4493 (  );
sky130_fd_sc_hd__tap_1 TAP_4494 (  );
sky130_fd_sc_hd__tap_1 TAP_4495 (  );
sky130_fd_sc_hd__tap_1 TAP_4496 (  );
sky130_fd_sc_hd__tap_1 TAP_4497 (  );
sky130_fd_sc_hd__tap_1 TAP_4498 (  );
sky130_fd_sc_hd__tap_1 TAP_4499 (  );
sky130_fd_sc_hd__tap_1 TAP_4500 (  );
sky130_fd_sc_hd__tap_1 TAP_4501 (  );
sky130_fd_sc_hd__tap_1 TAP_4502 (  );
sky130_fd_sc_hd__tap_1 TAP_4503 (  );
sky130_fd_sc_hd__tap_1 TAP_4504 (  );
sky130_fd_sc_hd__tap_1 TAP_4505 (  );
sky130_fd_sc_hd__tap_1 TAP_4506 (  );
sky130_fd_sc_hd__tap_1 TAP_4507 (  );
sky130_fd_sc_hd__tap_1 TAP_4508 (  );
sky130_fd_sc_hd__tap_1 TAP_4509 (  );
sky130_fd_sc_hd__tap_1 TAP_4510 (  );
sky130_fd_sc_hd__tap_1 TAP_4511 (  );
sky130_fd_sc_hd__tap_1 TAP_4512 (  );
sky130_fd_sc_hd__tap_1 TAP_4513 (  );
sky130_fd_sc_hd__tap_1 TAP_4514 (  );
sky130_fd_sc_hd__tap_1 TAP_4515 (  );
sky130_fd_sc_hd__tap_1 TAP_4516 (  );
sky130_fd_sc_hd__tap_1 TAP_4517 (  );
sky130_fd_sc_hd__tap_1 TAP_4518 (  );
sky130_fd_sc_hd__tap_1 TAP_4519 (  );
sky130_fd_sc_hd__tap_1 TAP_4520 (  );
sky130_fd_sc_hd__tap_1 TAP_4521 (  );
sky130_fd_sc_hd__tap_1 TAP_4522 (  );
sky130_fd_sc_hd__tap_1 TAP_4523 (  );
sky130_fd_sc_hd__tap_1 TAP_4524 (  );
sky130_fd_sc_hd__tap_1 TAP_4525 (  );
sky130_fd_sc_hd__tap_1 TAP_4526 (  );
sky130_fd_sc_hd__tap_1 TAP_4527 (  );
sky130_fd_sc_hd__tap_1 TAP_4528 (  );
sky130_fd_sc_hd__tap_1 TAP_4529 (  );
sky130_fd_sc_hd__tap_1 TAP_4530 (  );
sky130_fd_sc_hd__tap_1 TAP_4531 (  );
sky130_fd_sc_hd__tap_1 TAP_4532 (  );
sky130_fd_sc_hd__tap_1 TAP_4533 (  );
sky130_fd_sc_hd__tap_1 TAP_4534 (  );
sky130_fd_sc_hd__tap_1 TAP_4535 (  );
sky130_fd_sc_hd__tap_1 TAP_4536 (  );
sky130_fd_sc_hd__tap_1 TAP_4537 (  );
sky130_fd_sc_hd__tap_1 TAP_4538 (  );
sky130_fd_sc_hd__tap_1 TAP_4539 (  );
sky130_fd_sc_hd__tap_1 TAP_4540 (  );
sky130_fd_sc_hd__tap_1 TAP_4541 (  );
sky130_fd_sc_hd__tap_1 TAP_4542 (  );
sky130_fd_sc_hd__tap_1 TAP_4543 (  );
sky130_fd_sc_hd__tap_1 TAP_4544 (  );
sky130_fd_sc_hd__tap_1 TAP_4545 (  );
sky130_fd_sc_hd__tap_1 TAP_4546 (  );
sky130_fd_sc_hd__tap_1 TAP_4547 (  );
sky130_fd_sc_hd__tap_1 TAP_4548 (  );
sky130_fd_sc_hd__tap_1 TAP_4549 (  );
sky130_fd_sc_hd__tap_1 TAP_4550 (  );
sky130_fd_sc_hd__tap_1 TAP_4551 (  );
sky130_fd_sc_hd__tap_1 TAP_4552 (  );
sky130_fd_sc_hd__tap_1 TAP_4553 (  );
sky130_fd_sc_hd__tap_1 TAP_4554 (  );
sky130_fd_sc_hd__tap_1 TAP_4555 (  );
sky130_fd_sc_hd__tap_1 TAP_4556 (  );
sky130_fd_sc_hd__tap_1 TAP_4557 (  );
sky130_fd_sc_hd__tap_1 TAP_4558 (  );
sky130_fd_sc_hd__tap_1 TAP_4559 (  );
sky130_fd_sc_hd__tap_1 TAP_4560 (  );
sky130_fd_sc_hd__tap_1 TAP_4561 (  );
sky130_fd_sc_hd__tap_1 TAP_4562 (  );
sky130_fd_sc_hd__tap_1 TAP_4563 (  );
sky130_fd_sc_hd__tap_1 TAP_4564 (  );
sky130_fd_sc_hd__tap_1 TAP_4565 (  );
sky130_fd_sc_hd__tap_1 TAP_4566 (  );
sky130_fd_sc_hd__tap_1 TAP_4567 (  );
sky130_fd_sc_hd__tap_1 TAP_4568 (  );
sky130_fd_sc_hd__tap_1 TAP_4569 (  );
sky130_fd_sc_hd__tap_1 TAP_4570 (  );
sky130_fd_sc_hd__tap_1 TAP_4571 (  );
sky130_fd_sc_hd__tap_1 TAP_4572 (  );
sky130_fd_sc_hd__tap_1 TAP_4573 (  );
sky130_fd_sc_hd__tap_1 TAP_4574 (  );
sky130_fd_sc_hd__tap_1 TAP_4575 (  );
sky130_fd_sc_hd__tap_1 TAP_4576 (  );
sky130_fd_sc_hd__tap_1 TAP_4577 (  );
sky130_fd_sc_hd__tap_1 TAP_4578 (  );
sky130_fd_sc_hd__tap_1 TAP_4579 (  );
sky130_fd_sc_hd__tap_1 TAP_4580 (  );
sky130_fd_sc_hd__tap_1 TAP_4581 (  );
sky130_fd_sc_hd__tap_1 TAP_4582 (  );
sky130_fd_sc_hd__tap_1 TAP_4583 (  );
sky130_fd_sc_hd__tap_1 TAP_4584 (  );
sky130_fd_sc_hd__tap_1 TAP_4585 (  );
sky130_fd_sc_hd__tap_1 TAP_4586 (  );
sky130_fd_sc_hd__tap_1 TAP_4587 (  );
sky130_fd_sc_hd__tap_1 TAP_4588 (  );
sky130_fd_sc_hd__tap_1 TAP_4589 (  );
sky130_fd_sc_hd__tap_1 TAP_4590 (  );
sky130_fd_sc_hd__tap_1 TAP_4591 (  );
sky130_fd_sc_hd__tap_1 TAP_4592 (  );
sky130_fd_sc_hd__tap_1 TAP_4593 (  );
sky130_fd_sc_hd__tap_1 TAP_4594 (  );
sky130_fd_sc_hd__tap_1 TAP_4595 (  );
sky130_fd_sc_hd__tap_1 TAP_4596 (  );
sky130_fd_sc_hd__tap_1 TAP_4597 (  );
sky130_fd_sc_hd__tap_1 TAP_4598 (  );
sky130_fd_sc_hd__tap_1 TAP_4599 (  );
sky130_fd_sc_hd__tap_1 TAP_4600 (  );
sky130_fd_sc_hd__tap_1 TAP_4601 (  );
sky130_fd_sc_hd__tap_1 TAP_4602 (  );
sky130_fd_sc_hd__tap_1 TAP_4603 (  );
sky130_fd_sc_hd__tap_1 TAP_4604 (  );
sky130_fd_sc_hd__tap_1 TAP_4605 (  );
sky130_fd_sc_hd__tap_1 TAP_4606 (  );
sky130_fd_sc_hd__tap_1 TAP_4607 (  );
sky130_fd_sc_hd__tap_1 TAP_4608 (  );
sky130_fd_sc_hd__tap_1 TAP_4609 (  );
sky130_fd_sc_hd__tap_1 TAP_4610 (  );
sky130_fd_sc_hd__tap_1 TAP_4611 (  );
sky130_fd_sc_hd__tap_1 TAP_4612 (  );
sky130_fd_sc_hd__tap_1 TAP_4613 (  );
sky130_fd_sc_hd__tap_1 TAP_4614 (  );
sky130_fd_sc_hd__tap_1 TAP_4615 (  );
sky130_fd_sc_hd__tap_1 TAP_4616 (  );
sky130_fd_sc_hd__tap_1 TAP_4617 (  );
sky130_fd_sc_hd__tap_1 TAP_4618 (  );
sky130_fd_sc_hd__tap_1 TAP_4619 (  );
sky130_fd_sc_hd__tap_1 TAP_4620 (  );
sky130_fd_sc_hd__tap_1 TAP_4621 (  );
sky130_fd_sc_hd__tap_1 TAP_4622 (  );
sky130_fd_sc_hd__tap_1 TAP_4623 (  );
sky130_fd_sc_hd__tap_1 TAP_4624 (  );
sky130_fd_sc_hd__tap_1 TAP_4625 (  );
sky130_fd_sc_hd__tap_1 TAP_4626 (  );
sky130_fd_sc_hd__tap_1 TAP_4627 (  );
sky130_fd_sc_hd__tap_1 TAP_4628 (  );
sky130_fd_sc_hd__tap_1 TAP_4629 (  );
sky130_fd_sc_hd__tap_1 TAP_4630 (  );
sky130_fd_sc_hd__tap_1 TAP_4631 (  );
sky130_fd_sc_hd__tap_1 TAP_4632 (  );
sky130_fd_sc_hd__tap_1 TAP_4633 (  );
sky130_fd_sc_hd__tap_1 TAP_4634 (  );
sky130_fd_sc_hd__tap_1 TAP_4635 (  );
sky130_fd_sc_hd__tap_1 TAP_4636 (  );
sky130_fd_sc_hd__tap_1 TAP_4637 (  );
sky130_fd_sc_hd__tap_1 TAP_4638 (  );
sky130_fd_sc_hd__tap_1 TAP_4639 (  );
sky130_fd_sc_hd__tap_1 TAP_4640 (  );
sky130_fd_sc_hd__tap_1 TAP_4641 (  );
sky130_fd_sc_hd__tap_1 TAP_4642 (  );
sky130_fd_sc_hd__tap_1 TAP_4643 (  );
sky130_fd_sc_hd__tap_1 TAP_4644 (  );
sky130_fd_sc_hd__tap_1 TAP_4645 (  );
sky130_fd_sc_hd__tap_1 TAP_4646 (  );
sky130_fd_sc_hd__tap_1 TAP_4647 (  );
sky130_fd_sc_hd__tap_1 TAP_4648 (  );
sky130_fd_sc_hd__tap_1 TAP_4649 (  );
sky130_fd_sc_hd__tap_1 TAP_4650 (  );
sky130_fd_sc_hd__tap_1 TAP_4651 (  );
sky130_fd_sc_hd__tap_1 TAP_4652 (  );
sky130_fd_sc_hd__tap_1 TAP_4653 (  );
sky130_fd_sc_hd__tap_1 TAP_4654 (  );
sky130_fd_sc_hd__tap_1 TAP_4655 (  );
sky130_fd_sc_hd__tap_1 TAP_4656 (  );
sky130_fd_sc_hd__tap_1 TAP_4657 (  );
sky130_fd_sc_hd__tap_1 TAP_4658 (  );
sky130_fd_sc_hd__tap_1 TAP_4659 (  );
sky130_fd_sc_hd__tap_1 TAP_4660 (  );
sky130_fd_sc_hd__tap_1 TAP_4661 (  );
sky130_fd_sc_hd__tap_1 TAP_4662 (  );
sky130_fd_sc_hd__tap_1 TAP_4663 (  );
sky130_fd_sc_hd__tap_1 TAP_4664 (  );
sky130_fd_sc_hd__tap_1 TAP_4665 (  );
sky130_fd_sc_hd__tap_1 TAP_4666 (  );
sky130_fd_sc_hd__tap_1 TAP_4667 (  );
sky130_fd_sc_hd__tap_1 TAP_4668 (  );
sky130_fd_sc_hd__tap_1 TAP_4669 (  );
sky130_fd_sc_hd__tap_1 TAP_4670 (  );
sky130_fd_sc_hd__tap_1 TAP_4671 (  );
sky130_fd_sc_hd__tap_1 TAP_4672 (  );
sky130_fd_sc_hd__tap_1 TAP_4673 (  );
sky130_fd_sc_hd__tap_1 TAP_4674 (  );
sky130_fd_sc_hd__tap_1 TAP_4675 (  );
sky130_fd_sc_hd__tap_1 TAP_4676 (  );
sky130_fd_sc_hd__tap_1 TAP_4677 (  );
sky130_fd_sc_hd__tap_1 TAP_4678 (  );
sky130_fd_sc_hd__tap_1 TAP_4679 (  );
sky130_fd_sc_hd__tap_1 TAP_4680 (  );
sky130_fd_sc_hd__tap_1 TAP_4681 (  );
sky130_fd_sc_hd__tap_1 TAP_4682 (  );
sky130_fd_sc_hd__tap_1 TAP_4683 (  );
sky130_fd_sc_hd__tap_1 TAP_4684 (  );
sky130_fd_sc_hd__tap_1 TAP_4685 (  );
sky130_fd_sc_hd__tap_1 TAP_4686 (  );
sky130_fd_sc_hd__tap_1 TAP_4687 (  );
sky130_fd_sc_hd__tap_1 TAP_4688 (  );
sky130_fd_sc_hd__tap_1 TAP_4689 (  );
sky130_fd_sc_hd__tap_1 TAP_4690 (  );
sky130_fd_sc_hd__tap_1 TAP_4691 (  );
sky130_fd_sc_hd__tap_1 TAP_4692 (  );
sky130_fd_sc_hd__tap_1 TAP_4693 (  );
sky130_fd_sc_hd__tap_1 TAP_4694 (  );
sky130_fd_sc_hd__tap_1 TAP_4695 (  );
sky130_fd_sc_hd__tap_1 TAP_4696 (  );
sky130_fd_sc_hd__tap_1 TAP_4697 (  );
sky130_fd_sc_hd__tap_1 TAP_4698 (  );
sky130_fd_sc_hd__tap_1 TAP_4699 (  );
sky130_fd_sc_hd__tap_1 TAP_4700 (  );
sky130_fd_sc_hd__tap_1 TAP_4701 (  );
sky130_fd_sc_hd__tap_1 TAP_4702 (  );
sky130_fd_sc_hd__tap_1 TAP_4703 (  );
sky130_fd_sc_hd__tap_1 TAP_4704 (  );
sky130_fd_sc_hd__tap_1 TAP_4705 (  );
sky130_fd_sc_hd__tap_1 TAP_4706 (  );
sky130_fd_sc_hd__tap_1 TAP_4707 (  );
sky130_fd_sc_hd__tap_1 TAP_4708 (  );
sky130_fd_sc_hd__tap_1 TAP_4709 (  );
sky130_fd_sc_hd__tap_1 TAP_4710 (  );
sky130_fd_sc_hd__tap_1 TAP_4711 (  );
sky130_fd_sc_hd__tap_1 TAP_4712 (  );
sky130_fd_sc_hd__tap_1 TAP_4713 (  );
sky130_fd_sc_hd__tap_1 TAP_4714 (  );
sky130_fd_sc_hd__tap_1 TAP_4715 (  );
sky130_fd_sc_hd__tap_1 TAP_4716 (  );
sky130_fd_sc_hd__tap_1 TAP_4717 (  );
sky130_fd_sc_hd__tap_1 TAP_4718 (  );
sky130_fd_sc_hd__tap_1 TAP_4719 (  );
sky130_fd_sc_hd__tap_1 TAP_4720 (  );
sky130_fd_sc_hd__tap_1 TAP_4721 (  );
sky130_fd_sc_hd__tap_1 TAP_4722 (  );
sky130_fd_sc_hd__tap_1 TAP_4723 (  );
sky130_fd_sc_hd__tap_1 TAP_4724 (  );
sky130_fd_sc_hd__tap_1 TAP_4725 (  );
sky130_fd_sc_hd__tap_1 TAP_4726 (  );
sky130_fd_sc_hd__tap_1 TAP_4727 (  );
sky130_fd_sc_hd__tap_1 TAP_4728 (  );
sky130_fd_sc_hd__tap_1 TAP_4729 (  );
sky130_fd_sc_hd__tap_1 TAP_4730 (  );
sky130_fd_sc_hd__tap_1 TAP_4731 (  );
sky130_fd_sc_hd__tap_1 TAP_4732 (  );
sky130_fd_sc_hd__tap_1 TAP_4733 (  );
sky130_fd_sc_hd__tap_1 TAP_4734 (  );
sky130_fd_sc_hd__tap_1 TAP_4735 (  );
sky130_fd_sc_hd__tap_1 TAP_4736 (  );
sky130_fd_sc_hd__tap_1 TAP_4737 (  );
sky130_fd_sc_hd__tap_1 TAP_4738 (  );
sky130_fd_sc_hd__tap_1 TAP_4739 (  );
sky130_fd_sc_hd__tap_1 TAP_4740 (  );
sky130_fd_sc_hd__tap_1 TAP_4741 (  );
sky130_fd_sc_hd__tap_1 TAP_4742 (  );
sky130_fd_sc_hd__tap_1 TAP_4743 (  );
sky130_fd_sc_hd__tap_1 TAP_4744 (  );
sky130_fd_sc_hd__tap_1 TAP_4745 (  );
sky130_fd_sc_hd__tap_1 TAP_4746 (  );
sky130_fd_sc_hd__tap_1 TAP_4747 (  );
sky130_fd_sc_hd__tap_1 TAP_4748 (  );
sky130_fd_sc_hd__tap_1 TAP_4749 (  );
sky130_fd_sc_hd__tap_1 TAP_4750 (  );
sky130_fd_sc_hd__tap_1 TAP_4751 (  );
sky130_fd_sc_hd__tap_1 TAP_4752 (  );
sky130_fd_sc_hd__tap_1 TAP_4753 (  );
sky130_fd_sc_hd__tap_1 TAP_4754 (  );
sky130_fd_sc_hd__tap_1 TAP_4755 (  );
sky130_fd_sc_hd__tap_1 TAP_4756 (  );
sky130_fd_sc_hd__tap_1 TAP_4757 (  );
sky130_fd_sc_hd__tap_1 TAP_4758 (  );
sky130_fd_sc_hd__tap_1 TAP_4759 (  );
sky130_fd_sc_hd__tap_1 TAP_4760 (  );
sky130_fd_sc_hd__tap_1 TAP_4761 (  );
sky130_fd_sc_hd__tap_1 TAP_4762 (  );
sky130_fd_sc_hd__tap_1 TAP_4763 (  );
sky130_fd_sc_hd__tap_1 TAP_4764 (  );
sky130_fd_sc_hd__tap_1 TAP_4765 (  );
sky130_fd_sc_hd__tap_1 TAP_4766 (  );
sky130_fd_sc_hd__tap_1 TAP_4767 (  );
sky130_fd_sc_hd__tap_1 TAP_4768 (  );
sky130_fd_sc_hd__tap_1 TAP_4769 (  );
sky130_fd_sc_hd__tap_1 TAP_4770 (  );
sky130_fd_sc_hd__tap_1 TAP_4771 (  );
sky130_fd_sc_hd__tap_1 TAP_4772 (  );
sky130_fd_sc_hd__tap_1 TAP_4773 (  );
sky130_fd_sc_hd__tap_1 TAP_4774 (  );
sky130_fd_sc_hd__tap_1 TAP_4775 (  );
sky130_fd_sc_hd__tap_1 TAP_4776 (  );
sky130_fd_sc_hd__tap_1 TAP_4777 (  );
sky130_fd_sc_hd__tap_1 TAP_4778 (  );
sky130_fd_sc_hd__tap_1 TAP_4779 (  );
sky130_fd_sc_hd__tap_1 TAP_4780 (  );
sky130_fd_sc_hd__tap_1 TAP_4781 (  );
sky130_fd_sc_hd__tap_1 TAP_4782 (  );
sky130_fd_sc_hd__tap_1 TAP_4783 (  );
sky130_fd_sc_hd__tap_1 TAP_4784 (  );
sky130_fd_sc_hd__tap_1 TAP_4785 (  );
sky130_fd_sc_hd__tap_1 TAP_4786 (  );
sky130_fd_sc_hd__tap_1 TAP_4787 (  );
sky130_fd_sc_hd__tap_1 TAP_4788 (  );
sky130_fd_sc_hd__tap_1 TAP_4789 (  );
sky130_fd_sc_hd__tap_1 TAP_4790 (  );
sky130_fd_sc_hd__tap_1 TAP_4791 (  );
sky130_fd_sc_hd__tap_1 TAP_4792 (  );
sky130_fd_sc_hd__tap_1 TAP_4793 (  );
sky130_fd_sc_hd__tap_1 TAP_4794 (  );
sky130_fd_sc_hd__tap_1 TAP_4795 (  );
sky130_fd_sc_hd__tap_1 TAP_4796 (  );
sky130_fd_sc_hd__tap_1 TAP_4797 (  );
sky130_fd_sc_hd__tap_1 TAP_4798 (  );
sky130_fd_sc_hd__tap_1 TAP_4799 (  );
sky130_fd_sc_hd__tap_1 TAP_4800 (  );
sky130_fd_sc_hd__tap_1 TAP_4801 (  );
sky130_fd_sc_hd__tap_1 TAP_4802 (  );
sky130_fd_sc_hd__tap_1 TAP_4803 (  );
sky130_fd_sc_hd__tap_1 TAP_4804 (  );
sky130_fd_sc_hd__tap_1 TAP_4805 (  );
sky130_fd_sc_hd__tap_1 TAP_4806 (  );
sky130_fd_sc_hd__tap_1 TAP_4807 (  );
sky130_fd_sc_hd__tap_1 TAP_4808 (  );
sky130_fd_sc_hd__tap_1 TAP_4809 (  );
sky130_fd_sc_hd__tap_1 TAP_4810 (  );
sky130_fd_sc_hd__tap_1 TAP_4811 (  );
sky130_fd_sc_hd__tap_1 TAP_4812 (  );
sky130_fd_sc_hd__tap_1 TAP_4813 (  );
sky130_fd_sc_hd__tap_1 TAP_4814 (  );
sky130_fd_sc_hd__tap_1 TAP_4815 (  );
sky130_fd_sc_hd__tap_1 TAP_4816 (  );
sky130_fd_sc_hd__tap_1 TAP_4817 (  );
sky130_fd_sc_hd__tap_1 TAP_4818 (  );
sky130_fd_sc_hd__tap_1 TAP_4819 (  );
sky130_fd_sc_hd__tap_1 TAP_4820 (  );
sky130_fd_sc_hd__tap_1 TAP_4821 (  );
sky130_fd_sc_hd__tap_1 TAP_4822 (  );
sky130_fd_sc_hd__tap_1 TAP_4823 (  );
sky130_fd_sc_hd__tap_1 TAP_4824 (  );
sky130_fd_sc_hd__tap_1 TAP_4825 (  );
sky130_fd_sc_hd__tap_1 TAP_4826 (  );
sky130_fd_sc_hd__tap_1 TAP_4827 (  );
sky130_fd_sc_hd__tap_1 TAP_4828 (  );
sky130_fd_sc_hd__tap_1 TAP_4829 (  );
sky130_fd_sc_hd__tap_1 TAP_4830 (  );
sky130_fd_sc_hd__tap_1 TAP_4831 (  );
sky130_fd_sc_hd__tap_1 TAP_4832 (  );
sky130_fd_sc_hd__tap_1 TAP_4833 (  );
sky130_fd_sc_hd__tap_1 TAP_4834 (  );
sky130_fd_sc_hd__tap_1 TAP_4835 (  );
sky130_fd_sc_hd__tap_1 TAP_4836 (  );
sky130_fd_sc_hd__tap_1 TAP_4837 (  );
sky130_fd_sc_hd__tap_1 TAP_4838 (  );
sky130_fd_sc_hd__tap_1 TAP_4839 (  );
sky130_fd_sc_hd__tap_1 TAP_4840 (  );
sky130_fd_sc_hd__tap_1 TAP_4841 (  );
sky130_fd_sc_hd__tap_1 TAP_4842 (  );
sky130_fd_sc_hd__tap_1 TAP_4843 (  );
sky130_fd_sc_hd__tap_1 TAP_4844 (  );
sky130_fd_sc_hd__tap_1 TAP_4845 (  );
sky130_fd_sc_hd__tap_1 TAP_4846 (  );
sky130_fd_sc_hd__tap_1 TAP_4847 (  );
sky130_fd_sc_hd__tap_1 TAP_4848 (  );
sky130_fd_sc_hd__tap_1 TAP_4849 (  );
sky130_fd_sc_hd__tap_1 TAP_4850 (  );
sky130_fd_sc_hd__tap_1 TAP_4851 (  );
sky130_fd_sc_hd__tap_1 TAP_4852 (  );
sky130_fd_sc_hd__tap_1 TAP_4853 (  );
sky130_fd_sc_hd__tap_1 TAP_4854 (  );
sky130_fd_sc_hd__tap_1 TAP_4855 (  );
sky130_fd_sc_hd__tap_1 TAP_4856 (  );
sky130_fd_sc_hd__tap_1 TAP_4857 (  );
sky130_fd_sc_hd__tap_1 TAP_4858 (  );
sky130_fd_sc_hd__tap_1 TAP_4859 (  );
sky130_fd_sc_hd__tap_1 TAP_4860 (  );
sky130_fd_sc_hd__tap_1 TAP_4861 (  );
sky130_fd_sc_hd__tap_1 TAP_4862 (  );
sky130_fd_sc_hd__tap_1 TAP_4863 (  );
sky130_fd_sc_hd__tap_1 TAP_4864 (  );
sky130_fd_sc_hd__tap_1 TAP_4865 (  );
sky130_fd_sc_hd__tap_1 TAP_4866 (  );
sky130_fd_sc_hd__tap_1 TAP_4867 (  );
sky130_fd_sc_hd__tap_1 TAP_4868 (  );
sky130_fd_sc_hd__tap_1 TAP_4869 (  );
sky130_fd_sc_hd__tap_1 TAP_4870 (  );
sky130_fd_sc_hd__tap_1 TAP_4871 (  );
sky130_fd_sc_hd__tap_1 TAP_4872 (  );
sky130_fd_sc_hd__tap_1 TAP_4873 (  );
sky130_fd_sc_hd__tap_1 TAP_4874 (  );
sky130_fd_sc_hd__tap_1 TAP_4875 (  );
sky130_fd_sc_hd__tap_1 TAP_4876 (  );
sky130_fd_sc_hd__tap_1 TAP_4877 (  );
sky130_fd_sc_hd__tap_1 TAP_4878 (  );
sky130_fd_sc_hd__tap_1 TAP_4879 (  );
sky130_fd_sc_hd__tap_1 TAP_4880 (  );
sky130_fd_sc_hd__tap_1 TAP_4881 (  );
sky130_fd_sc_hd__tap_1 TAP_4882 (  );
sky130_fd_sc_hd__tap_1 TAP_4883 (  );
sky130_fd_sc_hd__tap_1 TAP_4884 (  );
sky130_fd_sc_hd__tap_1 TAP_4885 (  );
sky130_fd_sc_hd__tap_1 TAP_4886 (  );
sky130_fd_sc_hd__tap_1 TAP_4887 (  );
sky130_fd_sc_hd__tap_1 TAP_4888 (  );
sky130_fd_sc_hd__tap_1 TAP_4889 (  );
sky130_fd_sc_hd__tap_1 TAP_4890 (  );
sky130_fd_sc_hd__tap_1 TAP_4891 (  );
sky130_fd_sc_hd__tap_1 TAP_4892 (  );
sky130_fd_sc_hd__tap_1 TAP_4893 (  );
sky130_fd_sc_hd__tap_1 TAP_4894 (  );
sky130_fd_sc_hd__tap_1 TAP_4895 (  );
sky130_fd_sc_hd__tap_1 TAP_4896 (  );
sky130_fd_sc_hd__tap_1 TAP_4897 (  );
sky130_fd_sc_hd__tap_1 TAP_4898 (  );
sky130_fd_sc_hd__tap_1 TAP_4899 (  );
sky130_fd_sc_hd__tap_1 TAP_4900 (  );
sky130_fd_sc_hd__tap_1 TAP_4901 (  );
sky130_fd_sc_hd__tap_1 TAP_4902 (  );
sky130_fd_sc_hd__tap_1 TAP_4903 (  );
sky130_fd_sc_hd__tap_1 TAP_4904 (  );
sky130_fd_sc_hd__tap_1 TAP_4905 (  );
sky130_fd_sc_hd__tap_1 TAP_4906 (  );
sky130_fd_sc_hd__tap_1 TAP_4907 (  );
sky130_fd_sc_hd__tap_1 TAP_4908 (  );
sky130_fd_sc_hd__tap_1 TAP_4909 (  );
sky130_fd_sc_hd__tap_1 TAP_4910 (  );
sky130_fd_sc_hd__tap_1 TAP_4911 (  );
sky130_fd_sc_hd__tap_1 TAP_4912 (  );
sky130_fd_sc_hd__tap_1 TAP_4913 (  );
sky130_fd_sc_hd__tap_1 TAP_4914 (  );
sky130_fd_sc_hd__tap_1 TAP_4915 (  );
sky130_fd_sc_hd__tap_1 TAP_4916 (  );
sky130_fd_sc_hd__tap_1 TAP_4917 (  );
sky130_fd_sc_hd__tap_1 TAP_4918 (  );
sky130_fd_sc_hd__tap_1 TAP_4919 (  );
sky130_fd_sc_hd__tap_1 TAP_4920 (  );
sky130_fd_sc_hd__tap_1 TAP_4921 (  );
sky130_fd_sc_hd__tap_1 TAP_4922 (  );
sky130_fd_sc_hd__tap_1 TAP_4923 (  );
sky130_fd_sc_hd__tap_1 TAP_4924 (  );
sky130_fd_sc_hd__tap_1 TAP_4925 (  );
sky130_fd_sc_hd__tap_1 TAP_4926 (  );
sky130_fd_sc_hd__tap_1 TAP_4927 (  );
sky130_fd_sc_hd__tap_1 TAP_4928 (  );
sky130_fd_sc_hd__tap_1 TAP_4929 (  );
sky130_fd_sc_hd__tap_1 TAP_4930 (  );
sky130_fd_sc_hd__tap_1 TAP_4931 (  );
sky130_fd_sc_hd__tap_1 TAP_4932 (  );
sky130_fd_sc_hd__tap_1 TAP_4933 (  );
sky130_fd_sc_hd__tap_1 TAP_4934 (  );
sky130_fd_sc_hd__tap_1 TAP_4935 (  );
sky130_fd_sc_hd__tap_1 TAP_4936 (  );
sky130_fd_sc_hd__tap_1 TAP_4937 (  );
sky130_fd_sc_hd__tap_1 TAP_4938 (  );
sky130_fd_sc_hd__tap_1 TAP_4939 (  );
sky130_fd_sc_hd__tap_1 TAP_4940 (  );
sky130_fd_sc_hd__tap_1 TAP_4941 (  );
sky130_fd_sc_hd__tap_1 TAP_4942 (  );
sky130_fd_sc_hd__tap_1 TAP_4943 (  );
sky130_fd_sc_hd__tap_1 TAP_4944 (  );
sky130_fd_sc_hd__tap_1 TAP_4945 (  );
sky130_fd_sc_hd__tap_1 TAP_4946 (  );
sky130_fd_sc_hd__tap_1 TAP_4947 (  );
sky130_fd_sc_hd__tap_1 TAP_4948 (  );
sky130_fd_sc_hd__tap_1 TAP_4949 (  );
sky130_fd_sc_hd__tap_1 TAP_4950 (  );
sky130_fd_sc_hd__tap_1 TAP_4951 (  );
sky130_fd_sc_hd__tap_1 TAP_4952 (  );
sky130_fd_sc_hd__tap_1 TAP_4953 (  );
sky130_fd_sc_hd__tap_1 TAP_4954 (  );
sky130_fd_sc_hd__tap_1 TAP_4955 (  );
sky130_fd_sc_hd__tap_1 TAP_4956 (  );
sky130_fd_sc_hd__tap_1 TAP_4957 (  );
sky130_fd_sc_hd__tap_1 TAP_4958 (  );
sky130_fd_sc_hd__tap_1 TAP_4959 (  );
sky130_fd_sc_hd__tap_1 TAP_4960 (  );
sky130_fd_sc_hd__tap_1 TAP_4961 (  );
sky130_fd_sc_hd__tap_1 TAP_4962 (  );
sky130_fd_sc_hd__tap_1 TAP_4963 (  );
sky130_fd_sc_hd__tap_1 TAP_4964 (  );
sky130_fd_sc_hd__tap_1 TAP_4965 (  );
sky130_fd_sc_hd__tap_1 TAP_4966 (  );
sky130_fd_sc_hd__tap_1 TAP_4967 (  );
sky130_fd_sc_hd__tap_1 TAP_4968 (  );
sky130_fd_sc_hd__tap_1 TAP_4969 (  );
sky130_fd_sc_hd__tap_1 TAP_4970 (  );
sky130_fd_sc_hd__tap_1 TAP_4971 (  );
sky130_fd_sc_hd__tap_1 TAP_4972 (  );
sky130_fd_sc_hd__tap_1 TAP_4973 (  );
sky130_fd_sc_hd__tap_1 TAP_4974 (  );
sky130_fd_sc_hd__tap_1 TAP_4975 (  );
sky130_fd_sc_hd__tap_1 TAP_4976 (  );
sky130_fd_sc_hd__tap_1 TAP_4977 (  );
sky130_fd_sc_hd__tap_1 TAP_4978 (  );
sky130_fd_sc_hd__tap_1 TAP_4979 (  );
sky130_fd_sc_hd__tap_1 TAP_4980 (  );
sky130_fd_sc_hd__tap_1 TAP_4981 (  );
sky130_fd_sc_hd__tap_1 TAP_4982 (  );
sky130_fd_sc_hd__tap_1 TAP_4983 (  );
sky130_fd_sc_hd__tap_1 TAP_4984 (  );
sky130_fd_sc_hd__tap_1 TAP_4985 (  );
sky130_fd_sc_hd__tap_1 TAP_4986 (  );
sky130_fd_sc_hd__tap_1 TAP_4987 (  );
sky130_fd_sc_hd__tap_1 TAP_4988 (  );
sky130_fd_sc_hd__tap_1 TAP_4989 (  );
sky130_fd_sc_hd__tap_1 TAP_4990 (  );
sky130_fd_sc_hd__tap_1 TAP_4991 (  );
sky130_fd_sc_hd__tap_1 TAP_4992 (  );
sky130_fd_sc_hd__tap_1 TAP_4993 (  );
sky130_fd_sc_hd__tap_1 TAP_4994 (  );
sky130_fd_sc_hd__tap_1 TAP_4995 (  );
sky130_fd_sc_hd__tap_1 TAP_4996 (  );
sky130_fd_sc_hd__tap_1 TAP_4997 (  );
sky130_fd_sc_hd__tap_1 TAP_4998 (  );
sky130_fd_sc_hd__tap_1 TAP_4999 (  );
sky130_fd_sc_hd__tap_1 TAP_5000 (  );
sky130_fd_sc_hd__tap_1 TAP_5001 (  );
sky130_fd_sc_hd__tap_1 TAP_5002 (  );
sky130_fd_sc_hd__tap_1 TAP_5003 (  );
sky130_fd_sc_hd__tap_1 TAP_5004 (  );
sky130_fd_sc_hd__tap_1 TAP_5005 (  );
sky130_fd_sc_hd__tap_1 TAP_5006 (  );
sky130_fd_sc_hd__tap_1 TAP_5007 (  );
sky130_fd_sc_hd__tap_1 TAP_5008 (  );
sky130_fd_sc_hd__tap_1 TAP_5009 (  );
sky130_fd_sc_hd__tap_1 TAP_5010 (  );
sky130_fd_sc_hd__tap_1 TAP_5011 (  );
sky130_fd_sc_hd__tap_1 TAP_5012 (  );
sky130_fd_sc_hd__tap_1 TAP_5013 (  );
sky130_fd_sc_hd__tap_1 TAP_5014 (  );
sky130_fd_sc_hd__tap_1 TAP_5015 (  );
sky130_fd_sc_hd__tap_1 TAP_5016 (  );
sky130_fd_sc_hd__tap_1 TAP_5017 (  );
sky130_fd_sc_hd__tap_1 TAP_5018 (  );
sky130_fd_sc_hd__tap_1 TAP_5019 (  );
sky130_fd_sc_hd__tap_1 TAP_5020 (  );
sky130_fd_sc_hd__tap_1 TAP_5021 (  );
sky130_fd_sc_hd__tap_1 TAP_5022 (  );
sky130_fd_sc_hd__tap_1 TAP_5023 (  );
sky130_fd_sc_hd__tap_1 TAP_5024 (  );
sky130_fd_sc_hd__tap_1 TAP_5025 (  );
sky130_fd_sc_hd__tap_1 TAP_5026 (  );
sky130_fd_sc_hd__tap_1 TAP_5027 (  );
sky130_fd_sc_hd__tap_1 TAP_5028 (  );
sky130_fd_sc_hd__tap_1 TAP_5029 (  );
sky130_fd_sc_hd__tap_1 TAP_5030 (  );
sky130_fd_sc_hd__tap_1 TAP_5031 (  );
sky130_fd_sc_hd__tap_1 TAP_5032 (  );
sky130_fd_sc_hd__tap_1 TAP_5033 (  );
sky130_fd_sc_hd__tap_1 TAP_5034 (  );
sky130_fd_sc_hd__tap_1 TAP_5035 (  );
sky130_fd_sc_hd__tap_1 TAP_5036 (  );
sky130_fd_sc_hd__tap_1 TAP_5037 (  );
sky130_fd_sc_hd__tap_1 TAP_5038 (  );
sky130_fd_sc_hd__tap_1 TAP_5039 (  );
sky130_fd_sc_hd__tap_1 TAP_5040 (  );
sky130_fd_sc_hd__tap_1 TAP_5041 (  );
sky130_fd_sc_hd__tap_1 TAP_5042 (  );
sky130_fd_sc_hd__tap_1 TAP_5043 (  );
sky130_fd_sc_hd__tap_1 TAP_5044 (  );
sky130_fd_sc_hd__tap_1 TAP_5045 (  );
sky130_fd_sc_hd__tap_1 TAP_5046 (  );
sky130_fd_sc_hd__tap_1 TAP_5047 (  );
sky130_fd_sc_hd__tap_1 TAP_5048 (  );
sky130_fd_sc_hd__tap_1 TAP_5049 (  );
sky130_fd_sc_hd__tap_1 TAP_5050 (  );
sky130_fd_sc_hd__tap_1 TAP_5051 (  );
sky130_fd_sc_hd__tap_1 TAP_5052 (  );
sky130_fd_sc_hd__tap_1 TAP_5053 (  );
sky130_fd_sc_hd__tap_1 TAP_5054 (  );
sky130_fd_sc_hd__tap_1 TAP_5055 (  );
sky130_fd_sc_hd__tap_1 TAP_5056 (  );
sky130_fd_sc_hd__tap_1 TAP_5057 (  );
sky130_fd_sc_hd__tap_1 TAP_5058 (  );
sky130_fd_sc_hd__tap_1 TAP_5059 (  );
sky130_fd_sc_hd__tap_1 TAP_5060 (  );
sky130_fd_sc_hd__tap_1 TAP_5061 (  );
sky130_fd_sc_hd__tap_1 TAP_5062 (  );
sky130_fd_sc_hd__tap_1 TAP_5063 (  );
sky130_fd_sc_hd__tap_1 TAP_5064 (  );
sky130_fd_sc_hd__tap_1 TAP_5065 (  );
sky130_fd_sc_hd__tap_1 TAP_5066 (  );
sky130_fd_sc_hd__tap_1 TAP_5067 (  );
sky130_fd_sc_hd__tap_1 TAP_5068 (  );
sky130_fd_sc_hd__tap_1 TAP_5069 (  );
sky130_fd_sc_hd__tap_1 TAP_5070 (  );
sky130_fd_sc_hd__tap_1 TAP_5071 (  );
sky130_fd_sc_hd__tap_1 TAP_5072 (  );
sky130_fd_sc_hd__tap_1 TAP_5073 (  );
sky130_fd_sc_hd__tap_1 TAP_5074 (  );
sky130_fd_sc_hd__tap_1 TAP_5075 (  );
sky130_fd_sc_hd__tap_1 TAP_5076 (  );
sky130_fd_sc_hd__tap_1 TAP_5077 (  );
sky130_fd_sc_hd__tap_1 TAP_5078 (  );
sky130_fd_sc_hd__tap_1 TAP_5079 (  );
sky130_fd_sc_hd__tap_1 TAP_5080 (  );
sky130_fd_sc_hd__tap_1 TAP_5081 (  );
sky130_fd_sc_hd__tap_1 TAP_5082 (  );
sky130_fd_sc_hd__tap_1 TAP_5083 (  );
sky130_fd_sc_hd__tap_1 TAP_5084 (  );
sky130_fd_sc_hd__tap_1 TAP_5085 (  );
sky130_fd_sc_hd__tap_1 TAP_5086 (  );
sky130_fd_sc_hd__tap_1 TAP_5087 (  );
sky130_fd_sc_hd__tap_1 TAP_5088 (  );
sky130_fd_sc_hd__tap_1 TAP_5089 (  );
sky130_fd_sc_hd__tap_1 TAP_5090 (  );
sky130_fd_sc_hd__tap_1 TAP_5091 (  );
sky130_fd_sc_hd__tap_1 TAP_5092 (  );
sky130_fd_sc_hd__tap_1 TAP_5093 (  );
sky130_fd_sc_hd__tap_1 TAP_5094 (  );
sky130_fd_sc_hd__tap_1 TAP_5095 (  );
sky130_fd_sc_hd__tap_1 TAP_5096 (  );
sky130_fd_sc_hd__tap_1 TAP_5097 (  );
sky130_fd_sc_hd__tap_1 TAP_5098 (  );
sky130_fd_sc_hd__tap_1 TAP_5099 (  );
sky130_fd_sc_hd__tap_1 TAP_5100 (  );
sky130_fd_sc_hd__tap_1 TAP_5101 (  );
sky130_fd_sc_hd__tap_1 TAP_5102 (  );
sky130_fd_sc_hd__tap_1 TAP_5103 (  );
sky130_fd_sc_hd__tap_1 TAP_5104 (  );
sky130_fd_sc_hd__tap_1 TAP_5105 (  );
sky130_fd_sc_hd__tap_1 TAP_5106 (  );
sky130_fd_sc_hd__tap_1 TAP_5107 (  );
sky130_fd_sc_hd__tap_1 TAP_5108 (  );
sky130_fd_sc_hd__tap_1 TAP_5109 (  );
sky130_fd_sc_hd__tap_1 TAP_5110 (  );
sky130_fd_sc_hd__tap_1 TAP_5111 (  );
sky130_fd_sc_hd__tap_1 TAP_5112 (  );
sky130_fd_sc_hd__tap_1 TAP_5113 (  );
sky130_fd_sc_hd__tap_1 TAP_5114 (  );
sky130_fd_sc_hd__tap_1 TAP_5115 (  );
sky130_fd_sc_hd__tap_1 TAP_5116 (  );
sky130_fd_sc_hd__tap_1 TAP_5117 (  );
sky130_fd_sc_hd__tap_1 TAP_5118 (  );
sky130_fd_sc_hd__tap_1 TAP_5119 (  );
sky130_fd_sc_hd__tap_1 TAP_5120 (  );
sky130_fd_sc_hd__tap_1 TAP_5121 (  );
sky130_fd_sc_hd__tap_1 TAP_5122 (  );
sky130_fd_sc_hd__tap_1 TAP_5123 (  );
sky130_fd_sc_hd__tap_1 TAP_5124 (  );
sky130_fd_sc_hd__tap_1 TAP_5125 (  );
sky130_fd_sc_hd__tap_1 TAP_5126 (  );
sky130_fd_sc_hd__tap_1 TAP_5127 (  );
sky130_fd_sc_hd__tap_1 TAP_5128 (  );
sky130_fd_sc_hd__tap_1 TAP_5129 (  );
sky130_fd_sc_hd__tap_1 TAP_5130 (  );
sky130_fd_sc_hd__tap_1 TAP_5131 (  );
sky130_fd_sc_hd__tap_1 TAP_5132 (  );
sky130_fd_sc_hd__tap_1 TAP_5133 (  );
sky130_fd_sc_hd__tap_1 TAP_5134 (  );
sky130_fd_sc_hd__tap_1 TAP_5135 (  );
sky130_fd_sc_hd__tap_1 TAP_5136 (  );
sky130_fd_sc_hd__tap_1 TAP_5137 (  );
sky130_fd_sc_hd__tap_1 TAP_5138 (  );
sky130_fd_sc_hd__tap_1 TAP_5139 (  );
sky130_fd_sc_hd__tap_1 TAP_5140 (  );
sky130_fd_sc_hd__tap_1 TAP_5141 (  );
sky130_fd_sc_hd__tap_1 TAP_5142 (  );
sky130_fd_sc_hd__tap_1 TAP_5143 (  );
sky130_fd_sc_hd__tap_1 TAP_5144 (  );
sky130_fd_sc_hd__tap_1 TAP_5145 (  );
sky130_fd_sc_hd__tap_1 TAP_5146 (  );
sky130_fd_sc_hd__tap_1 TAP_5147 (  );
sky130_fd_sc_hd__tap_1 TAP_5148 (  );
sky130_fd_sc_hd__tap_1 TAP_5149 (  );
sky130_fd_sc_hd__tap_1 TAP_5150 (  );
sky130_fd_sc_hd__tap_1 TAP_5151 (  );
sky130_fd_sc_hd__tap_1 TAP_5152 (  );
sky130_fd_sc_hd__tap_1 TAP_5153 (  );
sky130_fd_sc_hd__tap_1 TAP_5154 (  );
sky130_fd_sc_hd__tap_1 TAP_5155 (  );
sky130_fd_sc_hd__tap_1 TAP_5156 (  );
sky130_fd_sc_hd__tap_1 TAP_5157 (  );
sky130_fd_sc_hd__tap_1 TAP_5158 (  );
sky130_fd_sc_hd__tap_1 TAP_5159 (  );
sky130_fd_sc_hd__tap_1 TAP_5160 (  );
sky130_fd_sc_hd__tap_1 TAP_5161 (  );
sky130_fd_sc_hd__tap_1 TAP_5162 (  );
sky130_fd_sc_hd__tap_1 TAP_5163 (  );
sky130_fd_sc_hd__tap_1 TAP_5164 (  );
sky130_fd_sc_hd__tap_1 TAP_5165 (  );
sky130_fd_sc_hd__tap_1 TAP_5166 (  );
sky130_fd_sc_hd__tap_1 TAP_5167 (  );
sky130_fd_sc_hd__tap_1 TAP_5168 (  );
sky130_fd_sc_hd__tap_1 TAP_5169 (  );
sky130_fd_sc_hd__tap_1 TAP_5170 (  );
sky130_fd_sc_hd__tap_1 TAP_5171 (  );
sky130_fd_sc_hd__tap_1 TAP_5172 (  );
sky130_fd_sc_hd__tap_1 TAP_5173 (  );
sky130_fd_sc_hd__tap_1 TAP_5174 (  );
sky130_fd_sc_hd__tap_1 TAP_5175 (  );
sky130_fd_sc_hd__tap_1 TAP_5176 (  );
sky130_fd_sc_hd__tap_1 TAP_5177 (  );
sky130_fd_sc_hd__tap_1 TAP_5178 (  );
sky130_fd_sc_hd__tap_1 TAP_5179 (  );
sky130_fd_sc_hd__tap_1 TAP_5180 (  );
sky130_fd_sc_hd__tap_1 TAP_5181 (  );
sky130_fd_sc_hd__tap_1 TAP_5182 (  );
sky130_fd_sc_hd__tap_1 TAP_5183 (  );
sky130_fd_sc_hd__tap_1 TAP_5184 (  );
sky130_fd_sc_hd__tap_1 TAP_5185 (  );
sky130_fd_sc_hd__tap_1 TAP_5186 (  );
sky130_fd_sc_hd__tap_1 TAP_5187 (  );
sky130_fd_sc_hd__tap_1 TAP_5188 (  );
sky130_fd_sc_hd__tap_1 TAP_5189 (  );
sky130_fd_sc_hd__tap_1 TAP_5190 (  );
sky130_fd_sc_hd__tap_1 TAP_5191 (  );
sky130_fd_sc_hd__tap_1 TAP_5192 (  );
sky130_fd_sc_hd__tap_1 TAP_5193 (  );
sky130_fd_sc_hd__tap_1 TAP_5194 (  );
sky130_fd_sc_hd__tap_1 TAP_5195 (  );
sky130_fd_sc_hd__tap_1 TAP_5196 (  );
sky130_fd_sc_hd__tap_1 TAP_5197 (  );
sky130_fd_sc_hd__tap_1 TAP_5198 (  );
sky130_fd_sc_hd__tap_1 TAP_5199 (  );
sky130_fd_sc_hd__tap_1 TAP_5200 (  );
sky130_fd_sc_hd__tap_1 TAP_5201 (  );
sky130_fd_sc_hd__tap_1 TAP_5202 (  );
sky130_fd_sc_hd__tap_1 TAP_5203 (  );
sky130_fd_sc_hd__tap_1 TAP_5204 (  );
sky130_fd_sc_hd__tap_1 TAP_5205 (  );
sky130_fd_sc_hd__tap_1 TAP_5206 (  );
sky130_fd_sc_hd__tap_1 TAP_5207 (  );
sky130_fd_sc_hd__tap_1 TAP_5208 (  );
sky130_fd_sc_hd__tap_1 TAP_5209 (  );
sky130_fd_sc_hd__tap_1 TAP_5210 (  );
sky130_fd_sc_hd__tap_1 TAP_5211 (  );
sky130_fd_sc_hd__tap_1 TAP_5212 (  );
sky130_fd_sc_hd__tap_1 TAP_5213 (  );
sky130_fd_sc_hd__tap_1 TAP_5214 (  );
sky130_fd_sc_hd__tap_1 TAP_5215 (  );
sky130_fd_sc_hd__tap_1 TAP_5216 (  );
sky130_fd_sc_hd__tap_1 TAP_5217 (  );
sky130_fd_sc_hd__tap_1 TAP_5218 (  );
sky130_fd_sc_hd__tap_1 TAP_5219 (  );
sky130_fd_sc_hd__tap_1 TAP_5220 (  );
sky130_fd_sc_hd__tap_1 TAP_5221 (  );
sky130_fd_sc_hd__tap_1 TAP_5222 (  );
sky130_fd_sc_hd__tap_1 TAP_5223 (  );
sky130_fd_sc_hd__tap_1 TAP_5224 (  );
sky130_fd_sc_hd__tap_1 TAP_5225 (  );
sky130_fd_sc_hd__tap_1 TAP_5226 (  );
sky130_fd_sc_hd__tap_1 TAP_5227 (  );
sky130_fd_sc_hd__tap_1 TAP_5228 (  );
sky130_fd_sc_hd__tap_1 TAP_5229 (  );
sky130_fd_sc_hd__tap_1 TAP_5230 (  );
sky130_fd_sc_hd__tap_1 TAP_5231 (  );
sky130_fd_sc_hd__tap_1 TAP_5232 (  );
sky130_fd_sc_hd__tap_1 TAP_5233 (  );
sky130_fd_sc_hd__tap_1 TAP_5234 (  );
sky130_fd_sc_hd__tap_1 TAP_5235 (  );
sky130_fd_sc_hd__tap_1 TAP_5236 (  );
sky130_fd_sc_hd__tap_1 TAP_5237 (  );
sky130_fd_sc_hd__tap_1 TAP_5238 (  );
sky130_fd_sc_hd__tap_1 TAP_5239 (  );
sky130_fd_sc_hd__tap_1 TAP_5240 (  );
sky130_fd_sc_hd__tap_1 TAP_5241 (  );
sky130_fd_sc_hd__tap_1 TAP_5242 (  );
sky130_fd_sc_hd__tap_1 TAP_5243 (  );
sky130_fd_sc_hd__tap_1 TAP_5244 (  );
sky130_fd_sc_hd__tap_1 TAP_5245 (  );
sky130_fd_sc_hd__tap_1 TAP_5246 (  );
sky130_fd_sc_hd__tap_1 TAP_5247 (  );
sky130_fd_sc_hd__tap_1 TAP_5248 (  );
sky130_fd_sc_hd__tap_1 TAP_5249 (  );
sky130_fd_sc_hd__tap_1 TAP_5250 (  );
sky130_fd_sc_hd__tap_1 TAP_5251 (  );
sky130_fd_sc_hd__tap_1 TAP_5252 (  );
sky130_fd_sc_hd__tap_1 TAP_5253 (  );
sky130_fd_sc_hd__tap_1 TAP_5254 (  );
sky130_fd_sc_hd__tap_1 TAP_5255 (  );
sky130_fd_sc_hd__tap_1 TAP_5256 (  );
sky130_fd_sc_hd__tap_1 TAP_5257 (  );
sky130_fd_sc_hd__tap_1 TAP_5258 (  );
sky130_fd_sc_hd__tap_1 TAP_5259 (  );
sky130_fd_sc_hd__tap_1 TAP_5260 (  );
sky130_fd_sc_hd__tap_1 TAP_5261 (  );
sky130_fd_sc_hd__tap_1 TAP_5262 (  );
sky130_fd_sc_hd__tap_1 TAP_5263 (  );
sky130_fd_sc_hd__tap_1 TAP_5264 (  );
sky130_fd_sc_hd__tap_1 TAP_5265 (  );
sky130_fd_sc_hd__tap_1 TAP_5266 (  );
sky130_fd_sc_hd__tap_1 TAP_5267 (  );
sky130_fd_sc_hd__tap_1 TAP_5268 (  );
sky130_fd_sc_hd__tap_1 TAP_5269 (  );
sky130_fd_sc_hd__tap_1 TAP_5270 (  );
sky130_fd_sc_hd__tap_1 TAP_5271 (  );
sky130_fd_sc_hd__tap_1 TAP_5272 (  );
sky130_fd_sc_hd__tap_1 TAP_5273 (  );
sky130_fd_sc_hd__tap_1 TAP_5274 (  );
sky130_fd_sc_hd__tap_1 TAP_5275 (  );
sky130_fd_sc_hd__tap_1 TAP_5276 (  );
sky130_fd_sc_hd__tap_1 TAP_5277 (  );
sky130_fd_sc_hd__tap_1 TAP_5278 (  );
sky130_fd_sc_hd__tap_1 TAP_5279 (  );
sky130_fd_sc_hd__tap_1 TAP_5280 (  );
sky130_fd_sc_hd__tap_1 TAP_5281 (  );
sky130_fd_sc_hd__tap_1 TAP_5282 (  );
sky130_fd_sc_hd__tap_1 TAP_5283 (  );
sky130_fd_sc_hd__tap_1 TAP_5284 (  );
sky130_fd_sc_hd__tap_1 TAP_5285 (  );
sky130_fd_sc_hd__tap_1 TAP_5286 (  );
sky130_fd_sc_hd__tap_1 TAP_5287 (  );
sky130_fd_sc_hd__tap_1 TAP_5288 (  );
sky130_fd_sc_hd__tap_1 TAP_5289 (  );
sky130_fd_sc_hd__tap_1 TAP_5290 (  );
sky130_fd_sc_hd__tap_1 TAP_5291 (  );
sky130_fd_sc_hd__tap_1 TAP_5292 (  );
sky130_fd_sc_hd__tap_1 TAP_5293 (  );
sky130_fd_sc_hd__tap_1 TAP_5294 (  );
sky130_fd_sc_hd__tap_1 TAP_5295 (  );
sky130_fd_sc_hd__tap_1 TAP_5296 (  );
sky130_fd_sc_hd__tap_1 TAP_5297 (  );
sky130_fd_sc_hd__tap_1 TAP_5298 (  );
sky130_fd_sc_hd__tap_1 TAP_5299 (  );
sky130_fd_sc_hd__tap_1 TAP_5300 (  );
sky130_fd_sc_hd__tap_1 TAP_5301 (  );
sky130_fd_sc_hd__tap_1 TAP_5302 (  );
sky130_fd_sc_hd__tap_1 TAP_5303 (  );
sky130_fd_sc_hd__tap_1 TAP_5304 (  );
sky130_fd_sc_hd__tap_1 TAP_5305 (  );
sky130_fd_sc_hd__tap_1 TAP_5306 (  );
sky130_fd_sc_hd__tap_1 TAP_5307 (  );
sky130_fd_sc_hd__tap_1 TAP_5308 (  );
sky130_fd_sc_hd__tap_1 TAP_5309 (  );
sky130_fd_sc_hd__tap_1 TAP_5310 (  );
sky130_fd_sc_hd__tap_1 TAP_5311 (  );
sky130_fd_sc_hd__tap_1 TAP_5312 (  );
sky130_fd_sc_hd__tap_1 TAP_5313 (  );
sky130_fd_sc_hd__tap_1 TAP_5314 (  );
sky130_fd_sc_hd__tap_1 TAP_5315 (  );
sky130_fd_sc_hd__tap_1 TAP_5316 (  );
sky130_fd_sc_hd__tap_1 TAP_5317 (  );
sky130_fd_sc_hd__tap_1 TAP_5318 (  );
sky130_fd_sc_hd__tap_1 TAP_5319 (  );
sky130_fd_sc_hd__tap_1 TAP_5320 (  );
sky130_fd_sc_hd__tap_1 TAP_5321 (  );
sky130_fd_sc_hd__tap_1 TAP_5322 (  );
sky130_fd_sc_hd__tap_1 TAP_5323 (  );
sky130_fd_sc_hd__tap_1 TAP_5324 (  );
sky130_fd_sc_hd__tap_1 TAP_5325 (  );
sky130_fd_sc_hd__tap_1 TAP_5326 (  );
sky130_fd_sc_hd__tap_1 TAP_5327 (  );
sky130_fd_sc_hd__tap_1 TAP_5328 (  );
sky130_fd_sc_hd__tap_1 TAP_5329 (  );
sky130_fd_sc_hd__tap_1 TAP_5330 (  );
sky130_fd_sc_hd__tap_1 TAP_5331 (  );
sky130_fd_sc_hd__tap_1 TAP_5332 (  );
sky130_fd_sc_hd__tap_1 TAP_5333 (  );
sky130_fd_sc_hd__tap_1 TAP_5334 (  );
sky130_fd_sc_hd__tap_1 TAP_5335 (  );
sky130_fd_sc_hd__tap_1 TAP_5336 (  );
sky130_fd_sc_hd__tap_1 TAP_5337 (  );
sky130_fd_sc_hd__tap_1 TAP_5338 (  );
sky130_fd_sc_hd__tap_1 TAP_5339 (  );
sky130_fd_sc_hd__tap_1 TAP_5340 (  );
sky130_fd_sc_hd__tap_1 TAP_5341 (  );
sky130_fd_sc_hd__tap_1 TAP_5342 (  );
sky130_fd_sc_hd__tap_1 TAP_5343 (  );
sky130_fd_sc_hd__tap_1 TAP_5344 (  );
sky130_fd_sc_hd__tap_1 TAP_5345 (  );
sky130_fd_sc_hd__tap_1 TAP_5346 (  );
sky130_fd_sc_hd__tap_1 TAP_5347 (  );
sky130_fd_sc_hd__tap_1 TAP_5348 (  );
sky130_fd_sc_hd__tap_1 TAP_5349 (  );
sky130_fd_sc_hd__tap_1 TAP_5350 (  );
sky130_fd_sc_hd__tap_1 TAP_5351 (  );
sky130_fd_sc_hd__tap_1 TAP_5352 (  );
sky130_fd_sc_hd__tap_1 TAP_5353 (  );
sky130_fd_sc_hd__tap_1 TAP_5354 (  );
sky130_fd_sc_hd__tap_1 TAP_5355 (  );
sky130_fd_sc_hd__tap_1 TAP_5356 (  );
sky130_fd_sc_hd__tap_1 TAP_5357 (  );
sky130_fd_sc_hd__tap_1 TAP_5358 (  );
sky130_fd_sc_hd__tap_1 TAP_5359 (  );
sky130_fd_sc_hd__tap_1 TAP_5360 (  );
sky130_fd_sc_hd__tap_1 TAP_5361 (  );
sky130_fd_sc_hd__tap_1 TAP_5362 (  );
sky130_fd_sc_hd__tap_1 TAP_5363 (  );
sky130_fd_sc_hd__tap_1 TAP_5364 (  );
sky130_fd_sc_hd__tap_1 TAP_5365 (  );
sky130_fd_sc_hd__tap_1 TAP_5366 (  );
sky130_fd_sc_hd__tap_1 TAP_5367 (  );
sky130_fd_sc_hd__tap_1 TAP_5368 (  );
sky130_fd_sc_hd__tap_1 TAP_5369 (  );
sky130_fd_sc_hd__tap_1 TAP_5370 (  );
sky130_fd_sc_hd__tap_1 TAP_5371 (  );
sky130_fd_sc_hd__tap_1 TAP_5372 (  );
sky130_fd_sc_hd__tap_1 TAP_5373 (  );
sky130_fd_sc_hd__tap_1 TAP_5374 (  );
sky130_fd_sc_hd__tap_1 TAP_5375 (  );
sky130_fd_sc_hd__tap_1 TAP_5376 (  );
sky130_fd_sc_hd__tap_1 TAP_5377 (  );
sky130_fd_sc_hd__tap_1 TAP_5378 (  );
sky130_fd_sc_hd__tap_1 TAP_5379 (  );
sky130_fd_sc_hd__tap_1 TAP_5380 (  );
sky130_fd_sc_hd__tap_1 TAP_5381 (  );
sky130_fd_sc_hd__tap_1 TAP_5382 (  );
sky130_fd_sc_hd__tap_1 TAP_5383 (  );
sky130_fd_sc_hd__tap_1 TAP_5384 (  );
sky130_fd_sc_hd__tap_1 TAP_5385 (  );
sky130_fd_sc_hd__tap_1 TAP_5386 (  );
sky130_fd_sc_hd__tap_1 TAP_5387 (  );
sky130_fd_sc_hd__tap_1 TAP_5388 (  );
sky130_fd_sc_hd__tap_1 TAP_5389 (  );
sky130_fd_sc_hd__tap_1 TAP_5390 (  );
sky130_fd_sc_hd__tap_1 TAP_5391 (  );
sky130_fd_sc_hd__tap_1 TAP_5392 (  );
sky130_fd_sc_hd__tap_1 TAP_5393 (  );
sky130_fd_sc_hd__tap_1 TAP_5394 (  );
sky130_fd_sc_hd__tap_1 TAP_5395 (  );
sky130_fd_sc_hd__tap_1 TAP_5396 (  );
sky130_fd_sc_hd__tap_1 TAP_5397 (  );
sky130_fd_sc_hd__tap_1 TAP_5398 (  );
sky130_fd_sc_hd__tap_1 TAP_5399 (  );
sky130_fd_sc_hd__tap_1 TAP_5400 (  );
sky130_fd_sc_hd__tap_1 TAP_5401 (  );
sky130_fd_sc_hd__tap_1 TAP_5402 (  );
sky130_fd_sc_hd__tap_1 TAP_5403 (  );
sky130_fd_sc_hd__tap_1 TAP_5404 (  );
sky130_fd_sc_hd__tap_1 TAP_5405 (  );
sky130_fd_sc_hd__tap_1 TAP_5406 (  );
sky130_fd_sc_hd__tap_1 TAP_5407 (  );
sky130_fd_sc_hd__tap_1 TAP_5408 (  );
sky130_fd_sc_hd__tap_1 TAP_5409 (  );
sky130_fd_sc_hd__tap_1 TAP_5410 (  );
sky130_fd_sc_hd__tap_1 TAP_5411 (  );
sky130_fd_sc_hd__tap_1 TAP_5412 (  );
sky130_fd_sc_hd__tap_1 TAP_5413 (  );
sky130_fd_sc_hd__tap_1 TAP_5414 (  );
sky130_fd_sc_hd__tap_1 TAP_5415 (  );
sky130_fd_sc_hd__tap_1 TAP_5416 (  );
sky130_fd_sc_hd__tap_1 TAP_5417 (  );
sky130_fd_sc_hd__tap_1 TAP_5418 (  );
sky130_fd_sc_hd__tap_1 TAP_5419 (  );
sky130_fd_sc_hd__tap_1 TAP_5420 (  );
sky130_fd_sc_hd__tap_1 TAP_5421 (  );
sky130_fd_sc_hd__tap_1 TAP_5422 (  );
sky130_fd_sc_hd__tap_1 TAP_5423 (  );
sky130_fd_sc_hd__tap_1 TAP_5424 (  );
sky130_fd_sc_hd__tap_1 TAP_5425 (  );
sky130_fd_sc_hd__tap_1 TAP_5426 (  );
sky130_fd_sc_hd__tap_1 TAP_5427 (  );
sky130_fd_sc_hd__tap_1 TAP_5428 (  );
sky130_fd_sc_hd__tap_1 TAP_5429 (  );
sky130_fd_sc_hd__tap_1 TAP_5430 (  );
sky130_fd_sc_hd__tap_1 TAP_5431 (  );
sky130_fd_sc_hd__tap_1 TAP_5432 (  );
sky130_fd_sc_hd__tap_1 TAP_5433 (  );
sky130_fd_sc_hd__tap_1 TAP_5434 (  );
sky130_fd_sc_hd__tap_1 TAP_5435 (  );
sky130_fd_sc_hd__tap_1 TAP_5436 (  );
sky130_fd_sc_hd__tap_1 TAP_5437 (  );
sky130_fd_sc_hd__tap_1 TAP_5438 (  );
sky130_fd_sc_hd__tap_1 TAP_5439 (  );
sky130_fd_sc_hd__tap_1 TAP_5440 (  );
sky130_fd_sc_hd__tap_1 TAP_5441 (  );
sky130_fd_sc_hd__tap_1 TAP_5442 (  );
sky130_fd_sc_hd__tap_1 TAP_5443 (  );
sky130_fd_sc_hd__tap_1 TAP_5444 (  );
sky130_fd_sc_hd__tap_1 TAP_5445 (  );
sky130_fd_sc_hd__tap_1 TAP_5446 (  );
sky130_fd_sc_hd__tap_1 TAP_5447 (  );
sky130_fd_sc_hd__tap_1 TAP_5448 (  );
sky130_fd_sc_hd__tap_1 TAP_5449 (  );
sky130_fd_sc_hd__tap_1 TAP_5450 (  );
sky130_fd_sc_hd__tap_1 TAP_5451 (  );
sky130_fd_sc_hd__tap_1 TAP_5452 (  );
sky130_fd_sc_hd__tap_1 TAP_5453 (  );
sky130_fd_sc_hd__tap_1 TAP_5454 (  );
sky130_fd_sc_hd__tap_1 TAP_5455 (  );
sky130_fd_sc_hd__tap_1 TAP_5456 (  );
sky130_fd_sc_hd__tap_1 TAP_5457 (  );
sky130_fd_sc_hd__tap_1 TAP_5458 (  );
sky130_fd_sc_hd__tap_1 TAP_5459 (  );
sky130_fd_sc_hd__tap_1 TAP_5460 (  );
sky130_fd_sc_hd__tap_1 TAP_5461 (  );
sky130_fd_sc_hd__tap_1 TAP_5462 (  );
sky130_fd_sc_hd__tap_1 TAP_5463 (  );
sky130_fd_sc_hd__tap_1 TAP_5464 (  );
sky130_fd_sc_hd__tap_1 TAP_5465 (  );
sky130_fd_sc_hd__tap_1 TAP_5466 (  );
sky130_fd_sc_hd__tap_1 TAP_5467 (  );
sky130_fd_sc_hd__tap_1 TAP_5468 (  );
sky130_fd_sc_hd__tap_1 TAP_5469 (  );
sky130_fd_sc_hd__tap_1 TAP_5470 (  );
sky130_fd_sc_hd__tap_1 TAP_5471 (  );
sky130_fd_sc_hd__tap_1 TAP_5472 (  );
sky130_fd_sc_hd__tap_1 TAP_5473 (  );
sky130_fd_sc_hd__tap_1 TAP_5474 (  );
sky130_fd_sc_hd__tap_1 TAP_5475 (  );
sky130_fd_sc_hd__tap_1 TAP_5476 (  );
sky130_fd_sc_hd__tap_1 TAP_5477 (  );
sky130_fd_sc_hd__tap_1 TAP_5478 (  );
sky130_fd_sc_hd__tap_1 TAP_5479 (  );
sky130_fd_sc_hd__tap_1 TAP_5480 (  );
sky130_fd_sc_hd__tap_1 TAP_5481 (  );
sky130_fd_sc_hd__tap_1 TAP_5482 (  );
sky130_fd_sc_hd__tap_1 TAP_5483 (  );
sky130_fd_sc_hd__tap_1 TAP_5484 (  );
sky130_fd_sc_hd__tap_1 TAP_5485 (  );
sky130_fd_sc_hd__tap_1 TAP_5486 (  );
sky130_fd_sc_hd__tap_1 TAP_5487 (  );
sky130_fd_sc_hd__tap_1 TAP_5488 (  );
sky130_fd_sc_hd__tap_1 TAP_5489 (  );
sky130_fd_sc_hd__tap_1 TAP_5490 (  );
sky130_fd_sc_hd__tap_1 TAP_5491 (  );
sky130_fd_sc_hd__tap_1 TAP_5492 (  );
sky130_fd_sc_hd__tap_1 TAP_5493 (  );
sky130_fd_sc_hd__tap_1 TAP_5494 (  );
sky130_fd_sc_hd__tap_1 TAP_5495 (  );
sky130_fd_sc_hd__tap_1 TAP_5496 (  );
sky130_fd_sc_hd__tap_1 TAP_5497 (  );
sky130_fd_sc_hd__tap_1 TAP_5498 (  );
sky130_fd_sc_hd__tap_1 TAP_5499 (  );
sky130_fd_sc_hd__tap_1 TAP_5500 (  );
sky130_fd_sc_hd__tap_1 TAP_5501 (  );
sky130_fd_sc_hd__tap_1 TAP_5502 (  );
sky130_fd_sc_hd__tap_1 TAP_5503 (  );
sky130_fd_sc_hd__tap_1 TAP_5504 (  );
sky130_fd_sc_hd__tap_1 TAP_5505 (  );
sky130_fd_sc_hd__tap_1 TAP_5506 (  );
sky130_fd_sc_hd__tap_1 TAP_5507 (  );
sky130_fd_sc_hd__tap_1 TAP_5508 (  );
sky130_fd_sc_hd__tap_1 TAP_5509 (  );
sky130_fd_sc_hd__tap_1 TAP_5510 (  );
sky130_fd_sc_hd__tap_1 TAP_5511 (  );
sky130_fd_sc_hd__tap_1 TAP_5512 (  );
sky130_fd_sc_hd__tap_1 TAP_5513 (  );
sky130_fd_sc_hd__tap_1 TAP_5514 (  );
sky130_fd_sc_hd__tap_1 TAP_5515 (  );
sky130_fd_sc_hd__tap_1 TAP_5516 (  );
sky130_fd_sc_hd__tap_1 TAP_5517 (  );
sky130_fd_sc_hd__tap_1 TAP_5518 (  );
sky130_fd_sc_hd__tap_1 TAP_5519 (  );
sky130_fd_sc_hd__tap_1 TAP_5520 (  );
sky130_fd_sc_hd__tap_1 TAP_5521 (  );
sky130_fd_sc_hd__tap_1 TAP_5522 (  );
sky130_fd_sc_hd__tap_1 TAP_5523 (  );
sky130_fd_sc_hd__tap_1 TAP_5524 (  );
sky130_fd_sc_hd__tap_1 TAP_5525 (  );
sky130_fd_sc_hd__tap_1 TAP_5526 (  );
sky130_fd_sc_hd__tap_1 TAP_5527 (  );
sky130_fd_sc_hd__tap_1 TAP_5528 (  );
sky130_fd_sc_hd__tap_1 TAP_5529 (  );
sky130_fd_sc_hd__tap_1 TAP_5530 (  );
sky130_fd_sc_hd__tap_1 TAP_5531 (  );
sky130_fd_sc_hd__tap_1 TAP_5532 (  );
sky130_fd_sc_hd__tap_1 TAP_5533 (  );
sky130_fd_sc_hd__tap_1 TAP_5534 (  );
sky130_fd_sc_hd__tap_1 TAP_5535 (  );
sky130_fd_sc_hd__tap_1 TAP_5536 (  );
sky130_fd_sc_hd__tap_1 TAP_5537 (  );
sky130_fd_sc_hd__tap_1 TAP_5538 (  );
sky130_fd_sc_hd__tap_1 TAP_5539 (  );
sky130_fd_sc_hd__tap_1 TAP_5540 (  );
sky130_fd_sc_hd__tap_1 TAP_5541 (  );
sky130_fd_sc_hd__tap_1 TAP_5542 (  );
sky130_fd_sc_hd__tap_1 TAP_5543 (  );
sky130_fd_sc_hd__tap_1 TAP_5544 (  );
sky130_fd_sc_hd__tap_1 TAP_5545 (  );
sky130_fd_sc_hd__tap_1 TAP_5546 (  );
sky130_fd_sc_hd__tap_1 TAP_5547 (  );
sky130_fd_sc_hd__tap_1 TAP_5548 (  );
sky130_fd_sc_hd__tap_1 TAP_5549 (  );
sky130_fd_sc_hd__tap_1 TAP_5550 (  );
sky130_fd_sc_hd__tap_1 TAP_5551 (  );
sky130_fd_sc_hd__tap_1 TAP_5552 (  );
sky130_fd_sc_hd__tap_1 TAP_5553 (  );
sky130_fd_sc_hd__tap_1 TAP_5554 (  );
sky130_fd_sc_hd__tap_1 TAP_5555 (  );
sky130_fd_sc_hd__tap_1 TAP_5556 (  );
sky130_fd_sc_hd__tap_1 TAP_5557 (  );
sky130_fd_sc_hd__tap_1 TAP_5558 (  );
sky130_fd_sc_hd__tap_1 TAP_5559 (  );
sky130_fd_sc_hd__tap_1 TAP_5560 (  );
sky130_fd_sc_hd__tap_1 TAP_5561 (  );
sky130_fd_sc_hd__tap_1 TAP_5562 (  );
sky130_fd_sc_hd__tap_1 TAP_5563 (  );
sky130_fd_sc_hd__tap_1 TAP_5564 (  );
sky130_fd_sc_hd__tap_1 TAP_5565 (  );
sky130_fd_sc_hd__tap_1 TAP_5566 (  );
sky130_fd_sc_hd__tap_1 TAP_5567 (  );
sky130_fd_sc_hd__tap_1 TAP_5568 (  );
sky130_fd_sc_hd__tap_1 TAP_5569 (  );
sky130_fd_sc_hd__tap_1 TAP_5570 (  );
sky130_fd_sc_hd__tap_1 TAP_5571 (  );
sky130_fd_sc_hd__tap_1 TAP_5572 (  );
sky130_fd_sc_hd__tap_1 TAP_5573 (  );
sky130_fd_sc_hd__tap_1 TAP_5574 (  );
sky130_fd_sc_hd__tap_1 TAP_5575 (  );
sky130_fd_sc_hd__tap_1 TAP_5576 (  );
sky130_fd_sc_hd__tap_1 TAP_5577 (  );
sky130_fd_sc_hd__tap_1 TAP_5578 (  );
sky130_fd_sc_hd__tap_1 TAP_5579 (  );
sky130_fd_sc_hd__tap_1 TAP_5580 (  );
sky130_fd_sc_hd__tap_1 TAP_5581 (  );
sky130_fd_sc_hd__tap_1 TAP_5582 (  );
sky130_fd_sc_hd__tap_1 TAP_5583 (  );
sky130_fd_sc_hd__tap_1 TAP_5584 (  );
sky130_fd_sc_hd__tap_1 TAP_5585 (  );
sky130_fd_sc_hd__tap_1 TAP_5586 (  );
sky130_fd_sc_hd__tap_1 TAP_5587 (  );
sky130_fd_sc_hd__tap_1 TAP_5588 (  );
sky130_fd_sc_hd__tap_1 TAP_5589 (  );
sky130_fd_sc_hd__tap_1 TAP_5590 (  );
sky130_fd_sc_hd__tap_1 TAP_5591 (  );
sky130_fd_sc_hd__tap_1 TAP_5592 (  );
sky130_fd_sc_hd__tap_1 TAP_5593 (  );
sky130_fd_sc_hd__tap_1 TAP_5594 (  );
sky130_fd_sc_hd__tap_1 TAP_5595 (  );
sky130_fd_sc_hd__tap_1 TAP_5596 (  );
sky130_fd_sc_hd__tap_1 TAP_5597 (  );
sky130_fd_sc_hd__tap_1 TAP_5598 (  );
sky130_fd_sc_hd__tap_1 TAP_5599 (  );
sky130_fd_sc_hd__tap_1 TAP_5600 (  );
sky130_fd_sc_hd__tap_1 TAP_5601 (  );
sky130_fd_sc_hd__tap_1 TAP_5602 (  );
sky130_fd_sc_hd__tap_1 TAP_5603 (  );
sky130_fd_sc_hd__tap_1 TAP_5604 (  );
sky130_fd_sc_hd__tap_1 TAP_5605 (  );
sky130_fd_sc_hd__tap_1 TAP_5606 (  );
sky130_fd_sc_hd__tap_1 TAP_5607 (  );
sky130_fd_sc_hd__tap_1 TAP_5608 (  );
sky130_fd_sc_hd__tap_1 TAP_5609 (  );
sky130_fd_sc_hd__tap_1 TAP_5610 (  );
sky130_fd_sc_hd__tap_1 TAP_5611 (  );
sky130_fd_sc_hd__tap_1 TAP_5612 (  );
sky130_fd_sc_hd__tap_1 TAP_5613 (  );
sky130_fd_sc_hd__tap_1 TAP_5614 (  );
sky130_fd_sc_hd__tap_1 TAP_5615 (  );
sky130_fd_sc_hd__tap_1 TAP_5616 (  );
sky130_fd_sc_hd__tap_1 TAP_5617 (  );
sky130_fd_sc_hd__tap_1 TAP_5618 (  );
sky130_fd_sc_hd__tap_1 TAP_5619 (  );
sky130_fd_sc_hd__tap_1 TAP_5620 (  );
sky130_fd_sc_hd__tap_1 TAP_5621 (  );
sky130_fd_sc_hd__tap_1 TAP_5622 (  );
sky130_fd_sc_hd__tap_1 TAP_5623 (  );
sky130_fd_sc_hd__tap_1 TAP_5624 (  );
sky130_fd_sc_hd__tap_1 TAP_5625 (  );
sky130_fd_sc_hd__tap_1 TAP_5626 (  );
sky130_fd_sc_hd__tap_1 TAP_5627 (  );
sky130_fd_sc_hd__tap_1 TAP_5628 (  );
sky130_fd_sc_hd__tap_1 TAP_5629 (  );
sky130_fd_sc_hd__tap_1 TAP_5630 (  );
sky130_fd_sc_hd__tap_1 TAP_5631 (  );
sky130_fd_sc_hd__tap_1 TAP_5632 (  );
sky130_fd_sc_hd__tap_1 TAP_5633 (  );
sky130_fd_sc_hd__tap_1 TAP_5634 (  );
sky130_fd_sc_hd__tap_1 TAP_5635 (  );
sky130_fd_sc_hd__tap_1 TAP_5636 (  );
sky130_fd_sc_hd__tap_1 TAP_5637 (  );
sky130_fd_sc_hd__tap_1 TAP_5638 (  );
sky130_fd_sc_hd__tap_1 TAP_5639 (  );
sky130_fd_sc_hd__tap_1 TAP_5640 (  );
sky130_fd_sc_hd__tap_1 TAP_5641 (  );
sky130_fd_sc_hd__tap_1 TAP_5642 (  );
sky130_fd_sc_hd__tap_1 TAP_5643 (  );
sky130_fd_sc_hd__tap_1 TAP_5644 (  );
sky130_fd_sc_hd__tap_1 TAP_5645 (  );
sky130_fd_sc_hd__tap_1 TAP_5646 (  );
sky130_fd_sc_hd__tap_1 TAP_5647 (  );
sky130_fd_sc_hd__tap_1 TAP_5648 (  );
sky130_fd_sc_hd__tap_1 TAP_5649 (  );
sky130_fd_sc_hd__tap_1 TAP_5650 (  );
sky130_fd_sc_hd__tap_1 TAP_5651 (  );
sky130_fd_sc_hd__tap_1 TAP_5652 (  );
sky130_fd_sc_hd__tap_1 TAP_5653 (  );
sky130_fd_sc_hd__tap_1 TAP_5654 (  );
sky130_fd_sc_hd__tap_1 TAP_5655 (  );
sky130_fd_sc_hd__tap_1 TAP_5656 (  );
sky130_fd_sc_hd__tap_1 TAP_5657 (  );
sky130_fd_sc_hd__tap_1 TAP_5658 (  );
sky130_fd_sc_hd__tap_1 TAP_5659 (  );
sky130_fd_sc_hd__tap_1 TAP_5660 (  );
sky130_fd_sc_hd__tap_1 TAP_5661 (  );
sky130_fd_sc_hd__tap_1 TAP_5662 (  );
sky130_fd_sc_hd__tap_1 TAP_5663 (  );
sky130_fd_sc_hd__tap_1 TAP_5664 (  );
sky130_fd_sc_hd__tap_1 TAP_5665 (  );
sky130_fd_sc_hd__tap_1 TAP_5666 (  );
sky130_fd_sc_hd__tap_1 TAP_5667 (  );
sky130_fd_sc_hd__tap_1 TAP_5668 (  );
sky130_fd_sc_hd__tap_1 TAP_5669 (  );
sky130_fd_sc_hd__tap_1 TAP_5670 (  );
sky130_fd_sc_hd__tap_1 TAP_5671 (  );
sky130_fd_sc_hd__tap_1 TAP_5672 (  );
sky130_fd_sc_hd__tap_1 TAP_5673 (  );
sky130_fd_sc_hd__tap_1 TAP_5674 (  );
sky130_fd_sc_hd__tap_1 TAP_5675 (  );
sky130_fd_sc_hd__tap_1 TAP_5676 (  );
sky130_fd_sc_hd__tap_1 TAP_5677 (  );
sky130_fd_sc_hd__tap_1 TAP_5678 (  );
sky130_fd_sc_hd__tap_1 TAP_5679 (  );
sky130_fd_sc_hd__tap_1 TAP_5680 (  );
sky130_fd_sc_hd__tap_1 TAP_5681 (  );
sky130_fd_sc_hd__tap_1 TAP_5682 (  );
sky130_fd_sc_hd__tap_1 TAP_5683 (  );
sky130_fd_sc_hd__tap_1 TAP_5684 (  );
sky130_fd_sc_hd__tap_1 TAP_5685 (  );
sky130_fd_sc_hd__tap_1 TAP_5686 (  );
sky130_fd_sc_hd__tap_1 TAP_5687 (  );
sky130_fd_sc_hd__tap_1 TAP_5688 (  );
sky130_fd_sc_hd__tap_1 TAP_5689 (  );
sky130_fd_sc_hd__tap_1 TAP_5690 (  );
sky130_fd_sc_hd__tap_1 TAP_5691 (  );
sky130_fd_sc_hd__tap_1 TAP_5692 (  );
sky130_fd_sc_hd__tap_1 TAP_5693 (  );
sky130_fd_sc_hd__tap_1 TAP_5694 (  );
sky130_fd_sc_hd__tap_1 TAP_5695 (  );
sky130_fd_sc_hd__tap_1 TAP_5696 (  );
sky130_fd_sc_hd__tap_1 TAP_5697 (  );
sky130_fd_sc_hd__tap_1 TAP_5698 (  );
sky130_fd_sc_hd__tap_1 TAP_5699 (  );
sky130_fd_sc_hd__tap_1 TAP_5700 (  );
sky130_fd_sc_hd__tap_1 TAP_5701 (  );
sky130_fd_sc_hd__tap_1 TAP_5702 (  );
sky130_fd_sc_hd__tap_1 TAP_5703 (  );
sky130_fd_sc_hd__tap_1 TAP_5704 (  );
sky130_fd_sc_hd__tap_1 TAP_5705 (  );
sky130_fd_sc_hd__tap_1 TAP_5706 (  );
sky130_fd_sc_hd__tap_1 TAP_5707 (  );
sky130_fd_sc_hd__tap_1 TAP_5708 (  );
sky130_fd_sc_hd__tap_1 TAP_5709 (  );
sky130_fd_sc_hd__tap_1 TAP_5710 (  );
sky130_fd_sc_hd__tap_1 TAP_5711 (  );
sky130_fd_sc_hd__tap_1 TAP_5712 (  );
sky130_fd_sc_hd__tap_1 TAP_5713 (  );
sky130_fd_sc_hd__tap_1 TAP_5714 (  );
sky130_fd_sc_hd__tap_1 TAP_5715 (  );
sky130_fd_sc_hd__tap_1 TAP_5716 (  );
sky130_fd_sc_hd__tap_1 TAP_5717 (  );
sky130_fd_sc_hd__tap_1 TAP_5718 (  );
sky130_fd_sc_hd__tap_1 TAP_5719 (  );
sky130_fd_sc_hd__tap_1 TAP_5720 (  );
sky130_fd_sc_hd__tap_1 TAP_5721 (  );
sky130_fd_sc_hd__tap_1 TAP_5722 (  );
sky130_fd_sc_hd__tap_1 TAP_5723 (  );
sky130_fd_sc_hd__tap_1 TAP_5724 (  );
sky130_fd_sc_hd__tap_1 TAP_5725 (  );
sky130_fd_sc_hd__tap_1 TAP_5726 (  );
sky130_fd_sc_hd__tap_1 TAP_5727 (  );
sky130_fd_sc_hd__tap_1 TAP_5728 (  );
sky130_fd_sc_hd__tap_1 TAP_5729 (  );
sky130_fd_sc_hd__tap_1 TAP_5730 (  );
sky130_fd_sc_hd__tap_1 TAP_5731 (  );
sky130_fd_sc_hd__tap_1 TAP_5732 (  );
sky130_fd_sc_hd__tap_1 TAP_5733 (  );
sky130_fd_sc_hd__tap_1 TAP_5734 (  );
sky130_fd_sc_hd__tap_1 TAP_5735 (  );
sky130_fd_sc_hd__tap_1 TAP_5736 (  );
sky130_fd_sc_hd__tap_1 TAP_5737 (  );
sky130_fd_sc_hd__tap_1 TAP_5738 (  );
sky130_fd_sc_hd__tap_1 TAP_5739 (  );
sky130_fd_sc_hd__tap_1 TAP_5740 (  );
sky130_fd_sc_hd__tap_1 TAP_5741 (  );
sky130_fd_sc_hd__tap_1 TAP_5742 (  );
sky130_fd_sc_hd__tap_1 TAP_5743 (  );
sky130_fd_sc_hd__tap_1 TAP_5744 (  );
sky130_fd_sc_hd__tap_1 TAP_5745 (  );
sky130_fd_sc_hd__tap_1 TAP_5746 (  );
sky130_fd_sc_hd__tap_1 TAP_5747 (  );
sky130_fd_sc_hd__tap_1 TAP_5748 (  );
sky130_fd_sc_hd__tap_1 TAP_5749 (  );
sky130_fd_sc_hd__tap_1 TAP_5750 (  );
sky130_fd_sc_hd__tap_1 TAP_5751 (  );
sky130_fd_sc_hd__tap_1 TAP_5752 (  );
sky130_fd_sc_hd__tap_1 TAP_5753 (  );
sky130_fd_sc_hd__tap_1 TAP_5754 (  );
sky130_fd_sc_hd__tap_1 TAP_5755 (  );
sky130_fd_sc_hd__tap_1 TAP_5756 (  );
sky130_fd_sc_hd__tap_1 TAP_5757 (  );
sky130_fd_sc_hd__tap_1 TAP_5758 (  );
sky130_fd_sc_hd__tap_1 TAP_5759 (  );
sky130_fd_sc_hd__tap_1 TAP_5760 (  );
sky130_fd_sc_hd__tap_1 TAP_5761 (  );
sky130_fd_sc_hd__tap_1 TAP_5762 (  );
sky130_fd_sc_hd__tap_1 TAP_5763 (  );
sky130_fd_sc_hd__tap_1 TAP_5764 (  );
sky130_fd_sc_hd__tap_1 TAP_5765 (  );
sky130_fd_sc_hd__tap_1 TAP_5766 (  );
sky130_fd_sc_hd__tap_1 TAP_5767 (  );
sky130_fd_sc_hd__tap_1 TAP_5768 (  );
sky130_fd_sc_hd__tap_1 TAP_5769 (  );
sky130_fd_sc_hd__tap_1 TAP_5770 (  );
sky130_fd_sc_hd__tap_1 TAP_5771 (  );
sky130_fd_sc_hd__tap_1 TAP_5772 (  );
sky130_fd_sc_hd__tap_1 TAP_5773 (  );
sky130_fd_sc_hd__tap_1 TAP_5774 (  );
sky130_fd_sc_hd__tap_1 TAP_5775 (  );
sky130_fd_sc_hd__tap_1 TAP_5776 (  );
sky130_fd_sc_hd__tap_1 TAP_5777 (  );
sky130_fd_sc_hd__tap_1 TAP_5778 (  );
sky130_fd_sc_hd__tap_1 TAP_5779 (  );
sky130_fd_sc_hd__tap_1 TAP_5780 (  );
sky130_fd_sc_hd__tap_1 TAP_5781 (  );
sky130_fd_sc_hd__tap_1 TAP_5782 (  );
sky130_fd_sc_hd__tap_1 TAP_5783 (  );
sky130_fd_sc_hd__tap_1 TAP_5784 (  );
sky130_fd_sc_hd__tap_1 TAP_5785 (  );
sky130_fd_sc_hd__tap_1 TAP_5786 (  );
sky130_fd_sc_hd__tap_1 TAP_5787 (  );
sky130_fd_sc_hd__tap_1 TAP_5788 (  );
sky130_fd_sc_hd__tap_1 TAP_5789 (  );
sky130_fd_sc_hd__tap_1 TAP_5790 (  );
sky130_fd_sc_hd__tap_1 TAP_5791 (  );
sky130_fd_sc_hd__tap_1 TAP_5792 (  );
sky130_fd_sc_hd__tap_1 TAP_5793 (  );
sky130_fd_sc_hd__tap_1 TAP_5794 (  );
sky130_fd_sc_hd__tap_1 TAP_5795 (  );
sky130_fd_sc_hd__tap_1 TAP_5796 (  );
sky130_fd_sc_hd__tap_1 TAP_5797 (  );
sky130_fd_sc_hd__tap_1 TAP_5798 (  );
sky130_fd_sc_hd__tap_1 TAP_5799 (  );
sky130_fd_sc_hd__tap_1 TAP_5800 (  );
sky130_fd_sc_hd__tap_1 TAP_5801 (  );
sky130_fd_sc_hd__tap_1 TAP_5802 (  );
sky130_fd_sc_hd__tap_1 TAP_5803 (  );
sky130_fd_sc_hd__tap_1 TAP_5804 (  );
sky130_fd_sc_hd__tap_1 TAP_5805 (  );
sky130_fd_sc_hd__tap_1 TAP_5806 (  );
sky130_fd_sc_hd__tap_1 TAP_5807 (  );
sky130_fd_sc_hd__tap_1 TAP_5808 (  );
sky130_fd_sc_hd__tap_1 TAP_5809 (  );
sky130_fd_sc_hd__tap_1 TAP_5810 (  );
sky130_fd_sc_hd__tap_1 TAP_5811 (  );
sky130_fd_sc_hd__tap_1 TAP_5812 (  );
sky130_fd_sc_hd__tap_1 TAP_5813 (  );
sky130_fd_sc_hd__tap_1 TAP_5814 (  );
sky130_fd_sc_hd__tap_1 TAP_5815 (  );
sky130_fd_sc_hd__tap_1 TAP_5816 (  );
sky130_fd_sc_hd__tap_1 TAP_5817 (  );
sky130_fd_sc_hd__tap_1 TAP_5818 (  );
sky130_fd_sc_hd__tap_1 TAP_5819 (  );
sky130_fd_sc_hd__tap_1 TAP_5820 (  );
sky130_fd_sc_hd__tap_1 TAP_5821 (  );
sky130_fd_sc_hd__tap_1 TAP_5822 (  );
sky130_fd_sc_hd__tap_1 TAP_5823 (  );
sky130_fd_sc_hd__tap_1 TAP_5824 (  );
sky130_fd_sc_hd__tap_1 TAP_5825 (  );
sky130_fd_sc_hd__tap_1 TAP_5826 (  );
sky130_fd_sc_hd__tap_1 TAP_5827 (  );
sky130_fd_sc_hd__tap_1 TAP_5828 (  );
sky130_fd_sc_hd__tap_1 TAP_5829 (  );
sky130_fd_sc_hd__tap_1 TAP_5830 (  );
sky130_fd_sc_hd__tap_1 TAP_5831 (  );
sky130_fd_sc_hd__tap_1 TAP_5832 (  );
sky130_fd_sc_hd__tap_1 TAP_5833 (  );
sky130_fd_sc_hd__tap_1 TAP_5834 (  );
sky130_fd_sc_hd__tap_1 TAP_5835 (  );
sky130_fd_sc_hd__tap_1 TAP_5836 (  );
sky130_fd_sc_hd__tap_1 TAP_5837 (  );
sky130_fd_sc_hd__tap_1 TAP_5838 (  );
sky130_fd_sc_hd__tap_1 TAP_5839 (  );
sky130_fd_sc_hd__tap_1 TAP_5840 (  );
sky130_fd_sc_hd__tap_1 TAP_5841 (  );
sky130_fd_sc_hd__tap_1 TAP_5842 (  );
sky130_fd_sc_hd__tap_1 TAP_5843 (  );
sky130_fd_sc_hd__tap_1 TAP_5844 (  );
sky130_fd_sc_hd__tap_1 TAP_5845 (  );
sky130_fd_sc_hd__tap_1 TAP_5846 (  );
sky130_fd_sc_hd__tap_1 TAP_5847 (  );
sky130_fd_sc_hd__tap_1 TAP_5848 (  );
sky130_fd_sc_hd__tap_1 TAP_5849 (  );
sky130_fd_sc_hd__tap_1 TAP_5850 (  );
sky130_fd_sc_hd__tap_1 TAP_5851 (  );
sky130_fd_sc_hd__tap_1 TAP_5852 (  );
sky130_fd_sc_hd__tap_1 TAP_5853 (  );
sky130_fd_sc_hd__tap_1 TAP_5854 (  );
sky130_fd_sc_hd__tap_1 TAP_5855 (  );
sky130_fd_sc_hd__tap_1 TAP_5856 (  );
sky130_fd_sc_hd__tap_1 TAP_5857 (  );
sky130_fd_sc_hd__tap_1 TAP_5858 (  );
sky130_fd_sc_hd__tap_1 TAP_5859 (  );
sky130_fd_sc_hd__tap_1 TAP_5860 (  );
sky130_fd_sc_hd__tap_1 TAP_5861 (  );
sky130_fd_sc_hd__tap_1 TAP_5862 (  );
sky130_fd_sc_hd__tap_1 TAP_5863 (  );
sky130_fd_sc_hd__tap_1 TAP_5864 (  );
sky130_fd_sc_hd__tap_1 TAP_5865 (  );
sky130_fd_sc_hd__tap_1 TAP_5866 (  );
sky130_fd_sc_hd__tap_1 TAP_5867 (  );
sky130_fd_sc_hd__tap_1 TAP_5868 (  );
sky130_fd_sc_hd__tap_1 TAP_5869 (  );
sky130_fd_sc_hd__tap_1 TAP_5870 (  );
sky130_fd_sc_hd__tap_1 TAP_5871 (  );
sky130_fd_sc_hd__tap_1 TAP_5872 (  );
sky130_fd_sc_hd__tap_1 TAP_5873 (  );
sky130_fd_sc_hd__tap_1 TAP_5874 (  );
sky130_fd_sc_hd__tap_1 TAP_5875 (  );
sky130_fd_sc_hd__tap_1 TAP_5876 (  );
sky130_fd_sc_hd__tap_1 TAP_5877 (  );
sky130_fd_sc_hd__tap_1 TAP_5878 (  );
sky130_fd_sc_hd__tap_1 TAP_5879 (  );
sky130_fd_sc_hd__tap_1 TAP_5880 (  );
sky130_fd_sc_hd__tap_1 TAP_5881 (  );
sky130_fd_sc_hd__tap_1 TAP_5882 (  );
sky130_fd_sc_hd__tap_1 TAP_5883 (  );
sky130_fd_sc_hd__tap_1 TAP_5884 (  );
sky130_fd_sc_hd__tap_1 TAP_5885 (  );
sky130_fd_sc_hd__tap_1 TAP_5886 (  );
sky130_fd_sc_hd__tap_1 TAP_5887 (  );
sky130_fd_sc_hd__tap_1 TAP_5888 (  );
sky130_fd_sc_hd__tap_1 TAP_5889 (  );
sky130_fd_sc_hd__tap_1 TAP_5890 (  );
sky130_fd_sc_hd__tap_1 TAP_5891 (  );
sky130_fd_sc_hd__tap_1 TAP_5892 (  );
sky130_fd_sc_hd__tap_1 TAP_5893 (  );
sky130_fd_sc_hd__tap_1 TAP_5894 (  );
sky130_fd_sc_hd__tap_1 TAP_5895 (  );
sky130_fd_sc_hd__tap_1 TAP_5896 (  );
sky130_fd_sc_hd__tap_1 TAP_5897 (  );
sky130_fd_sc_hd__tap_1 TAP_5898 (  );
sky130_fd_sc_hd__tap_1 TAP_5899 (  );
sky130_fd_sc_hd__tap_1 TAP_5900 (  );
sky130_fd_sc_hd__tap_1 TAP_5901 (  );
sky130_fd_sc_hd__tap_1 TAP_5902 (  );
sky130_fd_sc_hd__tap_1 TAP_5903 (  );
sky130_fd_sc_hd__tap_1 TAP_5904 (  );
sky130_fd_sc_hd__tap_1 TAP_5905 (  );
sky130_fd_sc_hd__tap_1 TAP_5906 (  );
sky130_fd_sc_hd__tap_1 TAP_5907 (  );
sky130_fd_sc_hd__tap_1 TAP_5908 (  );
sky130_fd_sc_hd__tap_1 TAP_5909 (  );
sky130_fd_sc_hd__tap_1 TAP_5910 (  );
sky130_fd_sc_hd__tap_1 TAP_5911 (  );
sky130_fd_sc_hd__tap_1 TAP_5912 (  );
sky130_fd_sc_hd__tap_1 TAP_5913 (  );
sky130_fd_sc_hd__tap_1 TAP_5914 (  );
sky130_fd_sc_hd__tap_1 TAP_5915 (  );
sky130_fd_sc_hd__tap_1 TAP_5916 (  );
sky130_fd_sc_hd__tap_1 TAP_5917 (  );
sky130_fd_sc_hd__tap_1 TAP_5918 (  );
sky130_fd_sc_hd__tap_1 TAP_5919 (  );
sky130_fd_sc_hd__tap_1 TAP_5920 (  );
sky130_fd_sc_hd__tap_1 TAP_5921 (  );
sky130_fd_sc_hd__tap_1 TAP_5922 (  );
sky130_fd_sc_hd__tap_1 TAP_5923 (  );
sky130_fd_sc_hd__tap_1 TAP_5924 (  );
sky130_fd_sc_hd__tap_1 TAP_5925 (  );
sky130_fd_sc_hd__tap_1 TAP_5926 (  );
sky130_fd_sc_hd__tap_1 TAP_5927 (  );
sky130_fd_sc_hd__tap_1 TAP_5928 (  );
sky130_fd_sc_hd__tap_1 TAP_5929 (  );
sky130_fd_sc_hd__tap_1 TAP_5930 (  );
sky130_fd_sc_hd__tap_1 TAP_5931 (  );
sky130_fd_sc_hd__tap_1 TAP_5932 (  );
sky130_fd_sc_hd__tap_1 TAP_5933 (  );
sky130_fd_sc_hd__tap_1 TAP_5934 (  );
sky130_fd_sc_hd__tap_1 TAP_5935 (  );
sky130_fd_sc_hd__tap_1 TAP_5936 (  );
sky130_fd_sc_hd__tap_1 TAP_5937 (  );
sky130_fd_sc_hd__tap_1 TAP_5938 (  );
sky130_fd_sc_hd__tap_1 TAP_5939 (  );
sky130_fd_sc_hd__tap_1 TAP_5940 (  );
sky130_fd_sc_hd__tap_1 TAP_5941 (  );
sky130_fd_sc_hd__tap_1 TAP_5942 (  );
sky130_fd_sc_hd__tap_1 TAP_5943 (  );
sky130_fd_sc_hd__tap_1 TAP_5944 (  );
sky130_fd_sc_hd__tap_1 TAP_5945 (  );
sky130_fd_sc_hd__tap_1 TAP_5946 (  );
sky130_fd_sc_hd__tap_1 TAP_5947 (  );
sky130_fd_sc_hd__tap_1 TAP_5948 (  );
sky130_fd_sc_hd__tap_1 TAP_5949 (  );
sky130_fd_sc_hd__tap_1 TAP_5950 (  );
sky130_fd_sc_hd__tap_1 TAP_5951 (  );
sky130_fd_sc_hd__tap_1 TAP_5952 (  );
sky130_fd_sc_hd__tap_1 TAP_5953 (  );
sky130_fd_sc_hd__tap_1 TAP_5954 (  );
sky130_fd_sc_hd__tap_1 TAP_5955 (  );
sky130_fd_sc_hd__tap_1 TAP_5956 (  );
sky130_fd_sc_hd__tap_1 TAP_5957 (  );
sky130_fd_sc_hd__tap_1 TAP_5958 (  );
sky130_fd_sc_hd__tap_1 TAP_5959 (  );
sky130_fd_sc_hd__tap_1 TAP_5960 (  );
sky130_fd_sc_hd__tap_1 TAP_5961 (  );
sky130_fd_sc_hd__tap_1 TAP_5962 (  );
sky130_fd_sc_hd__tap_1 TAP_5963 (  );
sky130_fd_sc_hd__tap_1 TAP_5964 (  );
sky130_fd_sc_hd__tap_1 TAP_5965 (  );
sky130_fd_sc_hd__tap_1 TAP_5966 (  );
sky130_fd_sc_hd__tap_1 TAP_5967 (  );
sky130_fd_sc_hd__tap_1 TAP_5968 (  );
sky130_fd_sc_hd__tap_1 TAP_5969 (  );
sky130_fd_sc_hd__tap_1 TAP_5970 (  );
sky130_fd_sc_hd__tap_1 TAP_5971 (  );
sky130_fd_sc_hd__tap_1 TAP_5972 (  );
sky130_fd_sc_hd__tap_1 TAP_5973 (  );
sky130_fd_sc_hd__tap_1 TAP_5974 (  );
sky130_fd_sc_hd__tap_1 TAP_5975 (  );
sky130_fd_sc_hd__tap_1 TAP_5976 (  );
sky130_fd_sc_hd__tap_1 TAP_5977 (  );
sky130_fd_sc_hd__tap_1 TAP_5978 (  );
sky130_fd_sc_hd__tap_1 TAP_5979 (  );
sky130_fd_sc_hd__tap_1 TAP_5980 (  );
sky130_fd_sc_hd__tap_1 TAP_5981 (  );
sky130_fd_sc_hd__tap_1 TAP_5982 (  );
sky130_fd_sc_hd__tap_1 TAP_5983 (  );
sky130_fd_sc_hd__tap_1 TAP_5984 (  );
sky130_fd_sc_hd__tap_1 TAP_5985 (  );
sky130_fd_sc_hd__tap_1 TAP_5986 (  );
sky130_fd_sc_hd__tap_1 TAP_5987 (  );
sky130_fd_sc_hd__tap_1 TAP_5988 (  );
sky130_fd_sc_hd__tap_1 TAP_5989 (  );
sky130_fd_sc_hd__tap_1 TAP_5990 (  );
sky130_fd_sc_hd__tap_1 TAP_5991 (  );
sky130_fd_sc_hd__tap_1 TAP_5992 (  );
sky130_fd_sc_hd__tap_1 TAP_5993 (  );
sky130_fd_sc_hd__tap_1 TAP_5994 (  );
sky130_fd_sc_hd__tap_1 TAP_5995 (  );
sky130_fd_sc_hd__tap_1 TAP_5996 (  );
sky130_fd_sc_hd__tap_1 TAP_5997 (  );
sky130_fd_sc_hd__tap_1 TAP_5998 (  );
sky130_fd_sc_hd__tap_1 TAP_5999 (  );
sky130_fd_sc_hd__tap_1 TAP_6000 (  );
sky130_fd_sc_hd__tap_1 TAP_6001 (  );
sky130_fd_sc_hd__tap_1 TAP_6002 (  );
sky130_fd_sc_hd__tap_1 TAP_6003 (  );
sky130_fd_sc_hd__tap_1 TAP_6004 (  );
sky130_fd_sc_hd__tap_1 TAP_6005 (  );
sky130_fd_sc_hd__tap_1 TAP_6006 (  );
sky130_fd_sc_hd__tap_1 TAP_6007 (  );
sky130_fd_sc_hd__tap_1 TAP_6008 (  );
sky130_fd_sc_hd__tap_1 TAP_6009 (  );
sky130_fd_sc_hd__tap_1 TAP_6010 (  );
sky130_fd_sc_hd__tap_1 TAP_6011 (  );
sky130_fd_sc_hd__tap_1 TAP_6012 (  );
sky130_fd_sc_hd__tap_1 TAP_6013 (  );
sky130_fd_sc_hd__tap_1 TAP_6014 (  );
sky130_fd_sc_hd__tap_1 TAP_6015 (  );
sky130_fd_sc_hd__tap_1 TAP_6016 (  );
sky130_fd_sc_hd__tap_1 TAP_6017 (  );
sky130_fd_sc_hd__tap_1 TAP_6018 (  );
sky130_fd_sc_hd__tap_1 TAP_6019 (  );
sky130_fd_sc_hd__tap_1 TAP_6020 (  );
sky130_fd_sc_hd__tap_1 TAP_6021 (  );
sky130_fd_sc_hd__tap_1 TAP_6022 (  );
sky130_fd_sc_hd__tap_1 TAP_6023 (  );
sky130_fd_sc_hd__tap_1 TAP_6024 (  );
sky130_fd_sc_hd__tap_1 TAP_6025 (  );
sky130_fd_sc_hd__tap_1 TAP_6026 (  );
sky130_fd_sc_hd__tap_1 TAP_6027 (  );
sky130_fd_sc_hd__tap_1 TAP_6028 (  );
sky130_fd_sc_hd__tap_1 TAP_6029 (  );
sky130_fd_sc_hd__tap_1 TAP_6030 (  );
sky130_fd_sc_hd__tap_1 TAP_6031 (  );
sky130_fd_sc_hd__tap_1 TAP_6032 (  );
sky130_fd_sc_hd__tap_1 TAP_6033 (  );
sky130_fd_sc_hd__tap_1 TAP_6034 (  );
sky130_fd_sc_hd__tap_1 TAP_6035 (  );
sky130_fd_sc_hd__tap_1 TAP_6036 (  );
sky130_fd_sc_hd__tap_1 TAP_6037 (  );
sky130_fd_sc_hd__tap_1 TAP_6038 (  );
sky130_fd_sc_hd__tap_1 TAP_6039 (  );
sky130_fd_sc_hd__tap_1 TAP_6040 (  );
sky130_fd_sc_hd__tap_1 TAP_6041 (  );
sky130_fd_sc_hd__tap_1 TAP_6042 (  );
sky130_fd_sc_hd__tap_1 TAP_6043 (  );
sky130_fd_sc_hd__tap_1 TAP_6044 (  );
sky130_fd_sc_hd__tap_1 TAP_6045 (  );
sky130_fd_sc_hd__tap_1 TAP_6046 (  );
sky130_fd_sc_hd__tap_1 TAP_6047 (  );
sky130_fd_sc_hd__tap_1 TAP_6048 (  );
sky130_fd_sc_hd__tap_1 TAP_6049 (  );
sky130_fd_sc_hd__tap_1 TAP_6050 (  );
sky130_fd_sc_hd__tap_1 TAP_6051 (  );
sky130_fd_sc_hd__tap_1 TAP_6052 (  );
sky130_fd_sc_hd__tap_1 TAP_6053 (  );
sky130_fd_sc_hd__tap_1 TAP_6054 (  );
sky130_fd_sc_hd__tap_1 TAP_6055 (  );
sky130_fd_sc_hd__tap_1 TAP_6056 (  );
sky130_fd_sc_hd__tap_1 TAP_6057 (  );
sky130_fd_sc_hd__tap_1 TAP_6058 (  );
sky130_fd_sc_hd__tap_1 TAP_6059 (  );
sky130_fd_sc_hd__tap_1 TAP_6060 (  );
sky130_fd_sc_hd__tap_1 TAP_6061 (  );
sky130_fd_sc_hd__tap_1 TAP_6062 (  );
sky130_fd_sc_hd__tap_1 TAP_6063 (  );
sky130_fd_sc_hd__tap_1 TAP_6064 (  );
sky130_fd_sc_hd__tap_1 TAP_6065 (  );
sky130_fd_sc_hd__tap_1 TAP_6066 (  );
sky130_fd_sc_hd__tap_1 TAP_6067 (  );
sky130_fd_sc_hd__tap_1 TAP_6068 (  );
sky130_fd_sc_hd__tap_1 TAP_6069 (  );
sky130_fd_sc_hd__tap_1 TAP_6070 (  );
sky130_fd_sc_hd__tap_1 TAP_6071 (  );
sky130_fd_sc_hd__tap_1 TAP_6072 (  );
sky130_fd_sc_hd__tap_1 TAP_6073 (  );
sky130_fd_sc_hd__tap_1 TAP_6074 (  );
sky130_fd_sc_hd__tap_1 TAP_6075 (  );
sky130_fd_sc_hd__tap_1 TAP_6076 (  );
sky130_fd_sc_hd__tap_1 TAP_6077 (  );
sky130_fd_sc_hd__tap_1 TAP_6078 (  );
sky130_fd_sc_hd__tap_1 TAP_6079 (  );
sky130_fd_sc_hd__tap_1 TAP_6080 (  );
sky130_fd_sc_hd__tap_1 TAP_6081 (  );
sky130_fd_sc_hd__tap_1 TAP_6082 (  );
sky130_fd_sc_hd__tap_1 TAP_6083 (  );
sky130_fd_sc_hd__tap_1 TAP_6084 (  );
sky130_fd_sc_hd__tap_1 TAP_6085 (  );
sky130_fd_sc_hd__tap_1 TAP_6086 (  );
sky130_fd_sc_hd__tap_1 TAP_6087 (  );
sky130_fd_sc_hd__tap_1 TAP_6088 (  );
sky130_fd_sc_hd__tap_1 TAP_6089 (  );
sky130_fd_sc_hd__tap_1 TAP_6090 (  );
sky130_fd_sc_hd__tap_1 TAP_6091 (  );
sky130_fd_sc_hd__tap_1 TAP_6092 (  );
sky130_fd_sc_hd__tap_1 TAP_6093 (  );
sky130_fd_sc_hd__tap_1 TAP_6094 (  );
sky130_fd_sc_hd__tap_1 TAP_6095 (  );
sky130_fd_sc_hd__tap_1 TAP_6096 (  );
sky130_fd_sc_hd__tap_1 TAP_6097 (  );
sky130_fd_sc_hd__tap_1 TAP_6098 (  );
sky130_fd_sc_hd__tap_1 TAP_6099 (  );
sky130_fd_sc_hd__tap_1 TAP_6100 (  );
sky130_fd_sc_hd__tap_1 TAP_6101 (  );
sky130_fd_sc_hd__tap_1 TAP_6102 (  );
sky130_fd_sc_hd__tap_1 TAP_6103 (  );
sky130_fd_sc_hd__tap_1 TAP_6104 (  );
sky130_fd_sc_hd__tap_1 TAP_6105 (  );
sky130_fd_sc_hd__tap_1 TAP_6106 (  );
sky130_fd_sc_hd__tap_1 TAP_6107 (  );
sky130_fd_sc_hd__tap_1 TAP_6108 (  );
sky130_fd_sc_hd__tap_1 TAP_6109 (  );
sky130_fd_sc_hd__tap_1 TAP_6110 (  );
sky130_fd_sc_hd__tap_1 TAP_6111 (  );
sky130_fd_sc_hd__tap_1 TAP_6112 (  );
sky130_fd_sc_hd__tap_1 TAP_6113 (  );
sky130_fd_sc_hd__tap_1 TAP_6114 (  );
sky130_fd_sc_hd__tap_1 TAP_6115 (  );
sky130_fd_sc_hd__tap_1 TAP_6116 (  );
sky130_fd_sc_hd__tap_1 TAP_6117 (  );
sky130_fd_sc_hd__tap_1 TAP_6118 (  );
sky130_fd_sc_hd__tap_1 TAP_6119 (  );
sky130_fd_sc_hd__tap_1 TAP_6120 (  );
sky130_fd_sc_hd__tap_1 TAP_6121 (  );
sky130_fd_sc_hd__tap_1 TAP_6122 (  );
sky130_fd_sc_hd__tap_1 TAP_6123 (  );
sky130_fd_sc_hd__tap_1 TAP_6124 (  );
sky130_fd_sc_hd__tap_1 TAP_6125 (  );
sky130_fd_sc_hd__tap_1 TAP_6126 (  );
sky130_fd_sc_hd__tap_1 TAP_6127 (  );
sky130_fd_sc_hd__tap_1 TAP_6128 (  );
sky130_fd_sc_hd__tap_1 TAP_6129 (  );
sky130_fd_sc_hd__tap_1 TAP_6130 (  );
sky130_fd_sc_hd__tap_1 TAP_6131 (  );
sky130_fd_sc_hd__tap_1 TAP_6132 (  );
sky130_fd_sc_hd__tap_1 TAP_6133 (  );
sky130_fd_sc_hd__tap_1 TAP_6134 (  );
sky130_fd_sc_hd__tap_1 TAP_6135 (  );
sky130_fd_sc_hd__tap_1 TAP_6136 (  );
sky130_fd_sc_hd__tap_1 TAP_6137 (  );
sky130_fd_sc_hd__tap_1 TAP_6138 (  );
sky130_fd_sc_hd__tap_1 TAP_6139 (  );
sky130_fd_sc_hd__tap_1 TAP_6140 (  );
sky130_fd_sc_hd__tap_1 TAP_6141 (  );
sky130_fd_sc_hd__tap_1 TAP_6142 (  );
sky130_fd_sc_hd__tap_1 TAP_6143 (  );
sky130_fd_sc_hd__tap_1 TAP_6144 (  );
sky130_fd_sc_hd__tap_1 TAP_6145 (  );
sky130_fd_sc_hd__tap_1 TAP_6146 (  );
sky130_fd_sc_hd__tap_1 TAP_6147 (  );
sky130_fd_sc_hd__tap_1 TAP_6148 (  );
sky130_fd_sc_hd__tap_1 TAP_6149 (  );
sky130_fd_sc_hd__tap_1 TAP_6150 (  );
sky130_fd_sc_hd__tap_1 TAP_6151 (  );
sky130_fd_sc_hd__tap_1 TAP_6152 (  );
sky130_fd_sc_hd__tap_1 TAP_6153 (  );
sky130_fd_sc_hd__tap_1 TAP_6154 (  );
sky130_fd_sc_hd__tap_1 TAP_6155 (  );
sky130_fd_sc_hd__tap_1 TAP_6156 (  );
sky130_fd_sc_hd__tap_1 TAP_6157 (  );
sky130_fd_sc_hd__tap_1 TAP_6158 (  );
sky130_fd_sc_hd__tap_1 TAP_6159 (  );
sky130_fd_sc_hd__tap_1 TAP_6160 (  );
sky130_fd_sc_hd__tap_1 TAP_6161 (  );
sky130_fd_sc_hd__tap_1 TAP_6162 (  );
sky130_fd_sc_hd__tap_1 TAP_6163 (  );
sky130_fd_sc_hd__tap_1 TAP_6164 (  );
sky130_fd_sc_hd__tap_1 TAP_6165 (  );
sky130_fd_sc_hd__tap_1 TAP_6166 (  );
sky130_fd_sc_hd__tap_1 TAP_6167 (  );
sky130_fd_sc_hd__tap_1 TAP_6168 (  );
sky130_fd_sc_hd__tap_1 TAP_6169 (  );
sky130_fd_sc_hd__tap_1 TAP_6170 (  );
sky130_fd_sc_hd__tap_1 TAP_6171 (  );
sky130_fd_sc_hd__tap_1 TAP_6172 (  );
sky130_fd_sc_hd__tap_1 TAP_6173 (  );
sky130_fd_sc_hd__tap_1 TAP_6174 (  );
sky130_fd_sc_hd__tap_1 TAP_6175 (  );
sky130_fd_sc_hd__tap_1 TAP_6176 (  );
sky130_fd_sc_hd__tap_1 TAP_6177 (  );
sky130_fd_sc_hd__tap_1 TAP_6178 (  );
sky130_fd_sc_hd__tap_1 TAP_6179 (  );
sky130_fd_sc_hd__tap_1 TAP_6180 (  );
sky130_fd_sc_hd__tap_1 TAP_6181 (  );
sky130_fd_sc_hd__tap_1 TAP_6182 (  );
sky130_fd_sc_hd__tap_1 TAP_6183 (  );
sky130_fd_sc_hd__tap_1 TAP_6184 (  );
sky130_fd_sc_hd__tap_1 TAP_6185 (  );
sky130_fd_sc_hd__tap_1 TAP_6186 (  );
sky130_fd_sc_hd__tap_1 TAP_6187 (  );
sky130_fd_sc_hd__tap_1 TAP_6188 (  );
sky130_fd_sc_hd__tap_1 TAP_6189 (  );
sky130_fd_sc_hd__tap_1 TAP_6190 (  );
sky130_fd_sc_hd__tap_1 TAP_6191 (  );
sky130_fd_sc_hd__tap_1 TAP_6192 (  );
sky130_fd_sc_hd__tap_1 TAP_6193 (  );
sky130_fd_sc_hd__tap_1 TAP_6194 (  );
sky130_fd_sc_hd__tap_1 TAP_6195 (  );
sky130_fd_sc_hd__tap_1 TAP_6196 (  );
sky130_fd_sc_hd__tap_1 TAP_6197 (  );
sky130_fd_sc_hd__tap_1 TAP_6198 (  );
sky130_fd_sc_hd__tap_1 TAP_6199 (  );
sky130_fd_sc_hd__tap_1 TAP_6200 (  );
sky130_fd_sc_hd__tap_1 TAP_6201 (  );
sky130_fd_sc_hd__tap_1 TAP_6202 (  );
sky130_fd_sc_hd__tap_1 TAP_6203 (  );
sky130_fd_sc_hd__tap_1 TAP_6204 (  );
sky130_fd_sc_hd__tap_1 TAP_6205 (  );
sky130_fd_sc_hd__tap_1 TAP_6206 (  );
sky130_fd_sc_hd__tap_1 TAP_6207 (  );
sky130_fd_sc_hd__tap_1 TAP_6208 (  );
sky130_fd_sc_hd__tap_1 TAP_6209 (  );
sky130_fd_sc_hd__tap_1 TAP_6210 (  );
sky130_fd_sc_hd__tap_1 TAP_6211 (  );
sky130_fd_sc_hd__tap_1 TAP_6212 (  );
sky130_fd_sc_hd__tap_1 TAP_6213 (  );
sky130_fd_sc_hd__tap_1 TAP_6214 (  );
sky130_fd_sc_hd__tap_1 TAP_6215 (  );
sky130_fd_sc_hd__tap_1 TAP_6216 (  );
sky130_fd_sc_hd__tap_1 TAP_6217 (  );
sky130_fd_sc_hd__tap_1 TAP_6218 (  );
sky130_fd_sc_hd__tap_1 TAP_6219 (  );
sky130_fd_sc_hd__tap_1 TAP_6220 (  );
sky130_fd_sc_hd__tap_1 TAP_6221 (  );
sky130_fd_sc_hd__tap_1 TAP_6222 (  );
sky130_fd_sc_hd__tap_1 TAP_6223 (  );
sky130_fd_sc_hd__tap_1 TAP_6224 (  );
sky130_fd_sc_hd__tap_1 TAP_6225 (  );
sky130_fd_sc_hd__tap_1 TAP_6226 (  );
sky130_fd_sc_hd__tap_1 TAP_6227 (  );
sky130_fd_sc_hd__tap_1 TAP_6228 (  );
sky130_fd_sc_hd__tap_1 TAP_6229 (  );
sky130_fd_sc_hd__tap_1 TAP_6230 (  );
sky130_fd_sc_hd__tap_1 TAP_6231 (  );
sky130_fd_sc_hd__tap_1 TAP_6232 (  );
sky130_fd_sc_hd__tap_1 TAP_6233 (  );
sky130_fd_sc_hd__tap_1 TAP_6234 (  );
sky130_fd_sc_hd__tap_1 TAP_6235 (  );
sky130_fd_sc_hd__tap_1 TAP_6236 (  );
sky130_fd_sc_hd__tap_1 TAP_6237 (  );
sky130_fd_sc_hd__tap_1 TAP_6238 (  );
sky130_fd_sc_hd__tap_1 TAP_6239 (  );
sky130_fd_sc_hd__tap_1 TAP_6240 (  );
sky130_fd_sc_hd__tap_1 TAP_6241 (  );
sky130_fd_sc_hd__tap_1 TAP_6242 (  );
sky130_fd_sc_hd__tap_1 TAP_6243 (  );
sky130_fd_sc_hd__tap_1 TAP_6244 (  );
sky130_fd_sc_hd__tap_1 TAP_6245 (  );
sky130_fd_sc_hd__tap_1 TAP_6246 (  );
sky130_fd_sc_hd__tap_1 TAP_6247 (  );
sky130_fd_sc_hd__tap_1 TAP_6248 (  );
sky130_fd_sc_hd__tap_1 TAP_6249 (  );
sky130_fd_sc_hd__tap_1 TAP_6250 (  );
sky130_fd_sc_hd__tap_1 TAP_6251 (  );
sky130_fd_sc_hd__tap_1 TAP_6252 (  );
sky130_fd_sc_hd__tap_1 TAP_6253 (  );
sky130_fd_sc_hd__tap_1 TAP_6254 (  );
sky130_fd_sc_hd__tap_1 TAP_6255 (  );
sky130_fd_sc_hd__tap_1 TAP_6256 (  );
sky130_fd_sc_hd__tap_1 TAP_6257 (  );
sky130_fd_sc_hd__tap_1 TAP_6258 (  );
sky130_fd_sc_hd__tap_1 TAP_6259 (  );
sky130_fd_sc_hd__tap_1 TAP_6260 (  );
sky130_fd_sc_hd__tap_1 TAP_6261 (  );
sky130_fd_sc_hd__tap_1 TAP_6262 (  );
sky130_fd_sc_hd__tap_1 TAP_6263 (  );
sky130_fd_sc_hd__tap_1 TAP_6264 (  );
sky130_fd_sc_hd__tap_1 TAP_6265 (  );
sky130_fd_sc_hd__tap_1 TAP_6266 (  );
sky130_fd_sc_hd__tap_1 TAP_6267 (  );
sky130_fd_sc_hd__tap_1 TAP_6268 (  );
sky130_fd_sc_hd__tap_1 TAP_6269 (  );
sky130_fd_sc_hd__tap_1 TAP_6270 (  );
sky130_fd_sc_hd__tap_1 TAP_6271 (  );
sky130_fd_sc_hd__tap_1 TAP_6272 (  );
sky130_fd_sc_hd__tap_1 TAP_6273 (  );
sky130_fd_sc_hd__tap_1 TAP_6274 (  );
sky130_fd_sc_hd__tap_1 TAP_6275 (  );
sky130_fd_sc_hd__tap_1 TAP_6276 (  );
sky130_fd_sc_hd__tap_1 TAP_6277 (  );
sky130_fd_sc_hd__tap_1 TAP_6278 (  );
sky130_fd_sc_hd__tap_1 TAP_6279 (  );
sky130_fd_sc_hd__tap_1 TAP_6280 (  );
sky130_fd_sc_hd__tap_1 TAP_6281 (  );
sky130_fd_sc_hd__tap_1 TAP_6282 (  );
sky130_fd_sc_hd__tap_1 TAP_6283 (  );
sky130_fd_sc_hd__tap_1 TAP_6284 (  );
sky130_fd_sc_hd__tap_1 TAP_6285 (  );
sky130_fd_sc_hd__tap_1 TAP_6286 (  );
sky130_fd_sc_hd__tap_1 TAP_6287 (  );
sky130_fd_sc_hd__tap_1 TAP_6288 (  );
sky130_fd_sc_hd__tap_1 TAP_6289 (  );
sky130_fd_sc_hd__tap_1 TAP_6290 (  );
sky130_fd_sc_hd__tap_1 TAP_6291 (  );
sky130_fd_sc_hd__tap_1 TAP_6292 (  );
sky130_fd_sc_hd__tap_1 TAP_6293 (  );
sky130_fd_sc_hd__tap_1 TAP_6294 (  );
sky130_fd_sc_hd__tap_1 TAP_6295 (  );
sky130_fd_sc_hd__tap_1 TAP_6296 (  );
sky130_fd_sc_hd__tap_1 TAP_6297 (  );
sky130_fd_sc_hd__tap_1 TAP_6298 (  );
sky130_fd_sc_hd__tap_1 TAP_6299 (  );
sky130_fd_sc_hd__tap_1 TAP_6300 (  );
sky130_fd_sc_hd__tap_1 TAP_6301 (  );
sky130_fd_sc_hd__tap_1 TAP_6302 (  );
sky130_fd_sc_hd__tap_1 TAP_6303 (  );
sky130_fd_sc_hd__tap_1 TAP_6304 (  );
sky130_fd_sc_hd__tap_1 TAP_6305 (  );
sky130_fd_sc_hd__tap_1 TAP_6306 (  );
sky130_fd_sc_hd__tap_1 TAP_6307 (  );
sky130_fd_sc_hd__tap_1 TAP_6308 (  );
sky130_fd_sc_hd__tap_1 TAP_6309 (  );
sky130_fd_sc_hd__tap_1 TAP_6310 (  );
sky130_fd_sc_hd__tap_1 TAP_6311 (  );
sky130_fd_sc_hd__tap_1 TAP_6312 (  );
sky130_fd_sc_hd__tap_1 TAP_6313 (  );
sky130_fd_sc_hd__tap_1 TAP_6314 (  );
sky130_fd_sc_hd__tap_1 TAP_6315 (  );
sky130_fd_sc_hd__tap_1 TAP_6316 (  );
sky130_fd_sc_hd__tap_1 TAP_6317 (  );
sky130_fd_sc_hd__tap_1 TAP_6318 (  );
sky130_fd_sc_hd__tap_1 TAP_6319 (  );
sky130_fd_sc_hd__tap_1 TAP_6320 (  );
sky130_fd_sc_hd__tap_1 TAP_6321 (  );
sky130_fd_sc_hd__tap_1 TAP_6322 (  );
sky130_fd_sc_hd__tap_1 TAP_6323 (  );
sky130_fd_sc_hd__tap_1 TAP_6324 (  );
sky130_fd_sc_hd__tap_1 TAP_6325 (  );
sky130_fd_sc_hd__tap_1 TAP_6326 (  );
sky130_fd_sc_hd__tap_1 TAP_6327 (  );
sky130_fd_sc_hd__tap_1 TAP_6328 (  );
sky130_fd_sc_hd__tap_1 TAP_6329 (  );
sky130_fd_sc_hd__tap_1 TAP_6330 (  );
sky130_fd_sc_hd__tap_1 TAP_6331 (  );
sky130_fd_sc_hd__tap_1 TAP_6332 (  );
sky130_fd_sc_hd__tap_1 TAP_6333 (  );
sky130_fd_sc_hd__tap_1 TAP_6334 (  );
sky130_fd_sc_hd__tap_1 TAP_6335 (  );
sky130_fd_sc_hd__tap_1 TAP_6336 (  );
sky130_fd_sc_hd__tap_1 TAP_6337 (  );
sky130_fd_sc_hd__tap_1 TAP_6338 (  );
sky130_fd_sc_hd__tap_1 TAP_6339 (  );
sky130_fd_sc_hd__tap_1 TAP_6340 (  );
sky130_fd_sc_hd__tap_1 TAP_6341 (  );
sky130_fd_sc_hd__tap_1 TAP_6342 (  );
sky130_fd_sc_hd__tap_1 TAP_6343 (  );
sky130_fd_sc_hd__tap_1 TAP_6344 (  );
sky130_fd_sc_hd__tap_1 TAP_6345 (  );
sky130_fd_sc_hd__tap_1 TAP_6346 (  );
sky130_fd_sc_hd__tap_1 TAP_6347 (  );
sky130_fd_sc_hd__tap_1 TAP_6348 (  );
sky130_fd_sc_hd__tap_1 TAP_6349 (  );
sky130_fd_sc_hd__tap_1 TAP_6350 (  );
sky130_fd_sc_hd__tap_1 TAP_6351 (  );
sky130_fd_sc_hd__tap_1 TAP_6352 (  );
sky130_fd_sc_hd__tap_1 TAP_6353 (  );
sky130_fd_sc_hd__tap_1 TAP_6354 (  );
sky130_fd_sc_hd__tap_1 TAP_6355 (  );
sky130_fd_sc_hd__tap_1 TAP_6356 (  );
sky130_fd_sc_hd__tap_1 TAP_6357 (  );
sky130_fd_sc_hd__tap_1 TAP_6358 (  );
sky130_fd_sc_hd__tap_1 TAP_6359 (  );
sky130_fd_sc_hd__tap_1 TAP_6360 (  );
sky130_fd_sc_hd__tap_1 TAP_6361 (  );
sky130_fd_sc_hd__tap_1 TAP_6362 (  );
sky130_fd_sc_hd__tap_1 TAP_6363 (  );
sky130_fd_sc_hd__tap_1 TAP_6364 (  );
sky130_fd_sc_hd__tap_1 TAP_6365 (  );
sky130_fd_sc_hd__tap_1 TAP_6366 (  );
sky130_fd_sc_hd__tap_1 TAP_6367 (  );
sky130_fd_sc_hd__tap_1 TAP_6368 (  );
sky130_fd_sc_hd__tap_1 TAP_6369 (  );
sky130_fd_sc_hd__tap_1 TAP_6370 (  );
sky130_fd_sc_hd__tap_1 TAP_6371 (  );
sky130_fd_sc_hd__tap_1 TAP_6372 (  );
sky130_fd_sc_hd__tap_1 TAP_6373 (  );
sky130_fd_sc_hd__tap_1 TAP_6374 (  );
sky130_fd_sc_hd__tap_1 TAP_6375 (  );
sky130_fd_sc_hd__tap_1 TAP_6376 (  );
sky130_fd_sc_hd__tap_1 TAP_6377 (  );
sky130_fd_sc_hd__tap_1 TAP_6378 (  );
sky130_fd_sc_hd__tap_1 TAP_6379 (  );
sky130_fd_sc_hd__tap_1 TAP_6380 (  );
sky130_fd_sc_hd__tap_1 TAP_6381 (  );
sky130_fd_sc_hd__tap_1 TAP_6382 (  );
sky130_fd_sc_hd__tap_1 TAP_6383 (  );
sky130_fd_sc_hd__tap_1 TAP_6384 (  );
sky130_fd_sc_hd__tap_1 TAP_6385 (  );
sky130_fd_sc_hd__tap_1 TAP_6386 (  );
sky130_fd_sc_hd__tap_1 TAP_6387 (  );
sky130_fd_sc_hd__tap_1 TAP_6388 (  );
sky130_fd_sc_hd__tap_1 TAP_6389 (  );
sky130_fd_sc_hd__tap_1 TAP_6390 (  );
sky130_fd_sc_hd__tap_1 TAP_6391 (  );
sky130_fd_sc_hd__tap_1 TAP_6392 (  );
sky130_fd_sc_hd__tap_1 TAP_6393 (  );
sky130_fd_sc_hd__tap_1 TAP_6394 (  );
sky130_fd_sc_hd__tap_1 TAP_6395 (  );
sky130_fd_sc_hd__tap_1 TAP_6396 (  );
sky130_fd_sc_hd__tap_1 TAP_6397 (  );
sky130_fd_sc_hd__tap_1 TAP_6398 (  );
sky130_fd_sc_hd__tap_1 TAP_6399 (  );
sky130_fd_sc_hd__tap_1 TAP_6400 (  );
sky130_fd_sc_hd__tap_1 TAP_6401 (  );
sky130_fd_sc_hd__tap_1 TAP_6402 (  );
sky130_fd_sc_hd__tap_1 TAP_6403 (  );
sky130_fd_sc_hd__tap_1 TAP_6404 (  );
sky130_fd_sc_hd__tap_1 TAP_6405 (  );
sky130_fd_sc_hd__tap_1 TAP_6406 (  );
sky130_fd_sc_hd__tap_1 TAP_6407 (  );
sky130_fd_sc_hd__tap_1 TAP_6408 (  );
sky130_fd_sc_hd__tap_1 TAP_6409 (  );
sky130_fd_sc_hd__tap_1 TAP_6410 (  );
sky130_fd_sc_hd__tap_1 TAP_6411 (  );
sky130_fd_sc_hd__tap_1 TAP_6412 (  );
sky130_fd_sc_hd__tap_1 TAP_6413 (  );
sky130_fd_sc_hd__tap_1 TAP_6414 (  );
sky130_fd_sc_hd__tap_1 TAP_6415 (  );
sky130_fd_sc_hd__tap_1 TAP_6416 (  );
sky130_fd_sc_hd__tap_1 TAP_6417 (  );
sky130_fd_sc_hd__tap_1 TAP_6418 (  );
sky130_fd_sc_hd__tap_1 TAP_6419 (  );
sky130_fd_sc_hd__tap_1 TAP_6420 (  );
sky130_fd_sc_hd__tap_1 TAP_6421 (  );
sky130_fd_sc_hd__tap_1 TAP_6422 (  );
sky130_fd_sc_hd__tap_1 TAP_6423 (  );
sky130_fd_sc_hd__tap_1 TAP_6424 (  );
sky130_fd_sc_hd__tap_1 TAP_6425 (  );
sky130_fd_sc_hd__tap_1 TAP_6426 (  );
sky130_fd_sc_hd__tap_1 TAP_6427 (  );
sky130_fd_sc_hd__tap_1 TAP_6428 (  );
sky130_fd_sc_hd__tap_1 TAP_6429 (  );
sky130_fd_sc_hd__tap_1 TAP_6430 (  );
sky130_fd_sc_hd__tap_1 TAP_6431 (  );
sky130_fd_sc_hd__tap_1 TAP_6432 (  );
sky130_fd_sc_hd__tap_1 TAP_6433 (  );
sky130_fd_sc_hd__tap_1 TAP_6434 (  );
sky130_fd_sc_hd__tap_1 TAP_6435 (  );
sky130_fd_sc_hd__tap_1 TAP_6436 (  );
sky130_fd_sc_hd__tap_1 TAP_6437 (  );
sky130_fd_sc_hd__tap_1 TAP_6438 (  );
sky130_fd_sc_hd__tap_1 TAP_6439 (  );
sky130_fd_sc_hd__tap_1 TAP_6440 (  );
sky130_fd_sc_hd__tap_1 TAP_6441 (  );
sky130_fd_sc_hd__tap_1 TAP_6442 (  );
sky130_fd_sc_hd__tap_1 TAP_6443 (  );
sky130_fd_sc_hd__tap_1 TAP_6444 (  );
sky130_fd_sc_hd__tap_1 TAP_6445 (  );
sky130_fd_sc_hd__tap_1 TAP_6446 (  );
sky130_fd_sc_hd__tap_1 TAP_6447 (  );
sky130_fd_sc_hd__tap_1 TAP_6448 (  );
sky130_fd_sc_hd__tap_1 TAP_6449 (  );
sky130_fd_sc_hd__tap_1 TAP_6450 (  );
sky130_fd_sc_hd__tap_1 TAP_6451 (  );
sky130_fd_sc_hd__tap_1 TAP_6452 (  );
sky130_fd_sc_hd__tap_1 TAP_6453 (  );
sky130_fd_sc_hd__tap_1 TAP_6454 (  );
sky130_fd_sc_hd__tap_1 TAP_6455 (  );
sky130_fd_sc_hd__tap_1 TAP_6456 (  );
sky130_fd_sc_hd__tap_1 TAP_6457 (  );
sky130_fd_sc_hd__tap_1 TAP_6458 (  );
sky130_fd_sc_hd__tap_1 TAP_6459 (  );
sky130_fd_sc_hd__tap_1 TAP_6460 (  );
sky130_fd_sc_hd__tap_1 TAP_6461 (  );
sky130_fd_sc_hd__tap_1 TAP_6462 (  );
sky130_fd_sc_hd__tap_1 TAP_6463 (  );
sky130_fd_sc_hd__tap_1 TAP_6464 (  );
sky130_fd_sc_hd__tap_1 TAP_6465 (  );
sky130_fd_sc_hd__tap_1 TAP_6466 (  );
sky130_fd_sc_hd__tap_1 TAP_6467 (  );
sky130_fd_sc_hd__tap_1 TAP_6468 (  );
sky130_fd_sc_hd__tap_1 TAP_6469 (  );
sky130_fd_sc_hd__tap_1 TAP_6470 (  );
sky130_fd_sc_hd__tap_1 TAP_6471 (  );
sky130_fd_sc_hd__tap_1 TAP_6472 (  );
sky130_fd_sc_hd__tap_1 TAP_6473 (  );
sky130_fd_sc_hd__tap_1 TAP_6474 (  );
sky130_fd_sc_hd__tap_1 TAP_6475 (  );
sky130_fd_sc_hd__tap_1 TAP_6476 (  );
sky130_fd_sc_hd__tap_1 TAP_6477 (  );
sky130_fd_sc_hd__tap_1 TAP_6478 (  );
sky130_fd_sc_hd__tap_1 TAP_6479 (  );
sky130_fd_sc_hd__tap_1 TAP_6480 (  );
sky130_fd_sc_hd__tap_1 TAP_6481 (  );
sky130_fd_sc_hd__tap_1 TAP_6482 (  );
sky130_fd_sc_hd__tap_1 TAP_6483 (  );
sky130_fd_sc_hd__tap_1 TAP_6484 (  );
sky130_fd_sc_hd__tap_1 TAP_6485 (  );
sky130_fd_sc_hd__tap_1 TAP_6486 (  );
sky130_fd_sc_hd__tap_1 TAP_6487 (  );
sky130_fd_sc_hd__tap_1 TAP_6488 (  );
sky130_fd_sc_hd__tap_1 TAP_6489 (  );
sky130_fd_sc_hd__tap_1 TAP_6490 (  );
sky130_fd_sc_hd__tap_1 TAP_6491 (  );
sky130_fd_sc_hd__tap_1 TAP_6492 (  );
sky130_fd_sc_hd__tap_1 TAP_6493 (  );
sky130_fd_sc_hd__tap_1 TAP_6494 (  );
sky130_fd_sc_hd__tap_1 TAP_6495 (  );
sky130_fd_sc_hd__tap_1 TAP_6496 (  );
sky130_fd_sc_hd__tap_1 TAP_6497 (  );
sky130_fd_sc_hd__tap_1 TAP_6498 (  );
sky130_fd_sc_hd__tap_1 TAP_6499 (  );
sky130_fd_sc_hd__tap_1 TAP_6500 (  );
sky130_fd_sc_hd__tap_1 TAP_6501 (  );
sky130_fd_sc_hd__tap_1 TAP_6502 (  );
sky130_fd_sc_hd__tap_1 TAP_6503 (  );
sky130_fd_sc_hd__tap_1 TAP_6504 (  );
sky130_fd_sc_hd__tap_1 TAP_6505 (  );
sky130_fd_sc_hd__tap_1 TAP_6506 (  );
sky130_fd_sc_hd__tap_1 TAP_6507 (  );
sky130_fd_sc_hd__tap_1 TAP_6508 (  );
sky130_fd_sc_hd__tap_1 TAP_6509 (  );
sky130_fd_sc_hd__tap_1 TAP_6510 (  );
sky130_fd_sc_hd__tap_1 TAP_6511 (  );
sky130_fd_sc_hd__tap_1 TAP_6512 (  );
sky130_fd_sc_hd__tap_1 TAP_6513 (  );
sky130_fd_sc_hd__tap_1 TAP_6514 (  );
sky130_fd_sc_hd__tap_1 TAP_6515 (  );
sky130_fd_sc_hd__tap_1 TAP_6516 (  );
sky130_fd_sc_hd__tap_1 TAP_6517 (  );
sky130_fd_sc_hd__tap_1 TAP_6518 (  );
sky130_fd_sc_hd__tap_1 TAP_6519 (  );
sky130_fd_sc_hd__tap_1 TAP_6520 (  );
sky130_fd_sc_hd__tap_1 TAP_6521 (  );
sky130_fd_sc_hd__tap_1 TAP_6522 (  );
sky130_fd_sc_hd__tap_1 TAP_6523 (  );
sky130_fd_sc_hd__tap_1 TAP_6524 (  );
sky130_fd_sc_hd__tap_1 TAP_6525 (  );
sky130_fd_sc_hd__tap_1 TAP_6526 (  );
sky130_fd_sc_hd__tap_1 TAP_6527 (  );
sky130_fd_sc_hd__tap_1 TAP_6528 (  );
sky130_fd_sc_hd__tap_1 TAP_6529 (  );
sky130_fd_sc_hd__tap_1 TAP_6530 (  );
sky130_fd_sc_hd__tap_1 TAP_6531 (  );
sky130_fd_sc_hd__tap_1 TAP_6532 (  );
sky130_fd_sc_hd__tap_1 TAP_6533 (  );
sky130_fd_sc_hd__tap_1 TAP_6534 (  );
sky130_fd_sc_hd__tap_1 TAP_6535 (  );
sky130_fd_sc_hd__tap_1 TAP_6536 (  );
sky130_fd_sc_hd__tap_1 TAP_6537 (  );
sky130_fd_sc_hd__tap_1 TAP_6538 (  );
sky130_fd_sc_hd__tap_1 TAP_6539 (  );
sky130_fd_sc_hd__tap_1 TAP_6540 (  );
sky130_fd_sc_hd__tap_1 TAP_6541 (  );
sky130_fd_sc_hd__tap_1 TAP_6542 (  );
sky130_fd_sc_hd__tap_1 TAP_6543 (  );
sky130_fd_sc_hd__tap_1 TAP_6544 (  );
sky130_fd_sc_hd__tap_1 TAP_6545 (  );
sky130_fd_sc_hd__tap_1 TAP_6546 (  );
sky130_fd_sc_hd__tap_1 TAP_6547 (  );
sky130_fd_sc_hd__tap_1 TAP_6548 (  );
sky130_fd_sc_hd__tap_1 TAP_6549 (  );
sky130_fd_sc_hd__tap_1 TAP_6550 (  );
sky130_fd_sc_hd__tap_1 TAP_6551 (  );
sky130_fd_sc_hd__tap_1 TAP_6552 (  );
sky130_fd_sc_hd__tap_1 TAP_6553 (  );
sky130_fd_sc_hd__tap_1 TAP_6554 (  );
sky130_fd_sc_hd__tap_1 TAP_6555 (  );
sky130_fd_sc_hd__tap_1 TAP_6556 (  );
sky130_fd_sc_hd__tap_1 TAP_6557 (  );
sky130_fd_sc_hd__tap_1 TAP_6558 (  );
sky130_fd_sc_hd__tap_1 TAP_6559 (  );
sky130_fd_sc_hd__tap_1 TAP_6560 (  );
sky130_fd_sc_hd__tap_1 TAP_6561 (  );
sky130_fd_sc_hd__tap_1 TAP_6562 (  );
sky130_fd_sc_hd__tap_1 TAP_6563 (  );
sky130_fd_sc_hd__tap_1 TAP_6564 (  );
sky130_fd_sc_hd__tap_1 TAP_6565 (  );
sky130_fd_sc_hd__tap_1 TAP_6566 (  );
sky130_fd_sc_hd__tap_1 TAP_6567 (  );
sky130_fd_sc_hd__tap_1 TAP_6568 (  );
sky130_fd_sc_hd__tap_1 TAP_6569 (  );
sky130_fd_sc_hd__tap_1 TAP_6570 (  );
sky130_fd_sc_hd__tap_1 TAP_6571 (  );
sky130_fd_sc_hd__tap_1 TAP_6572 (  );
sky130_fd_sc_hd__tap_1 TAP_6573 (  );
sky130_fd_sc_hd__tap_1 TAP_6574 (  );
sky130_fd_sc_hd__tap_1 TAP_6575 (  );
sky130_fd_sc_hd__tap_1 TAP_6576 (  );
sky130_fd_sc_hd__tap_1 TAP_6577 (  );
sky130_fd_sc_hd__tap_1 TAP_6578 (  );
sky130_fd_sc_hd__tap_1 TAP_6579 (  );
sky130_fd_sc_hd__tap_1 TAP_6580 (  );
sky130_fd_sc_hd__tap_1 TAP_6581 (  );
sky130_fd_sc_hd__tap_1 TAP_6582 (  );
sky130_fd_sc_hd__tap_1 TAP_6583 (  );
sky130_fd_sc_hd__tap_1 TAP_6584 (  );
sky130_fd_sc_hd__tap_1 TAP_6585 (  );
sky130_fd_sc_hd__tap_1 TAP_6586 (  );
sky130_fd_sc_hd__tap_1 TAP_6587 (  );
sky130_fd_sc_hd__tap_1 TAP_6588 (  );
sky130_fd_sc_hd__tap_1 TAP_6589 (  );
sky130_fd_sc_hd__tap_1 TAP_6590 (  );
sky130_fd_sc_hd__tap_1 TAP_6591 (  );
sky130_fd_sc_hd__tap_1 TAP_6592 (  );
sky130_fd_sc_hd__tap_1 TAP_6593 (  );
sky130_fd_sc_hd__tap_1 TAP_6594 (  );
sky130_fd_sc_hd__tap_1 TAP_6595 (  );
sky130_fd_sc_hd__tap_1 TAP_6596 (  );
sky130_fd_sc_hd__tap_1 TAP_6597 (  );
sky130_fd_sc_hd__tap_1 TAP_6598 (  );
sky130_fd_sc_hd__tap_1 TAP_6599 (  );
sky130_fd_sc_hd__tap_1 TAP_6600 (  );
sky130_fd_sc_hd__tap_1 TAP_6601 (  );
sky130_fd_sc_hd__tap_1 TAP_6602 (  );
sky130_fd_sc_hd__tap_1 TAP_6603 (  );
sky130_fd_sc_hd__tap_1 TAP_6604 (  );
sky130_fd_sc_hd__tap_1 TAP_6605 (  );
sky130_fd_sc_hd__tap_1 TAP_6606 (  );
sky130_fd_sc_hd__tap_1 TAP_6607 (  );
sky130_fd_sc_hd__tap_1 TAP_6608 (  );
sky130_fd_sc_hd__tap_1 TAP_6609 (  );
sky130_fd_sc_hd__tap_1 TAP_6610 (  );
sky130_fd_sc_hd__tap_1 TAP_6611 (  );
sky130_fd_sc_hd__tap_1 TAP_6612 (  );
sky130_fd_sc_hd__tap_1 TAP_6613 (  );
sky130_fd_sc_hd__tap_1 TAP_6614 (  );
sky130_fd_sc_hd__tap_1 TAP_6615 (  );
sky130_fd_sc_hd__tap_1 TAP_6616 (  );
sky130_fd_sc_hd__tap_1 TAP_6617 (  );
sky130_fd_sc_hd__tap_1 TAP_6618 (  );
sky130_fd_sc_hd__tap_1 TAP_6619 (  );
sky130_fd_sc_hd__tap_1 TAP_6620 (  );
sky130_fd_sc_hd__tap_1 TAP_6621 (  );
sky130_fd_sc_hd__tap_1 TAP_6622 (  );
sky130_fd_sc_hd__tap_1 TAP_6623 (  );
sky130_fd_sc_hd__tap_1 TAP_6624 (  );
sky130_fd_sc_hd__tap_1 TAP_6625 (  );
sky130_fd_sc_hd__tap_1 TAP_6626 (  );
sky130_fd_sc_hd__tap_1 TAP_6627 (  );
sky130_fd_sc_hd__tap_1 TAP_6628 (  );
sky130_fd_sc_hd__tap_1 TAP_6629 (  );
sky130_fd_sc_hd__tap_1 TAP_6630 (  );
sky130_fd_sc_hd__tap_1 TAP_6631 (  );
sky130_fd_sc_hd__tap_1 TAP_6632 (  );
sky130_fd_sc_hd__tap_1 TAP_6633 (  );
sky130_fd_sc_hd__tap_1 TAP_6634 (  );
sky130_fd_sc_hd__tap_1 TAP_6635 (  );
sky130_fd_sc_hd__tap_1 TAP_6636 (  );
sky130_fd_sc_hd__tap_1 TAP_6637 (  );
sky130_fd_sc_hd__tap_1 TAP_6638 (  );
sky130_fd_sc_hd__tap_1 TAP_6639 (  );
sky130_fd_sc_hd__tap_1 TAP_6640 (  );
sky130_fd_sc_hd__tap_1 TAP_6641 (  );
sky130_fd_sc_hd__tap_1 TAP_6642 (  );
sky130_fd_sc_hd__tap_1 TAP_6643 (  );
sky130_fd_sc_hd__tap_1 TAP_6644 (  );
sky130_fd_sc_hd__tap_1 TAP_6645 (  );
sky130_fd_sc_hd__tap_1 TAP_6646 (  );
sky130_fd_sc_hd__tap_1 TAP_6647 (  );
sky130_fd_sc_hd__tap_1 TAP_6648 (  );
sky130_fd_sc_hd__tap_1 TAP_6649 (  );
sky130_fd_sc_hd__tap_1 TAP_6650 (  );
sky130_fd_sc_hd__tap_1 TAP_6651 (  );
sky130_fd_sc_hd__tap_1 TAP_6652 (  );
sky130_fd_sc_hd__tap_1 TAP_6653 (  );
sky130_fd_sc_hd__tap_1 TAP_6654 (  );
sky130_fd_sc_hd__tap_1 TAP_6655 (  );
sky130_fd_sc_hd__tap_1 TAP_6656 (  );
sky130_fd_sc_hd__tap_1 TAP_6657 (  );
sky130_fd_sc_hd__tap_1 TAP_6658 (  );
sky130_fd_sc_hd__tap_1 TAP_6659 (  );
sky130_fd_sc_hd__tap_1 TAP_6660 (  );
sky130_fd_sc_hd__tap_1 TAP_6661 (  );
sky130_fd_sc_hd__tap_1 TAP_6662 (  );
sky130_fd_sc_hd__tap_1 TAP_6663 (  );
sky130_fd_sc_hd__tap_1 TAP_6664 (  );
sky130_fd_sc_hd__tap_1 TAP_6665 (  );
sky130_fd_sc_hd__tap_1 TAP_6666 (  );
sky130_fd_sc_hd__tap_1 TAP_6667 (  );
sky130_fd_sc_hd__tap_1 TAP_6668 (  );
sky130_fd_sc_hd__tap_1 TAP_6669 (  );
sky130_fd_sc_hd__tap_1 TAP_6670 (  );
sky130_fd_sc_hd__tap_1 TAP_6671 (  );
sky130_fd_sc_hd__tap_1 TAP_6672 (  );
sky130_fd_sc_hd__tap_1 TAP_6673 (  );
sky130_fd_sc_hd__tap_1 TAP_6674 (  );
sky130_fd_sc_hd__tap_1 TAP_6675 (  );
sky130_fd_sc_hd__tap_1 TAP_6676 (  );
sky130_fd_sc_hd__tap_1 TAP_6677 (  );
sky130_fd_sc_hd__tap_1 TAP_6678 (  );
sky130_fd_sc_hd__tap_1 TAP_6679 (  );
sky130_fd_sc_hd__tap_1 TAP_6680 (  );
sky130_fd_sc_hd__tap_1 TAP_6681 (  );
sky130_fd_sc_hd__tap_1 TAP_6682 (  );
sky130_fd_sc_hd__tap_1 TAP_6683 (  );
sky130_fd_sc_hd__tap_1 TAP_6684 (  );
sky130_fd_sc_hd__tap_1 TAP_6685 (  );
sky130_fd_sc_hd__tap_1 TAP_6686 (  );
sky130_fd_sc_hd__tap_1 TAP_6687 (  );
sky130_fd_sc_hd__tap_1 TAP_6688 (  );
sky130_fd_sc_hd__tap_1 TAP_6689 (  );
sky130_fd_sc_hd__tap_1 TAP_6690 (  );
sky130_fd_sc_hd__tap_1 TAP_6691 (  );
sky130_fd_sc_hd__tap_1 TAP_6692 (  );
sky130_fd_sc_hd__tap_1 TAP_6693 (  );
sky130_fd_sc_hd__tap_1 TAP_6694 (  );
sky130_fd_sc_hd__tap_1 TAP_6695 (  );
sky130_fd_sc_hd__tap_1 TAP_6696 (  );
sky130_fd_sc_hd__tap_1 TAP_6697 (  );
sky130_fd_sc_hd__tap_1 TAP_6698 (  );
sky130_fd_sc_hd__tap_1 TAP_6699 (  );
sky130_fd_sc_hd__tap_1 TAP_6700 (  );
sky130_fd_sc_hd__tap_1 TAP_6701 (  );
sky130_fd_sc_hd__tap_1 TAP_6702 (  );
sky130_fd_sc_hd__tap_1 TAP_6703 (  );
sky130_fd_sc_hd__tap_1 TAP_6704 (  );
sky130_fd_sc_hd__tap_1 TAP_6705 (  );
sky130_fd_sc_hd__tap_1 TAP_6706 (  );
sky130_fd_sc_hd__tap_1 TAP_6707 (  );
sky130_fd_sc_hd__tap_1 TAP_6708 (  );
sky130_fd_sc_hd__tap_1 TAP_6709 (  );
sky130_fd_sc_hd__tap_1 TAP_6710 (  );
sky130_fd_sc_hd__tap_1 TAP_6711 (  );
sky130_fd_sc_hd__tap_1 TAP_6712 (  );
sky130_fd_sc_hd__tap_1 TAP_6713 (  );
sky130_fd_sc_hd__tap_1 TAP_6714 (  );
sky130_fd_sc_hd__tap_1 TAP_6715 (  );
sky130_fd_sc_hd__tap_1 TAP_6716 (  );
sky130_fd_sc_hd__tap_1 TAP_6717 (  );
sky130_fd_sc_hd__tap_1 TAP_6718 (  );
sky130_fd_sc_hd__tap_1 TAP_6719 (  );
sky130_fd_sc_hd__tap_1 TAP_6720 (  );
sky130_fd_sc_hd__tap_1 TAP_6721 (  );
sky130_fd_sc_hd__tap_1 TAP_6722 (  );
sky130_fd_sc_hd__tap_1 TAP_6723 (  );
sky130_fd_sc_hd__tap_1 TAP_6724 (  );
sky130_fd_sc_hd__tap_1 TAP_6725 (  );
sky130_fd_sc_hd__tap_1 TAP_6726 (  );
sky130_fd_sc_hd__tap_1 TAP_6727 (  );
sky130_fd_sc_hd__tap_1 TAP_6728 (  );
sky130_fd_sc_hd__tap_1 TAP_6729 (  );
sky130_fd_sc_hd__tap_1 TAP_6730 (  );
sky130_fd_sc_hd__tap_1 TAP_6731 (  );
sky130_fd_sc_hd__tap_1 TAP_6732 (  );
sky130_fd_sc_hd__tap_1 TAP_6733 (  );
sky130_fd_sc_hd__tap_1 TAP_6734 (  );
sky130_fd_sc_hd__tap_1 TAP_6735 (  );
sky130_fd_sc_hd__tap_1 TAP_6736 (  );
sky130_fd_sc_hd__tap_1 TAP_6737 (  );
sky130_fd_sc_hd__tap_1 TAP_6738 (  );
sky130_fd_sc_hd__tap_1 TAP_6739 (  );
sky130_fd_sc_hd__tap_1 TAP_6740 (  );
sky130_fd_sc_hd__tap_1 TAP_6741 (  );
sky130_fd_sc_hd__tap_1 TAP_6742 (  );
sky130_fd_sc_hd__tap_1 TAP_6743 (  );
sky130_fd_sc_hd__tap_1 TAP_6744 (  );
sky130_fd_sc_hd__tap_1 TAP_6745 (  );
sky130_fd_sc_hd__tap_1 TAP_6746 (  );
sky130_fd_sc_hd__tap_1 TAP_6747 (  );
sky130_fd_sc_hd__tap_1 TAP_6748 (  );
sky130_fd_sc_hd__tap_1 TAP_6749 (  );
sky130_fd_sc_hd__tap_1 TAP_6750 (  );
sky130_fd_sc_hd__tap_1 TAP_6751 (  );
sky130_fd_sc_hd__tap_1 TAP_6752 (  );
sky130_fd_sc_hd__tap_1 TAP_6753 (  );
sky130_fd_sc_hd__tap_1 TAP_6754 (  );
sky130_fd_sc_hd__tap_1 TAP_6755 (  );
sky130_fd_sc_hd__tap_1 TAP_6756 (  );
sky130_fd_sc_hd__tap_1 TAP_6757 (  );
sky130_fd_sc_hd__tap_1 TAP_6758 (  );
sky130_fd_sc_hd__tap_1 TAP_6759 (  );
sky130_fd_sc_hd__tap_1 TAP_6760 (  );
sky130_fd_sc_hd__tap_1 TAP_6761 (  );
sky130_fd_sc_hd__tap_1 TAP_6762 (  );
sky130_fd_sc_hd__tap_1 TAP_6763 (  );
sky130_fd_sc_hd__tap_1 TAP_6764 (  );
sky130_fd_sc_hd__tap_1 TAP_6765 (  );
sky130_fd_sc_hd__tap_1 TAP_6766 (  );
sky130_fd_sc_hd__tap_1 TAP_6767 (  );
sky130_fd_sc_hd__tap_1 TAP_6768 (  );
sky130_fd_sc_hd__tap_1 TAP_6769 (  );
sky130_fd_sc_hd__tap_1 TAP_6770 (  );
sky130_fd_sc_hd__tap_1 TAP_6771 (  );
sky130_fd_sc_hd__tap_1 TAP_6772 (  );
sky130_fd_sc_hd__tap_1 TAP_6773 (  );
sky130_fd_sc_hd__tap_1 TAP_6774 (  );
sky130_fd_sc_hd__tap_1 TAP_6775 (  );
sky130_fd_sc_hd__tap_1 TAP_6776 (  );
sky130_fd_sc_hd__tap_1 TAP_6777 (  );
sky130_fd_sc_hd__tap_1 TAP_6778 (  );
sky130_fd_sc_hd__tap_1 TAP_6779 (  );
sky130_fd_sc_hd__tap_1 TAP_6780 (  );
sky130_fd_sc_hd__tap_1 TAP_6781 (  );
sky130_fd_sc_hd__tap_1 TAP_6782 (  );
sky130_fd_sc_hd__tap_1 TAP_6783 (  );
sky130_fd_sc_hd__tap_1 TAP_6784 (  );
sky130_fd_sc_hd__tap_1 TAP_6785 (  );
sky130_fd_sc_hd__tap_1 TAP_6786 (  );
sky130_fd_sc_hd__tap_1 TAP_6787 (  );
sky130_fd_sc_hd__tap_1 TAP_6788 (  );
sky130_fd_sc_hd__tap_1 TAP_6789 (  );
sky130_fd_sc_hd__tap_1 TAP_6790 (  );
sky130_fd_sc_hd__tap_1 TAP_6791 (  );
sky130_fd_sc_hd__tap_1 TAP_6792 (  );
sky130_fd_sc_hd__tap_1 TAP_6793 (  );
sky130_fd_sc_hd__tap_1 TAP_6794 (  );
sky130_fd_sc_hd__tap_1 TAP_6795 (  );
sky130_fd_sc_hd__tap_1 TAP_6796 (  );
sky130_fd_sc_hd__tap_1 TAP_6797 (  );
sky130_fd_sc_hd__tap_1 TAP_6798 (  );
sky130_fd_sc_hd__tap_1 TAP_6799 (  );
sky130_fd_sc_hd__tap_1 TAP_6800 (  );
sky130_fd_sc_hd__tap_1 TAP_6801 (  );
sky130_fd_sc_hd__tap_1 TAP_6802 (  );
sky130_fd_sc_hd__tap_1 TAP_6803 (  );
sky130_fd_sc_hd__tap_1 TAP_6804 (  );
sky130_fd_sc_hd__tap_1 TAP_6805 (  );
sky130_fd_sc_hd__tap_1 TAP_6806 (  );
sky130_fd_sc_hd__tap_1 TAP_6807 (  );
sky130_fd_sc_hd__tap_1 TAP_6808 (  );
sky130_fd_sc_hd__tap_1 TAP_6809 (  );
sky130_fd_sc_hd__tap_1 TAP_6810 (  );
sky130_fd_sc_hd__tap_1 TAP_6811 (  );
sky130_fd_sc_hd__tap_1 TAP_6812 (  );
sky130_fd_sc_hd__tap_1 TAP_6813 (  );
sky130_fd_sc_hd__tap_1 TAP_6814 (  );
sky130_fd_sc_hd__tap_1 TAP_6815 (  );
sky130_fd_sc_hd__tap_1 TAP_6816 (  );
sky130_fd_sc_hd__tap_1 TAP_6817 (  );
sky130_fd_sc_hd__tap_1 TAP_6818 (  );
sky130_fd_sc_hd__tap_1 TAP_6819 (  );
sky130_fd_sc_hd__tap_1 TAP_6820 (  );
sky130_fd_sc_hd__tap_1 TAP_6821 (  );
sky130_fd_sc_hd__tap_1 TAP_6822 (  );
sky130_fd_sc_hd__tap_1 TAP_6823 (  );
sky130_fd_sc_hd__tap_1 TAP_6824 (  );
sky130_fd_sc_hd__tap_1 TAP_6825 (  );
sky130_fd_sc_hd__tap_1 TAP_6826 (  );
sky130_fd_sc_hd__tap_1 TAP_6827 (  );
sky130_fd_sc_hd__tap_1 TAP_6828 (  );
sky130_fd_sc_hd__tap_1 TAP_6829 (  );
sky130_fd_sc_hd__tap_1 TAP_6830 (  );
sky130_fd_sc_hd__tap_1 TAP_6831 (  );
sky130_fd_sc_hd__tap_1 TAP_6832 (  );
sky130_fd_sc_hd__tap_1 TAP_6833 (  );
sky130_fd_sc_hd__tap_1 TAP_6834 (  );
sky130_fd_sc_hd__tap_1 TAP_6835 (  );
sky130_fd_sc_hd__tap_1 TAP_6836 (  );
sky130_fd_sc_hd__tap_1 TAP_6837 (  );
sky130_fd_sc_hd__tap_1 TAP_6838 (  );
sky130_fd_sc_hd__tap_1 TAP_6839 (  );
sky130_fd_sc_hd__tap_1 TAP_6840 (  );
sky130_fd_sc_hd__tap_1 TAP_6841 (  );
sky130_fd_sc_hd__tap_1 TAP_6842 (  );
sky130_fd_sc_hd__tap_1 TAP_6843 (  );
sky130_fd_sc_hd__tap_1 TAP_6844 (  );
sky130_fd_sc_hd__tap_1 TAP_6845 (  );
sky130_fd_sc_hd__tap_1 TAP_6846 (  );
sky130_fd_sc_hd__tap_1 TAP_6847 (  );
sky130_fd_sc_hd__tap_1 TAP_6848 (  );
sky130_fd_sc_hd__tap_1 TAP_6849 (  );
sky130_fd_sc_hd__tap_1 TAP_6850 (  );
sky130_fd_sc_hd__tap_1 TAP_6851 (  );
sky130_fd_sc_hd__tap_1 TAP_6852 (  );
sky130_fd_sc_hd__tap_1 TAP_6853 (  );
sky130_fd_sc_hd__tap_1 TAP_6854 (  );
sky130_fd_sc_hd__tap_1 TAP_6855 (  );
sky130_fd_sc_hd__tap_1 TAP_6856 (  );
sky130_fd_sc_hd__tap_1 TAP_6857 (  );
sky130_fd_sc_hd__tap_1 TAP_6858 (  );
sky130_fd_sc_hd__tap_1 TAP_6859 (  );
sky130_fd_sc_hd__tap_1 TAP_6860 (  );
sky130_fd_sc_hd__tap_1 TAP_6861 (  );
sky130_fd_sc_hd__tap_1 TAP_6862 (  );
sky130_fd_sc_hd__tap_1 TAP_6863 (  );
sky130_fd_sc_hd__tap_1 TAP_6864 (  );
sky130_fd_sc_hd__tap_1 TAP_6865 (  );
sky130_fd_sc_hd__tap_1 TAP_6866 (  );
sky130_fd_sc_hd__tap_1 TAP_6867 (  );
sky130_fd_sc_hd__tap_1 TAP_6868 (  );
sky130_fd_sc_hd__tap_1 TAP_6869 (  );
sky130_fd_sc_hd__tap_1 TAP_6870 (  );
sky130_fd_sc_hd__tap_1 TAP_6871 (  );
sky130_fd_sc_hd__tap_1 TAP_6872 (  );
sky130_fd_sc_hd__tap_1 TAP_6873 (  );
sky130_fd_sc_hd__tap_1 TAP_6874 (  );
sky130_fd_sc_hd__tap_1 TAP_6875 (  );
sky130_fd_sc_hd__tap_1 TAP_6876 (  );
sky130_fd_sc_hd__tap_1 TAP_6877 (  );
sky130_fd_sc_hd__tap_1 TAP_6878 (  );
sky130_fd_sc_hd__tap_1 TAP_6879 (  );
sky130_fd_sc_hd__tap_1 TAP_6880 (  );
sky130_fd_sc_hd__tap_1 TAP_6881 (  );
sky130_fd_sc_hd__tap_1 TAP_6882 (  );
sky130_fd_sc_hd__tap_1 TAP_6883 (  );
sky130_fd_sc_hd__tap_1 TAP_6884 (  );
sky130_fd_sc_hd__tap_1 TAP_6885 (  );
sky130_fd_sc_hd__tap_1 TAP_6886 (  );
sky130_fd_sc_hd__tap_1 TAP_6887 (  );
sky130_fd_sc_hd__tap_1 TAP_6888 (  );
sky130_fd_sc_hd__tap_1 TAP_6889 (  );
sky130_fd_sc_hd__tap_1 TAP_6890 (  );
sky130_fd_sc_hd__tap_1 TAP_6891 (  );
sky130_fd_sc_hd__tap_1 TAP_6892 (  );
sky130_fd_sc_hd__tap_1 TAP_6893 (  );
sky130_fd_sc_hd__tap_1 TAP_6894 (  );
sky130_fd_sc_hd__tap_1 TAP_6895 (  );
sky130_fd_sc_hd__tap_1 TAP_6896 (  );
sky130_fd_sc_hd__tap_1 TAP_6897 (  );
sky130_fd_sc_hd__tap_1 TAP_6898 (  );
sky130_fd_sc_hd__tap_1 TAP_6899 (  );
sky130_fd_sc_hd__tap_1 TAP_6900 (  );
sky130_fd_sc_hd__tap_1 TAP_6901 (  );
sky130_fd_sc_hd__tap_1 TAP_6902 (  );
sky130_fd_sc_hd__tap_1 TAP_6903 (  );
sky130_fd_sc_hd__tap_1 TAP_6904 (  );
sky130_fd_sc_hd__tap_1 TAP_6905 (  );
sky130_fd_sc_hd__tap_1 TAP_6906 (  );
sky130_fd_sc_hd__tap_1 TAP_6907 (  );
sky130_fd_sc_hd__tap_1 TAP_6908 (  );
sky130_fd_sc_hd__tap_1 TAP_6909 (  );
sky130_fd_sc_hd__tap_1 TAP_6910 (  );
sky130_fd_sc_hd__tap_1 TAP_6911 (  );
sky130_fd_sc_hd__tap_1 TAP_6912 (  );
sky130_fd_sc_hd__tap_1 TAP_6913 (  );
sky130_fd_sc_hd__tap_1 TAP_6914 (  );
sky130_fd_sc_hd__tap_1 TAP_6915 (  );
sky130_fd_sc_hd__tap_1 TAP_6916 (  );
sky130_fd_sc_hd__tap_1 TAP_6917 (  );
sky130_fd_sc_hd__tap_1 TAP_6918 (  );
sky130_fd_sc_hd__tap_1 TAP_6919 (  );
sky130_fd_sc_hd__tap_1 TAP_6920 (  );
sky130_fd_sc_hd__tap_1 TAP_6921 (  );
sky130_fd_sc_hd__tap_1 TAP_6922 (  );
sky130_fd_sc_hd__tap_1 TAP_6923 (  );
sky130_fd_sc_hd__tap_1 TAP_6924 (  );
sky130_fd_sc_hd__tap_1 TAP_6925 (  );
sky130_fd_sc_hd__tap_1 TAP_6926 (  );
sky130_fd_sc_hd__tap_1 TAP_6927 (  );
sky130_fd_sc_hd__tap_1 TAP_6928 (  );
sky130_fd_sc_hd__tap_1 TAP_6929 (  );
sky130_fd_sc_hd__tap_1 TAP_6930 (  );
sky130_fd_sc_hd__tap_1 TAP_6931 (  );
sky130_fd_sc_hd__tap_1 TAP_6932 (  );
sky130_fd_sc_hd__tap_1 TAP_6933 (  );
sky130_fd_sc_hd__tap_1 TAP_6934 (  );
sky130_fd_sc_hd__tap_1 TAP_6935 (  );
sky130_fd_sc_hd__tap_1 TAP_6936 (  );
sky130_fd_sc_hd__tap_1 TAP_6937 (  );
sky130_fd_sc_hd__tap_1 TAP_6938 (  );
sky130_fd_sc_hd__tap_1 TAP_6939 (  );
sky130_fd_sc_hd__tap_1 TAP_6940 (  );
sky130_fd_sc_hd__tap_1 TAP_6941 (  );
sky130_fd_sc_hd__tap_1 TAP_6942 (  );
sky130_fd_sc_hd__tap_1 TAP_6943 (  );
sky130_fd_sc_hd__tap_1 TAP_6944 (  );
sky130_fd_sc_hd__tap_1 TAP_6945 (  );
sky130_fd_sc_hd__tap_1 TAP_6946 (  );
sky130_fd_sc_hd__tap_1 TAP_6947 (  );
sky130_fd_sc_hd__tap_1 TAP_6948 (  );
sky130_fd_sc_hd__tap_1 TAP_6949 (  );
sky130_fd_sc_hd__tap_1 TAP_6950 (  );
sky130_fd_sc_hd__tap_1 TAP_6951 (  );
sky130_fd_sc_hd__tap_1 TAP_6952 (  );
sky130_fd_sc_hd__tap_1 TAP_6953 (  );
sky130_fd_sc_hd__tap_1 TAP_6954 (  );
sky130_fd_sc_hd__tap_1 TAP_6955 (  );
sky130_fd_sc_hd__tap_1 TAP_6956 (  );
sky130_fd_sc_hd__tap_1 TAP_6957 (  );
sky130_fd_sc_hd__tap_1 TAP_6958 (  );
sky130_fd_sc_hd__tap_1 TAP_6959 (  );
sky130_fd_sc_hd__tap_1 TAP_6960 (  );
sky130_fd_sc_hd__tap_1 TAP_6961 (  );
sky130_fd_sc_hd__tap_1 TAP_6962 (  );
sky130_fd_sc_hd__tap_1 TAP_6963 (  );
sky130_fd_sc_hd__tap_1 TAP_6964 (  );
sky130_fd_sc_hd__tap_1 TAP_6965 (  );
sky130_fd_sc_hd__tap_1 TAP_6966 (  );
sky130_fd_sc_hd__tap_1 TAP_6967 (  );
sky130_fd_sc_hd__tap_1 TAP_6968 (  );
sky130_fd_sc_hd__tap_1 TAP_6969 (  );
sky130_fd_sc_hd__tap_1 TAP_6970 (  );
sky130_fd_sc_hd__tap_1 TAP_6971 (  );
sky130_fd_sc_hd__tap_1 TAP_6972 (  );
sky130_fd_sc_hd__tap_1 TAP_6973 (  );
sky130_fd_sc_hd__tap_1 TAP_6974 (  );
sky130_fd_sc_hd__tap_1 TAP_6975 (  );
sky130_fd_sc_hd__tap_1 TAP_6976 (  );
sky130_fd_sc_hd__tap_1 TAP_6977 (  );
sky130_fd_sc_hd__tap_1 TAP_6978 (  );
sky130_fd_sc_hd__tap_1 TAP_6979 (  );
sky130_fd_sc_hd__tap_1 TAP_6980 (  );
sky130_fd_sc_hd__tap_1 TAP_6981 (  );
sky130_fd_sc_hd__tap_1 TAP_6982 (  );
sky130_fd_sc_hd__tap_1 TAP_6983 (  );
sky130_fd_sc_hd__tap_1 TAP_6984 (  );
sky130_fd_sc_hd__tap_1 TAP_6985 (  );
sky130_fd_sc_hd__tap_1 TAP_6986 (  );
sky130_fd_sc_hd__tap_1 TAP_6987 (  );
sky130_fd_sc_hd__tap_1 TAP_6988 (  );
sky130_fd_sc_hd__tap_1 TAP_6989 (  );
sky130_fd_sc_hd__tap_1 TAP_6990 (  );
sky130_fd_sc_hd__tap_1 TAP_6991 (  );
sky130_fd_sc_hd__tap_1 TAP_6992 (  );
sky130_fd_sc_hd__tap_1 TAP_6993 (  );
sky130_fd_sc_hd__tap_1 TAP_6994 (  );
sky130_fd_sc_hd__tap_1 TAP_6995 (  );
sky130_fd_sc_hd__tap_1 TAP_6996 (  );
sky130_fd_sc_hd__tap_1 TAP_6997 (  );
sky130_fd_sc_hd__tap_1 TAP_6998 (  );
sky130_fd_sc_hd__tap_1 TAP_6999 (  );
sky130_fd_sc_hd__tap_1 TAP_7000 (  );
sky130_fd_sc_hd__tap_1 TAP_7001 (  );
sky130_fd_sc_hd__tap_1 TAP_7002 (  );
sky130_fd_sc_hd__tap_1 TAP_7003 (  );
sky130_fd_sc_hd__tap_1 TAP_7004 (  );
sky130_fd_sc_hd__tap_1 TAP_7005 (  );
sky130_fd_sc_hd__tap_1 TAP_7006 (  );
sky130_fd_sc_hd__tap_1 TAP_7007 (  );
sky130_fd_sc_hd__tap_1 TAP_7008 (  );
sky130_fd_sc_hd__tap_1 TAP_7009 (  );
sky130_fd_sc_hd__tap_1 TAP_7010 (  );
sky130_fd_sc_hd__tap_1 TAP_7011 (  );
sky130_fd_sc_hd__tap_1 TAP_7012 (  );
sky130_fd_sc_hd__tap_1 TAP_7013 (  );
sky130_fd_sc_hd__tap_1 TAP_7014 (  );
sky130_fd_sc_hd__tap_1 TAP_7015 (  );
sky130_fd_sc_hd__tap_1 TAP_7016 (  );
sky130_fd_sc_hd__tap_1 TAP_7017 (  );
sky130_fd_sc_hd__tap_1 TAP_7018 (  );
sky130_fd_sc_hd__tap_1 TAP_7019 (  );
sky130_fd_sc_hd__tap_1 TAP_7020 (  );
sky130_fd_sc_hd__tap_1 TAP_7021 (  );
sky130_fd_sc_hd__tap_1 TAP_7022 (  );
sky130_fd_sc_hd__tap_1 TAP_7023 (  );
sky130_fd_sc_hd__tap_1 TAP_7024 (  );
sky130_fd_sc_hd__tap_1 TAP_7025 (  );
sky130_fd_sc_hd__tap_1 TAP_7026 (  );
sky130_fd_sc_hd__tap_1 TAP_7027 (  );
sky130_fd_sc_hd__tap_1 TAP_7028 (  );
sky130_fd_sc_hd__tap_1 TAP_7029 (  );
sky130_fd_sc_hd__tap_1 TAP_7030 (  );
sky130_fd_sc_hd__tap_1 TAP_7031 (  );
sky130_fd_sc_hd__tap_1 TAP_7032 (  );
sky130_fd_sc_hd__tap_1 TAP_7033 (  );
sky130_fd_sc_hd__tap_1 TAP_7034 (  );
sky130_fd_sc_hd__tap_1 TAP_7035 (  );
sky130_fd_sc_hd__tap_1 TAP_7036 (  );
sky130_fd_sc_hd__tap_1 TAP_7037 (  );
sky130_fd_sc_hd__tap_1 TAP_7038 (  );
sky130_fd_sc_hd__tap_1 TAP_7039 (  );
sky130_fd_sc_hd__tap_1 TAP_7040 (  );
sky130_fd_sc_hd__tap_1 TAP_7041 (  );
sky130_fd_sc_hd__tap_1 TAP_7042 (  );
sky130_fd_sc_hd__tap_1 TAP_7043 (  );
sky130_fd_sc_hd__tap_1 TAP_7044 (  );
sky130_fd_sc_hd__tap_1 TAP_7045 (  );
sky130_fd_sc_hd__tap_1 TAP_7046 (  );
sky130_fd_sc_hd__tap_1 TAP_7047 (  );
sky130_fd_sc_hd__tap_1 TAP_7048 (  );
sky130_fd_sc_hd__tap_1 TAP_7049 (  );
sky130_fd_sc_hd__tap_1 TAP_7050 (  );
sky130_fd_sc_hd__tap_1 TAP_7051 (  );
sky130_fd_sc_hd__tap_1 TAP_7052 (  );
sky130_fd_sc_hd__tap_1 TAP_7053 (  );
sky130_fd_sc_hd__tap_1 TAP_7054 (  );
sky130_fd_sc_hd__tap_1 TAP_7055 (  );
sky130_fd_sc_hd__tap_1 TAP_7056 (  );
sky130_fd_sc_hd__tap_1 TAP_7057 (  );
sky130_fd_sc_hd__tap_1 TAP_7058 (  );
sky130_fd_sc_hd__tap_1 TAP_7059 (  );
sky130_fd_sc_hd__tap_1 TAP_7060 (  );
sky130_fd_sc_hd__tap_1 TAP_7061 (  );
sky130_fd_sc_hd__tap_1 TAP_7062 (  );
sky130_fd_sc_hd__tap_1 TAP_7063 (  );
sky130_fd_sc_hd__tap_1 TAP_7064 (  );
sky130_fd_sc_hd__tap_1 TAP_7065 (  );
sky130_fd_sc_hd__tap_1 TAP_7066 (  );
sky130_fd_sc_hd__tap_1 TAP_7067 (  );
sky130_fd_sc_hd__tap_1 TAP_7068 (  );
sky130_fd_sc_hd__tap_1 TAP_7069 (  );
sky130_fd_sc_hd__tap_1 TAP_7070 (  );
sky130_fd_sc_hd__tap_1 TAP_7071 (  );
sky130_fd_sc_hd__tap_1 TAP_7072 (  );
sky130_fd_sc_hd__tap_1 TAP_7073 (  );
sky130_fd_sc_hd__tap_1 TAP_7074 (  );
sky130_fd_sc_hd__tap_1 TAP_7075 (  );
sky130_fd_sc_hd__tap_1 TAP_7076 (  );
sky130_fd_sc_hd__tap_1 TAP_7077 (  );
sky130_fd_sc_hd__tap_1 TAP_7078 (  );
sky130_fd_sc_hd__tap_1 TAP_7079 (  );
sky130_fd_sc_hd__tap_1 TAP_7080 (  );
sky130_fd_sc_hd__tap_1 TAP_7081 (  );
sky130_fd_sc_hd__tap_1 TAP_7082 (  );
sky130_fd_sc_hd__tap_1 TAP_7083 (  );
sky130_fd_sc_hd__tap_1 TAP_7084 (  );
sky130_fd_sc_hd__tap_1 TAP_7085 (  );
sky130_fd_sc_hd__tap_1 TAP_7086 (  );
sky130_fd_sc_hd__tap_1 TAP_7087 (  );
sky130_fd_sc_hd__tap_1 TAP_7088 (  );
sky130_fd_sc_hd__tap_1 TAP_7089 (  );
sky130_fd_sc_hd__tap_1 TAP_7090 (  );
sky130_fd_sc_hd__tap_1 TAP_7091 (  );
sky130_fd_sc_hd__tap_1 TAP_7092 (  );
sky130_fd_sc_hd__tap_1 TAP_7093 (  );
sky130_fd_sc_hd__tap_1 TAP_7094 (  );
sky130_fd_sc_hd__tap_1 TAP_7095 (  );
sky130_fd_sc_hd__tap_1 TAP_7096 (  );
sky130_fd_sc_hd__tap_1 TAP_7097 (  );
sky130_fd_sc_hd__tap_1 TAP_7098 (  );
sky130_fd_sc_hd__tap_1 TAP_7099 (  );
sky130_fd_sc_hd__tap_1 TAP_7100 (  );
sky130_fd_sc_hd__tap_1 TAP_7101 (  );
sky130_fd_sc_hd__tap_1 TAP_7102 (  );
sky130_fd_sc_hd__tap_1 TAP_7103 (  );
sky130_fd_sc_hd__tap_1 TAP_7104 (  );
sky130_fd_sc_hd__tap_1 TAP_7105 (  );
sky130_fd_sc_hd__tap_1 TAP_7106 (  );
sky130_fd_sc_hd__tap_1 TAP_7107 (  );
sky130_fd_sc_hd__tap_1 TAP_7108 (  );
sky130_fd_sc_hd__tap_1 TAP_7109 (  );
sky130_fd_sc_hd__tap_1 TAP_7110 (  );
sky130_fd_sc_hd__tap_1 TAP_7111 (  );
sky130_fd_sc_hd__tap_1 TAP_7112 (  );
sky130_fd_sc_hd__tap_1 TAP_7113 (  );
sky130_fd_sc_hd__tap_1 TAP_7114 (  );
sky130_fd_sc_hd__tap_1 TAP_7115 (  );
sky130_fd_sc_hd__tap_1 TAP_7116 (  );
sky130_fd_sc_hd__tap_1 TAP_7117 (  );
sky130_fd_sc_hd__tap_1 TAP_7118 (  );
sky130_fd_sc_hd__tap_1 TAP_7119 (  );
sky130_fd_sc_hd__tap_1 TAP_7120 (  );
sky130_fd_sc_hd__tap_1 TAP_7121 (  );
sky130_fd_sc_hd__tap_1 TAP_7122 (  );
sky130_fd_sc_hd__tap_1 TAP_7123 (  );
sky130_fd_sc_hd__tap_1 TAP_7124 (  );
sky130_fd_sc_hd__tap_1 TAP_7125 (  );
sky130_fd_sc_hd__tap_1 TAP_7126 (  );
sky130_fd_sc_hd__tap_1 TAP_7127 (  );
sky130_fd_sc_hd__tap_1 TAP_7128 (  );
sky130_fd_sc_hd__tap_1 TAP_7129 (  );
sky130_fd_sc_hd__tap_1 TAP_7130 (  );
sky130_fd_sc_hd__tap_1 TAP_7131 (  );
sky130_fd_sc_hd__tap_1 TAP_7132 (  );
sky130_fd_sc_hd__tap_1 TAP_7133 (  );
sky130_fd_sc_hd__tap_1 TAP_7134 (  );
sky130_fd_sc_hd__tap_1 TAP_7135 (  );
sky130_fd_sc_hd__tap_1 TAP_7136 (  );
sky130_fd_sc_hd__tap_1 TAP_7137 (  );
sky130_fd_sc_hd__tap_1 TAP_7138 (  );
sky130_fd_sc_hd__tap_1 TAP_7139 (  );
sky130_fd_sc_hd__tap_1 TAP_7140 (  );
sky130_fd_sc_hd__tap_1 TAP_7141 (  );
sky130_fd_sc_hd__tap_1 TAP_7142 (  );
sky130_fd_sc_hd__tap_1 TAP_7143 (  );
sky130_fd_sc_hd__tap_1 TAP_7144 (  );
sky130_fd_sc_hd__tap_1 TAP_7145 (  );
sky130_fd_sc_hd__tap_1 TAP_7146 (  );
sky130_fd_sc_hd__tap_1 TAP_7147 (  );
sky130_fd_sc_hd__tap_1 TAP_7148 (  );
sky130_fd_sc_hd__tap_1 TAP_7149 (  );
sky130_fd_sc_hd__tap_1 TAP_7150 (  );
sky130_fd_sc_hd__tap_1 TAP_7151 (  );
sky130_fd_sc_hd__tap_1 TAP_7152 (  );
sky130_fd_sc_hd__tap_1 TAP_7153 (  );
sky130_fd_sc_hd__tap_1 TAP_7154 (  );
sky130_fd_sc_hd__tap_1 TAP_7155 (  );
sky130_fd_sc_hd__tap_1 TAP_7156 (  );
sky130_fd_sc_hd__tap_1 TAP_7157 (  );
sky130_fd_sc_hd__tap_1 TAP_7158 (  );
sky130_fd_sc_hd__tap_1 TAP_7159 (  );
sky130_fd_sc_hd__tap_1 TAP_7160 (  );
sky130_fd_sc_hd__tap_1 TAP_7161 (  );
sky130_fd_sc_hd__tap_1 TAP_7162 (  );
sky130_fd_sc_hd__tap_1 TAP_7163 (  );
sky130_fd_sc_hd__tap_1 TAP_7164 (  );
sky130_fd_sc_hd__tap_1 TAP_7165 (  );
sky130_fd_sc_hd__tap_1 TAP_7166 (  );
sky130_fd_sc_hd__tap_1 TAP_7167 (  );
sky130_fd_sc_hd__tap_1 TAP_7168 (  );
sky130_fd_sc_hd__tap_1 TAP_7169 (  );
sky130_fd_sc_hd__tap_1 TAP_7170 (  );
sky130_fd_sc_hd__tap_1 TAP_7171 (  );
sky130_fd_sc_hd__tap_1 TAP_7172 (  );
sky130_fd_sc_hd__tap_1 TAP_7173 (  );
sky130_fd_sc_hd__tap_1 TAP_7174 (  );
sky130_fd_sc_hd__tap_1 TAP_7175 (  );
sky130_fd_sc_hd__tap_1 TAP_7176 (  );
sky130_fd_sc_hd__tap_1 TAP_7177 (  );
sky130_fd_sc_hd__tap_1 TAP_7178 (  );
sky130_fd_sc_hd__tap_1 TAP_7179 (  );
sky130_fd_sc_hd__tap_1 TAP_7180 (  );
sky130_fd_sc_hd__tap_1 TAP_7181 (  );
sky130_fd_sc_hd__tap_1 TAP_7182 (  );
sky130_fd_sc_hd__tap_1 TAP_7183 (  );
sky130_fd_sc_hd__tap_1 TAP_7184 (  );
sky130_fd_sc_hd__tap_1 TAP_7185 (  );
sky130_fd_sc_hd__tap_1 TAP_7186 (  );
sky130_fd_sc_hd__tap_1 TAP_7187 (  );
sky130_fd_sc_hd__tap_1 TAP_7188 (  );
sky130_fd_sc_hd__tap_1 TAP_7189 (  );
sky130_fd_sc_hd__tap_1 TAP_7190 (  );
sky130_fd_sc_hd__tap_1 TAP_7191 (  );
sky130_fd_sc_hd__tap_1 TAP_7192 (  );
sky130_fd_sc_hd__tap_1 TAP_7193 (  );
sky130_fd_sc_hd__tap_1 TAP_7194 (  );
sky130_fd_sc_hd__tap_1 TAP_7195 (  );
sky130_fd_sc_hd__tap_1 TAP_7196 (  );
sky130_fd_sc_hd__tap_1 TAP_7197 (  );
sky130_fd_sc_hd__tap_1 TAP_7198 (  );
sky130_fd_sc_hd__tap_1 TAP_7199 (  );
sky130_fd_sc_hd__tap_1 TAP_7200 (  );
sky130_fd_sc_hd__tap_1 TAP_7201 (  );
sky130_fd_sc_hd__tap_1 TAP_7202 (  );
sky130_fd_sc_hd__tap_1 TAP_7203 (  );
sky130_fd_sc_hd__tap_1 TAP_7204 (  );
sky130_fd_sc_hd__tap_1 TAP_7205 (  );
sky130_fd_sc_hd__tap_1 TAP_7206 (  );
sky130_fd_sc_hd__tap_1 TAP_7207 (  );
sky130_fd_sc_hd__tap_1 TAP_7208 (  );
sky130_fd_sc_hd__tap_1 TAP_7209 (  );
sky130_fd_sc_hd__tap_1 TAP_7210 (  );
sky130_fd_sc_hd__tap_1 TAP_7211 (  );
sky130_fd_sc_hd__tap_1 TAP_7212 (  );
sky130_fd_sc_hd__tap_1 TAP_7213 (  );
sky130_fd_sc_hd__tap_1 TAP_7214 (  );
sky130_fd_sc_hd__tap_1 TAP_7215 (  );
sky130_fd_sc_hd__tap_1 TAP_7216 (  );
sky130_fd_sc_hd__tap_1 TAP_7217 (  );
sky130_fd_sc_hd__tap_1 TAP_7218 (  );
sky130_fd_sc_hd__tap_1 TAP_7219 (  );
sky130_fd_sc_hd__tap_1 TAP_7220 (  );
sky130_fd_sc_hd__tap_1 TAP_7221 (  );
sky130_fd_sc_hd__tap_1 TAP_7222 (  );
sky130_fd_sc_hd__tap_1 TAP_7223 (  );
sky130_fd_sc_hd__tap_1 TAP_7224 (  );
sky130_fd_sc_hd__tap_1 TAP_7225 (  );
sky130_fd_sc_hd__tap_1 TAP_7226 (  );
sky130_fd_sc_hd__tap_1 TAP_7227 (  );
sky130_fd_sc_hd__tap_1 TAP_7228 (  );
sky130_fd_sc_hd__tap_1 TAP_7229 (  );
sky130_fd_sc_hd__tap_1 TAP_7230 (  );
sky130_fd_sc_hd__tap_1 TAP_7231 (  );
sky130_fd_sc_hd__tap_1 TAP_7232 (  );
sky130_fd_sc_hd__tap_1 TAP_7233 (  );
sky130_fd_sc_hd__tap_1 TAP_7234 (  );
sky130_fd_sc_hd__tap_1 TAP_7235 (  );
sky130_fd_sc_hd__tap_1 TAP_7236 (  );
sky130_fd_sc_hd__tap_1 TAP_7237 (  );
sky130_fd_sc_hd__tap_1 TAP_7238 (  );
sky130_fd_sc_hd__tap_1 TAP_7239 (  );
sky130_fd_sc_hd__tap_1 TAP_7240 (  );
sky130_fd_sc_hd__tap_1 TAP_7241 (  );
sky130_fd_sc_hd__tap_1 TAP_7242 (  );
sky130_fd_sc_hd__tap_1 TAP_7243 (  );
sky130_fd_sc_hd__tap_1 TAP_7244 (  );
sky130_fd_sc_hd__tap_1 TAP_7245 (  );
sky130_fd_sc_hd__tap_1 TAP_7246 (  );
sky130_fd_sc_hd__tap_1 TAP_7247 (  );
sky130_fd_sc_hd__tap_1 TAP_7248 (  );
sky130_fd_sc_hd__tap_1 TAP_7249 (  );
sky130_fd_sc_hd__tap_1 TAP_7250 (  );
sky130_fd_sc_hd__tap_1 TAP_7251 (  );
sky130_fd_sc_hd__tap_1 TAP_7252 (  );
sky130_fd_sc_hd__tap_1 TAP_7253 (  );
sky130_fd_sc_hd__tap_1 TAP_7254 (  );
sky130_fd_sc_hd__tap_1 TAP_7255 (  );
sky130_fd_sc_hd__tap_1 TAP_7256 (  );
sky130_fd_sc_hd__tap_1 TAP_7257 (  );
sky130_fd_sc_hd__tap_1 TAP_7258 (  );
sky130_fd_sc_hd__tap_1 TAP_7259 (  );
sky130_fd_sc_hd__tap_1 TAP_7260 (  );
sky130_fd_sc_hd__tap_1 TAP_7261 (  );
sky130_fd_sc_hd__tap_1 TAP_7262 (  );
sky130_fd_sc_hd__tap_1 TAP_7263 (  );
sky130_fd_sc_hd__tap_1 TAP_7264 (  );
sky130_fd_sc_hd__tap_1 TAP_7265 (  );
sky130_fd_sc_hd__tap_1 TAP_7266 (  );
sky130_fd_sc_hd__tap_1 TAP_7267 (  );
sky130_fd_sc_hd__tap_1 TAP_7268 (  );
sky130_fd_sc_hd__tap_1 TAP_7269 (  );
sky130_fd_sc_hd__tap_1 TAP_7270 (  );
sky130_fd_sc_hd__tap_1 TAP_7271 (  );
sky130_fd_sc_hd__tap_1 TAP_7272 (  );
sky130_fd_sc_hd__tap_1 TAP_7273 (  );
sky130_fd_sc_hd__tap_1 TAP_7274 (  );
sky130_fd_sc_hd__tap_1 TAP_7275 (  );
sky130_fd_sc_hd__tap_1 TAP_7276 (  );
sky130_fd_sc_hd__tap_1 TAP_7277 (  );
sky130_fd_sc_hd__tap_1 TAP_7278 (  );
sky130_fd_sc_hd__tap_1 TAP_7279 (  );
sky130_fd_sc_hd__tap_1 TAP_7280 (  );
sky130_fd_sc_hd__tap_1 TAP_7281 (  );
sky130_fd_sc_hd__tap_1 TAP_7282 (  );
sky130_fd_sc_hd__tap_1 TAP_7283 (  );
sky130_fd_sc_hd__tap_1 TAP_7284 (  );
sky130_fd_sc_hd__tap_1 TAP_7285 (  );
sky130_fd_sc_hd__tap_1 TAP_7286 (  );
sky130_fd_sc_hd__tap_1 TAP_7287 (  );
sky130_fd_sc_hd__tap_1 TAP_7288 (  );
sky130_fd_sc_hd__tap_1 TAP_7289 (  );
sky130_fd_sc_hd__tap_1 TAP_7290 (  );
sky130_fd_sc_hd__tap_1 TAP_7291 (  );
sky130_fd_sc_hd__tap_1 TAP_7292 (  );
sky130_fd_sc_hd__tap_1 TAP_7293 (  );
sky130_fd_sc_hd__tap_1 TAP_7294 (  );
sky130_fd_sc_hd__tap_1 TAP_7295 (  );
sky130_fd_sc_hd__tap_1 TAP_7296 (  );
sky130_fd_sc_hd__tap_1 TAP_7297 (  );
sky130_fd_sc_hd__tap_1 TAP_7298 (  );
sky130_fd_sc_hd__tap_1 TAP_7299 (  );
sky130_fd_sc_hd__tap_1 TAP_7300 (  );
sky130_fd_sc_hd__tap_1 TAP_7301 (  );
sky130_fd_sc_hd__tap_1 TAP_7302 (  );
sky130_fd_sc_hd__tap_1 TAP_7303 (  );
sky130_fd_sc_hd__tap_1 TAP_7304 (  );
sky130_fd_sc_hd__tap_1 TAP_7305 (  );
sky130_fd_sc_hd__tap_1 TAP_7306 (  );
sky130_fd_sc_hd__tap_1 TAP_7307 (  );
sky130_fd_sc_hd__tap_1 TAP_7308 (  );
sky130_fd_sc_hd__tap_1 TAP_7309 (  );
sky130_fd_sc_hd__tap_1 TAP_7310 (  );
sky130_fd_sc_hd__tap_1 TAP_7311 (  );
sky130_fd_sc_hd__tap_1 TAP_7312 (  );
sky130_fd_sc_hd__tap_1 TAP_7313 (  );
sky130_fd_sc_hd__tap_1 TAP_7314 (  );
sky130_fd_sc_hd__tap_1 TAP_7315 (  );
sky130_fd_sc_hd__tap_1 TAP_7316 (  );
sky130_fd_sc_hd__tap_1 TAP_7317 (  );
sky130_fd_sc_hd__tap_1 TAP_7318 (  );
sky130_fd_sc_hd__tap_1 TAP_7319 (  );
sky130_fd_sc_hd__tap_1 TAP_7320 (  );
sky130_fd_sc_hd__tap_1 TAP_7321 (  );
sky130_fd_sc_hd__tap_1 TAP_7322 (  );
sky130_fd_sc_hd__tap_1 TAP_7323 (  );
sky130_fd_sc_hd__tap_1 TAP_7324 (  );
sky130_fd_sc_hd__tap_1 TAP_7325 (  );
sky130_fd_sc_hd__tap_1 TAP_7326 (  );
sky130_fd_sc_hd__tap_1 TAP_7327 (  );
sky130_fd_sc_hd__tap_1 TAP_7328 (  );
sky130_fd_sc_hd__tap_1 TAP_7329 (  );
sky130_fd_sc_hd__tap_1 TAP_7330 (  );
sky130_fd_sc_hd__tap_1 TAP_7331 (  );
sky130_fd_sc_hd__tap_1 TAP_7332 (  );
sky130_fd_sc_hd__tap_1 TAP_7333 (  );
sky130_fd_sc_hd__tap_1 TAP_7334 (  );
sky130_fd_sc_hd__tap_1 TAP_7335 (  );
sky130_fd_sc_hd__tap_1 TAP_7336 (  );
sky130_fd_sc_hd__tap_1 TAP_7337 (  );
sky130_fd_sc_hd__tap_1 TAP_7338 (  );
sky130_fd_sc_hd__tap_1 TAP_7339 (  );
sky130_fd_sc_hd__tap_1 TAP_734 (  );
sky130_fd_sc_hd__tap_1 TAP_7340 (  );
sky130_fd_sc_hd__tap_1 TAP_7341 (  );
sky130_fd_sc_hd__tap_1 TAP_7342 (  );
sky130_fd_sc_hd__tap_1 TAP_7343 (  );
sky130_fd_sc_hd__tap_1 TAP_7344 (  );
sky130_fd_sc_hd__tap_1 TAP_7345 (  );
sky130_fd_sc_hd__tap_1 TAP_7346 (  );
sky130_fd_sc_hd__tap_1 TAP_7347 (  );
sky130_fd_sc_hd__tap_1 TAP_7348 (  );
sky130_fd_sc_hd__tap_1 TAP_7349 (  );
sky130_fd_sc_hd__tap_1 TAP_735 (  );
sky130_fd_sc_hd__tap_1 TAP_7350 (  );
sky130_fd_sc_hd__tap_1 TAP_7351 (  );
sky130_fd_sc_hd__tap_1 TAP_7352 (  );
sky130_fd_sc_hd__tap_1 TAP_7353 (  );
sky130_fd_sc_hd__tap_1 TAP_7354 (  );
sky130_fd_sc_hd__tap_1 TAP_7355 (  );
sky130_fd_sc_hd__tap_1 TAP_7356 (  );
sky130_fd_sc_hd__tap_1 TAP_7357 (  );
sky130_fd_sc_hd__tap_1 TAP_7358 (  );
sky130_fd_sc_hd__tap_1 TAP_7359 (  );
sky130_fd_sc_hd__tap_1 TAP_736 (  );
sky130_fd_sc_hd__tap_1 TAP_7360 (  );
sky130_fd_sc_hd__tap_1 TAP_7361 (  );
sky130_fd_sc_hd__tap_1 TAP_7362 (  );
sky130_fd_sc_hd__tap_1 TAP_7363 (  );
sky130_fd_sc_hd__tap_1 TAP_7364 (  );
sky130_fd_sc_hd__tap_1 TAP_7365 (  );
sky130_fd_sc_hd__tap_1 TAP_7366 (  );
sky130_fd_sc_hd__tap_1 TAP_7367 (  );
sky130_fd_sc_hd__tap_1 TAP_7368 (  );
sky130_fd_sc_hd__tap_1 TAP_7369 (  );
sky130_fd_sc_hd__tap_1 TAP_737 (  );
sky130_fd_sc_hd__tap_1 TAP_7370 (  );
sky130_fd_sc_hd__tap_1 TAP_7371 (  );
sky130_fd_sc_hd__tap_1 TAP_7372 (  );
sky130_fd_sc_hd__tap_1 TAP_7373 (  );
sky130_fd_sc_hd__tap_1 TAP_7374 (  );
sky130_fd_sc_hd__tap_1 TAP_7375 (  );
sky130_fd_sc_hd__tap_1 TAP_7376 (  );
sky130_fd_sc_hd__tap_1 TAP_7377 (  );
sky130_fd_sc_hd__tap_1 TAP_7378 (  );
sky130_fd_sc_hd__tap_1 TAP_7379 (  );
sky130_fd_sc_hd__tap_1 TAP_738 (  );
sky130_fd_sc_hd__tap_1 TAP_7380 (  );
sky130_fd_sc_hd__tap_1 TAP_7381 (  );
sky130_fd_sc_hd__tap_1 TAP_7382 (  );
sky130_fd_sc_hd__tap_1 TAP_7383 (  );
sky130_fd_sc_hd__tap_1 TAP_7384 (  );
sky130_fd_sc_hd__tap_1 TAP_7385 (  );
sky130_fd_sc_hd__tap_1 TAP_7386 (  );
sky130_fd_sc_hd__tap_1 TAP_7387 (  );
sky130_fd_sc_hd__tap_1 TAP_7388 (  );
sky130_fd_sc_hd__tap_1 TAP_7389 (  );
sky130_fd_sc_hd__tap_1 TAP_739 (  );
sky130_fd_sc_hd__tap_1 TAP_7390 (  );
sky130_fd_sc_hd__tap_1 TAP_7391 (  );
sky130_fd_sc_hd__tap_1 TAP_7392 (  );
sky130_fd_sc_hd__tap_1 TAP_7393 (  );
sky130_fd_sc_hd__tap_1 TAP_7394 (  );
sky130_fd_sc_hd__tap_1 TAP_7395 (  );
sky130_fd_sc_hd__tap_1 TAP_7396 (  );
sky130_fd_sc_hd__tap_1 TAP_7397 (  );
sky130_fd_sc_hd__tap_1 TAP_7398 (  );
sky130_fd_sc_hd__tap_1 TAP_7399 (  );
sky130_fd_sc_hd__tap_1 TAP_740 (  );
sky130_fd_sc_hd__tap_1 TAP_7400 (  );
sky130_fd_sc_hd__tap_1 TAP_7401 (  );
sky130_fd_sc_hd__tap_1 TAP_7402 (  );
sky130_fd_sc_hd__tap_1 TAP_7403 (  );
sky130_fd_sc_hd__tap_1 TAP_7404 (  );
sky130_fd_sc_hd__tap_1 TAP_7405 (  );
sky130_fd_sc_hd__tap_1 TAP_7406 (  );
sky130_fd_sc_hd__tap_1 TAP_7407 (  );
sky130_fd_sc_hd__tap_1 TAP_7408 (  );
sky130_fd_sc_hd__tap_1 TAP_7409 (  );
sky130_fd_sc_hd__tap_1 TAP_741 (  );
sky130_fd_sc_hd__tap_1 TAP_7410 (  );
sky130_fd_sc_hd__tap_1 TAP_7411 (  );
sky130_fd_sc_hd__tap_1 TAP_7412 (  );
sky130_fd_sc_hd__tap_1 TAP_7413 (  );
sky130_fd_sc_hd__tap_1 TAP_7414 (  );
sky130_fd_sc_hd__tap_1 TAP_7415 (  );
sky130_fd_sc_hd__tap_1 TAP_7416 (  );
sky130_fd_sc_hd__tap_1 TAP_7417 (  );
sky130_fd_sc_hd__tap_1 TAP_7418 (  );
sky130_fd_sc_hd__tap_1 TAP_7419 (  );
sky130_fd_sc_hd__tap_1 TAP_742 (  );
sky130_fd_sc_hd__tap_1 TAP_7420 (  );
sky130_fd_sc_hd__tap_1 TAP_7421 (  );
sky130_fd_sc_hd__tap_1 TAP_7422 (  );
sky130_fd_sc_hd__tap_1 TAP_7423 (  );
sky130_fd_sc_hd__tap_1 TAP_7424 (  );
sky130_fd_sc_hd__tap_1 TAP_7425 (  );
sky130_fd_sc_hd__tap_1 TAP_7426 (  );
sky130_fd_sc_hd__tap_1 TAP_7427 (  );
sky130_fd_sc_hd__tap_1 TAP_7428 (  );
sky130_fd_sc_hd__tap_1 TAP_7429 (  );
sky130_fd_sc_hd__tap_1 TAP_743 (  );
sky130_fd_sc_hd__tap_1 TAP_7430 (  );
sky130_fd_sc_hd__tap_1 TAP_7431 (  );
sky130_fd_sc_hd__tap_1 TAP_7432 (  );
sky130_fd_sc_hd__tap_1 TAP_7433 (  );
sky130_fd_sc_hd__tap_1 TAP_7434 (  );
sky130_fd_sc_hd__tap_1 TAP_7435 (  );
sky130_fd_sc_hd__tap_1 TAP_7436 (  );
sky130_fd_sc_hd__tap_1 TAP_7437 (  );
sky130_fd_sc_hd__tap_1 TAP_7438 (  );
sky130_fd_sc_hd__tap_1 TAP_7439 (  );
sky130_fd_sc_hd__tap_1 TAP_744 (  );
sky130_fd_sc_hd__tap_1 TAP_7440 (  );
sky130_fd_sc_hd__tap_1 TAP_7441 (  );
sky130_fd_sc_hd__tap_1 TAP_7442 (  );
sky130_fd_sc_hd__tap_1 TAP_7443 (  );
sky130_fd_sc_hd__tap_1 TAP_7444 (  );
sky130_fd_sc_hd__tap_1 TAP_7445 (  );
sky130_fd_sc_hd__tap_1 TAP_7446 (  );
sky130_fd_sc_hd__tap_1 TAP_7447 (  );
sky130_fd_sc_hd__tap_1 TAP_7448 (  );
sky130_fd_sc_hd__tap_1 TAP_7449 (  );
sky130_fd_sc_hd__tap_1 TAP_745 (  );
sky130_fd_sc_hd__tap_1 TAP_7450 (  );
sky130_fd_sc_hd__tap_1 TAP_7451 (  );
sky130_fd_sc_hd__tap_1 TAP_7452 (  );
sky130_fd_sc_hd__tap_1 TAP_7453 (  );
sky130_fd_sc_hd__tap_1 TAP_7454 (  );
sky130_fd_sc_hd__tap_1 TAP_7455 (  );
sky130_fd_sc_hd__tap_1 TAP_7456 (  );
sky130_fd_sc_hd__tap_1 TAP_7457 (  );
sky130_fd_sc_hd__tap_1 TAP_7458 (  );
sky130_fd_sc_hd__tap_1 TAP_7459 (  );
sky130_fd_sc_hd__tap_1 TAP_746 (  );
sky130_fd_sc_hd__tap_1 TAP_7460 (  );
sky130_fd_sc_hd__tap_1 TAP_7461 (  );
sky130_fd_sc_hd__tap_1 TAP_7462 (  );
sky130_fd_sc_hd__tap_1 TAP_7463 (  );
sky130_fd_sc_hd__tap_1 TAP_7464 (  );
sky130_fd_sc_hd__tap_1 TAP_7465 (  );
sky130_fd_sc_hd__tap_1 TAP_7466 (  );
sky130_fd_sc_hd__tap_1 TAP_7467 (  );
sky130_fd_sc_hd__tap_1 TAP_7468 (  );
sky130_fd_sc_hd__tap_1 TAP_7469 (  );
sky130_fd_sc_hd__tap_1 TAP_747 (  );
sky130_fd_sc_hd__tap_1 TAP_7470 (  );
sky130_fd_sc_hd__tap_1 TAP_7471 (  );
sky130_fd_sc_hd__tap_1 TAP_7472 (  );
sky130_fd_sc_hd__tap_1 TAP_7473 (  );
sky130_fd_sc_hd__tap_1 TAP_7474 (  );
sky130_fd_sc_hd__tap_1 TAP_7475 (  );
sky130_fd_sc_hd__tap_1 TAP_7476 (  );
sky130_fd_sc_hd__tap_1 TAP_7477 (  );
sky130_fd_sc_hd__tap_1 TAP_7478 (  );
sky130_fd_sc_hd__tap_1 TAP_7479 (  );
sky130_fd_sc_hd__tap_1 TAP_748 (  );
sky130_fd_sc_hd__tap_1 TAP_7480 (  );
sky130_fd_sc_hd__tap_1 TAP_7481 (  );
sky130_fd_sc_hd__tap_1 TAP_7482 (  );
sky130_fd_sc_hd__tap_1 TAP_7483 (  );
sky130_fd_sc_hd__tap_1 TAP_7484 (  );
sky130_fd_sc_hd__tap_1 TAP_7485 (  );
sky130_fd_sc_hd__tap_1 TAP_7486 (  );
sky130_fd_sc_hd__tap_1 TAP_7487 (  );
sky130_fd_sc_hd__tap_1 TAP_7488 (  );
sky130_fd_sc_hd__tap_1 TAP_7489 (  );
sky130_fd_sc_hd__tap_1 TAP_749 (  );
sky130_fd_sc_hd__tap_1 TAP_7490 (  );
sky130_fd_sc_hd__tap_1 TAP_7491 (  );
sky130_fd_sc_hd__tap_1 TAP_7492 (  );
sky130_fd_sc_hd__tap_1 TAP_7493 (  );
sky130_fd_sc_hd__tap_1 TAP_7494 (  );
sky130_fd_sc_hd__tap_1 TAP_7495 (  );
sky130_fd_sc_hd__tap_1 TAP_7496 (  );
sky130_fd_sc_hd__tap_1 TAP_7497 (  );
sky130_fd_sc_hd__tap_1 TAP_7498 (  );
sky130_fd_sc_hd__tap_1 TAP_7499 (  );
sky130_fd_sc_hd__tap_1 TAP_750 (  );
sky130_fd_sc_hd__tap_1 TAP_7500 (  );
sky130_fd_sc_hd__tap_1 TAP_7501 (  );
sky130_fd_sc_hd__tap_1 TAP_7502 (  );
sky130_fd_sc_hd__tap_1 TAP_7503 (  );
sky130_fd_sc_hd__tap_1 TAP_7504 (  );
sky130_fd_sc_hd__tap_1 TAP_7505 (  );
sky130_fd_sc_hd__tap_1 TAP_7506 (  );
sky130_fd_sc_hd__tap_1 TAP_7507 (  );
sky130_fd_sc_hd__tap_1 TAP_7508 (  );
sky130_fd_sc_hd__tap_1 TAP_7509 (  );
sky130_fd_sc_hd__tap_1 TAP_751 (  );
sky130_fd_sc_hd__tap_1 TAP_7510 (  );
sky130_fd_sc_hd__tap_1 TAP_7511 (  );
sky130_fd_sc_hd__tap_1 TAP_7512 (  );
sky130_fd_sc_hd__tap_1 TAP_7513 (  );
sky130_fd_sc_hd__tap_1 TAP_7514 (  );
sky130_fd_sc_hd__tap_1 TAP_7515 (  );
sky130_fd_sc_hd__tap_1 TAP_7516 (  );
sky130_fd_sc_hd__tap_1 TAP_7517 (  );
sky130_fd_sc_hd__tap_1 TAP_7518 (  );
sky130_fd_sc_hd__tap_1 TAP_7519 (  );
sky130_fd_sc_hd__tap_1 TAP_752 (  );
sky130_fd_sc_hd__tap_1 TAP_7520 (  );
sky130_fd_sc_hd__tap_1 TAP_7521 (  );
sky130_fd_sc_hd__tap_1 TAP_7522 (  );
sky130_fd_sc_hd__tap_1 TAP_7523 (  );
sky130_fd_sc_hd__tap_1 TAP_7524 (  );
sky130_fd_sc_hd__tap_1 TAP_7525 (  );
sky130_fd_sc_hd__tap_1 TAP_7526 (  );
sky130_fd_sc_hd__tap_1 TAP_7527 (  );
sky130_fd_sc_hd__tap_1 TAP_7528 (  );
sky130_fd_sc_hd__tap_1 TAP_7529 (  );
sky130_fd_sc_hd__tap_1 TAP_753 (  );
sky130_fd_sc_hd__tap_1 TAP_7530 (  );
sky130_fd_sc_hd__tap_1 TAP_7531 (  );
sky130_fd_sc_hd__tap_1 TAP_7532 (  );
sky130_fd_sc_hd__tap_1 TAP_7533 (  );
sky130_fd_sc_hd__tap_1 TAP_7534 (  );
sky130_fd_sc_hd__tap_1 TAP_7535 (  );
sky130_fd_sc_hd__tap_1 TAP_7536 (  );
sky130_fd_sc_hd__tap_1 TAP_7537 (  );
sky130_fd_sc_hd__tap_1 TAP_7538 (  );
sky130_fd_sc_hd__tap_1 TAP_7539 (  );
sky130_fd_sc_hd__tap_1 TAP_754 (  );
sky130_fd_sc_hd__tap_1 TAP_7540 (  );
sky130_fd_sc_hd__tap_1 TAP_7541 (  );
sky130_fd_sc_hd__tap_1 TAP_7542 (  );
sky130_fd_sc_hd__tap_1 TAP_7543 (  );
sky130_fd_sc_hd__tap_1 TAP_7544 (  );
sky130_fd_sc_hd__tap_1 TAP_7545 (  );
sky130_fd_sc_hd__tap_1 TAP_7546 (  );
sky130_fd_sc_hd__tap_1 TAP_7547 (  );
sky130_fd_sc_hd__tap_1 TAP_7548 (  );
sky130_fd_sc_hd__tap_1 TAP_7549 (  );
sky130_fd_sc_hd__tap_1 TAP_755 (  );
sky130_fd_sc_hd__tap_1 TAP_7550 (  );
sky130_fd_sc_hd__tap_1 TAP_7551 (  );
sky130_fd_sc_hd__tap_1 TAP_7552 (  );
sky130_fd_sc_hd__tap_1 TAP_7553 (  );
sky130_fd_sc_hd__tap_1 TAP_7554 (  );
sky130_fd_sc_hd__tap_1 TAP_7555 (  );
sky130_fd_sc_hd__tap_1 TAP_7556 (  );
sky130_fd_sc_hd__tap_1 TAP_7557 (  );
sky130_fd_sc_hd__tap_1 TAP_7558 (  );
sky130_fd_sc_hd__tap_1 TAP_7559 (  );
sky130_fd_sc_hd__tap_1 TAP_756 (  );
sky130_fd_sc_hd__tap_1 TAP_7560 (  );
sky130_fd_sc_hd__tap_1 TAP_7561 (  );
sky130_fd_sc_hd__tap_1 TAP_7562 (  );
sky130_fd_sc_hd__tap_1 TAP_7563 (  );
sky130_fd_sc_hd__tap_1 TAP_7564 (  );
sky130_fd_sc_hd__tap_1 TAP_7565 (  );
sky130_fd_sc_hd__tap_1 TAP_7566 (  );
sky130_fd_sc_hd__tap_1 TAP_7567 (  );
sky130_fd_sc_hd__tap_1 TAP_7568 (  );
sky130_fd_sc_hd__tap_1 TAP_7569 (  );
sky130_fd_sc_hd__tap_1 TAP_757 (  );
sky130_fd_sc_hd__tap_1 TAP_7570 (  );
sky130_fd_sc_hd__tap_1 TAP_7571 (  );
sky130_fd_sc_hd__tap_1 TAP_7572 (  );
sky130_fd_sc_hd__tap_1 TAP_7573 (  );
sky130_fd_sc_hd__tap_1 TAP_7574 (  );
sky130_fd_sc_hd__tap_1 TAP_7575 (  );
sky130_fd_sc_hd__tap_1 TAP_7576 (  );
sky130_fd_sc_hd__tap_1 TAP_7577 (  );
sky130_fd_sc_hd__tap_1 TAP_7578 (  );
sky130_fd_sc_hd__tap_1 TAP_7579 (  );
sky130_fd_sc_hd__tap_1 TAP_758 (  );
sky130_fd_sc_hd__tap_1 TAP_7580 (  );
sky130_fd_sc_hd__tap_1 TAP_7581 (  );
sky130_fd_sc_hd__tap_1 TAP_7582 (  );
sky130_fd_sc_hd__tap_1 TAP_7583 (  );
sky130_fd_sc_hd__tap_1 TAP_7584 (  );
sky130_fd_sc_hd__tap_1 TAP_7585 (  );
sky130_fd_sc_hd__tap_1 TAP_7586 (  );
sky130_fd_sc_hd__tap_1 TAP_7587 (  );
sky130_fd_sc_hd__tap_1 TAP_7588 (  );
sky130_fd_sc_hd__tap_1 TAP_7589 (  );
sky130_fd_sc_hd__tap_1 TAP_759 (  );
sky130_fd_sc_hd__tap_1 TAP_7590 (  );
sky130_fd_sc_hd__tap_1 TAP_7591 (  );
sky130_fd_sc_hd__tap_1 TAP_7592 (  );
sky130_fd_sc_hd__tap_1 TAP_7593 (  );
sky130_fd_sc_hd__tap_1 TAP_7594 (  );
sky130_fd_sc_hd__tap_1 TAP_7595 (  );
sky130_fd_sc_hd__tap_1 TAP_7596 (  );
sky130_fd_sc_hd__tap_1 TAP_7597 (  );
sky130_fd_sc_hd__tap_1 TAP_7598 (  );
sky130_fd_sc_hd__tap_1 TAP_7599 (  );
sky130_fd_sc_hd__tap_1 TAP_760 (  );
sky130_fd_sc_hd__tap_1 TAP_7600 (  );
sky130_fd_sc_hd__tap_1 TAP_7601 (  );
sky130_fd_sc_hd__tap_1 TAP_7602 (  );
sky130_fd_sc_hd__tap_1 TAP_7603 (  );
sky130_fd_sc_hd__tap_1 TAP_7604 (  );
sky130_fd_sc_hd__tap_1 TAP_7605 (  );
sky130_fd_sc_hd__tap_1 TAP_7606 (  );
sky130_fd_sc_hd__tap_1 TAP_7607 (  );
sky130_fd_sc_hd__tap_1 TAP_7608 (  );
sky130_fd_sc_hd__tap_1 TAP_7609 (  );
sky130_fd_sc_hd__tap_1 TAP_761 (  );
sky130_fd_sc_hd__tap_1 TAP_7610 (  );
sky130_fd_sc_hd__tap_1 TAP_7611 (  );
sky130_fd_sc_hd__tap_1 TAP_7612 (  );
sky130_fd_sc_hd__tap_1 TAP_7613 (  );
sky130_fd_sc_hd__tap_1 TAP_7614 (  );
sky130_fd_sc_hd__tap_1 TAP_7615 (  );
sky130_fd_sc_hd__tap_1 TAP_7616 (  );
sky130_fd_sc_hd__tap_1 TAP_7617 (  );
sky130_fd_sc_hd__tap_1 TAP_7618 (  );
sky130_fd_sc_hd__tap_1 TAP_7619 (  );
sky130_fd_sc_hd__tap_1 TAP_762 (  );
sky130_fd_sc_hd__tap_1 TAP_7620 (  );
sky130_fd_sc_hd__tap_1 TAP_7621 (  );
sky130_fd_sc_hd__tap_1 TAP_7622 (  );
sky130_fd_sc_hd__tap_1 TAP_7623 (  );
sky130_fd_sc_hd__tap_1 TAP_7624 (  );
sky130_fd_sc_hd__tap_1 TAP_7625 (  );
sky130_fd_sc_hd__tap_1 TAP_7626 (  );
sky130_fd_sc_hd__tap_1 TAP_7627 (  );
sky130_fd_sc_hd__tap_1 TAP_7628 (  );
sky130_fd_sc_hd__tap_1 TAP_7629 (  );
sky130_fd_sc_hd__tap_1 TAP_763 (  );
sky130_fd_sc_hd__tap_1 TAP_7630 (  );
sky130_fd_sc_hd__tap_1 TAP_7631 (  );
sky130_fd_sc_hd__tap_1 TAP_7632 (  );
sky130_fd_sc_hd__tap_1 TAP_7633 (  );
sky130_fd_sc_hd__tap_1 TAP_7634 (  );
sky130_fd_sc_hd__tap_1 TAP_7635 (  );
sky130_fd_sc_hd__tap_1 TAP_7636 (  );
sky130_fd_sc_hd__tap_1 TAP_7637 (  );
sky130_fd_sc_hd__tap_1 TAP_7638 (  );
sky130_fd_sc_hd__tap_1 TAP_7639 (  );
sky130_fd_sc_hd__tap_1 TAP_764 (  );
sky130_fd_sc_hd__tap_1 TAP_7640 (  );
sky130_fd_sc_hd__tap_1 TAP_7641 (  );
sky130_fd_sc_hd__tap_1 TAP_7642 (  );
sky130_fd_sc_hd__tap_1 TAP_7643 (  );
sky130_fd_sc_hd__tap_1 TAP_7644 (  );
sky130_fd_sc_hd__tap_1 TAP_7645 (  );
sky130_fd_sc_hd__tap_1 TAP_7646 (  );
sky130_fd_sc_hd__tap_1 TAP_7647 (  );
sky130_fd_sc_hd__tap_1 TAP_7648 (  );
sky130_fd_sc_hd__tap_1 TAP_7649 (  );
sky130_fd_sc_hd__tap_1 TAP_765 (  );
sky130_fd_sc_hd__tap_1 TAP_7650 (  );
sky130_fd_sc_hd__tap_1 TAP_7651 (  );
sky130_fd_sc_hd__tap_1 TAP_7652 (  );
sky130_fd_sc_hd__tap_1 TAP_7653 (  );
sky130_fd_sc_hd__tap_1 TAP_7654 (  );
sky130_fd_sc_hd__tap_1 TAP_7655 (  );
sky130_fd_sc_hd__tap_1 TAP_7656 (  );
sky130_fd_sc_hd__tap_1 TAP_7657 (  );
sky130_fd_sc_hd__tap_1 TAP_7658 (  );
sky130_fd_sc_hd__tap_1 TAP_7659 (  );
sky130_fd_sc_hd__tap_1 TAP_766 (  );
sky130_fd_sc_hd__tap_1 TAP_7660 (  );
sky130_fd_sc_hd__tap_1 TAP_7661 (  );
sky130_fd_sc_hd__tap_1 TAP_7662 (  );
sky130_fd_sc_hd__tap_1 TAP_7663 (  );
sky130_fd_sc_hd__tap_1 TAP_7664 (  );
sky130_fd_sc_hd__tap_1 TAP_7665 (  );
sky130_fd_sc_hd__tap_1 TAP_7666 (  );
sky130_fd_sc_hd__tap_1 TAP_7667 (  );
sky130_fd_sc_hd__tap_1 TAP_7668 (  );
sky130_fd_sc_hd__tap_1 TAP_7669 (  );
sky130_fd_sc_hd__tap_1 TAP_767 (  );
sky130_fd_sc_hd__tap_1 TAP_7670 (  );
sky130_fd_sc_hd__tap_1 TAP_7671 (  );
sky130_fd_sc_hd__tap_1 TAP_7672 (  );
sky130_fd_sc_hd__tap_1 TAP_7673 (  );
sky130_fd_sc_hd__tap_1 TAP_7674 (  );
sky130_fd_sc_hd__tap_1 TAP_7675 (  );
sky130_fd_sc_hd__tap_1 TAP_7676 (  );
sky130_fd_sc_hd__tap_1 TAP_7677 (  );
sky130_fd_sc_hd__tap_1 TAP_7678 (  );
sky130_fd_sc_hd__tap_1 TAP_7679 (  );
sky130_fd_sc_hd__tap_1 TAP_768 (  );
sky130_fd_sc_hd__tap_1 TAP_7680 (  );
sky130_fd_sc_hd__tap_1 TAP_7681 (  );
sky130_fd_sc_hd__tap_1 TAP_7682 (  );
sky130_fd_sc_hd__tap_1 TAP_7683 (  );
sky130_fd_sc_hd__tap_1 TAP_7684 (  );
sky130_fd_sc_hd__tap_1 TAP_7685 (  );
sky130_fd_sc_hd__tap_1 TAP_7686 (  );
sky130_fd_sc_hd__tap_1 TAP_7687 (  );
sky130_fd_sc_hd__tap_1 TAP_7688 (  );
sky130_fd_sc_hd__tap_1 TAP_7689 (  );
sky130_fd_sc_hd__tap_1 TAP_769 (  );
sky130_fd_sc_hd__tap_1 TAP_7690 (  );
sky130_fd_sc_hd__tap_1 TAP_7691 (  );
sky130_fd_sc_hd__tap_1 TAP_7692 (  );
sky130_fd_sc_hd__tap_1 TAP_7693 (  );
sky130_fd_sc_hd__tap_1 TAP_7694 (  );
sky130_fd_sc_hd__tap_1 TAP_7695 (  );
sky130_fd_sc_hd__tap_1 TAP_7696 (  );
sky130_fd_sc_hd__tap_1 TAP_7697 (  );
sky130_fd_sc_hd__tap_1 TAP_7698 (  );
sky130_fd_sc_hd__tap_1 TAP_7699 (  );
sky130_fd_sc_hd__tap_1 TAP_770 (  );
sky130_fd_sc_hd__tap_1 TAP_7700 (  );
sky130_fd_sc_hd__tap_1 TAP_7701 (  );
sky130_fd_sc_hd__tap_1 TAP_7702 (  );
sky130_fd_sc_hd__tap_1 TAP_7703 (  );
sky130_fd_sc_hd__tap_1 TAP_7704 (  );
sky130_fd_sc_hd__tap_1 TAP_7705 (  );
sky130_fd_sc_hd__tap_1 TAP_7706 (  );
sky130_fd_sc_hd__tap_1 TAP_7707 (  );
sky130_fd_sc_hd__tap_1 TAP_7708 (  );
sky130_fd_sc_hd__tap_1 TAP_7709 (  );
sky130_fd_sc_hd__tap_1 TAP_771 (  );
sky130_fd_sc_hd__tap_1 TAP_7710 (  );
sky130_fd_sc_hd__tap_1 TAP_7711 (  );
sky130_fd_sc_hd__tap_1 TAP_7712 (  );
sky130_fd_sc_hd__tap_1 TAP_7713 (  );
sky130_fd_sc_hd__tap_1 TAP_7714 (  );
sky130_fd_sc_hd__tap_1 TAP_7715 (  );
sky130_fd_sc_hd__tap_1 TAP_7716 (  );
sky130_fd_sc_hd__tap_1 TAP_7717 (  );
sky130_fd_sc_hd__tap_1 TAP_7718 (  );
sky130_fd_sc_hd__tap_1 TAP_7719 (  );
sky130_fd_sc_hd__tap_1 TAP_772 (  );
sky130_fd_sc_hd__tap_1 TAP_7720 (  );
sky130_fd_sc_hd__tap_1 TAP_7721 (  );
sky130_fd_sc_hd__tap_1 TAP_7722 (  );
sky130_fd_sc_hd__tap_1 TAP_7723 (  );
sky130_fd_sc_hd__tap_1 TAP_7724 (  );
sky130_fd_sc_hd__tap_1 TAP_7725 (  );
sky130_fd_sc_hd__tap_1 TAP_7726 (  );
sky130_fd_sc_hd__tap_1 TAP_7727 (  );
sky130_fd_sc_hd__tap_1 TAP_7728 (  );
sky130_fd_sc_hd__tap_1 TAP_7729 (  );
sky130_fd_sc_hd__tap_1 TAP_773 (  );
sky130_fd_sc_hd__tap_1 TAP_7730 (  );
sky130_fd_sc_hd__tap_1 TAP_7731 (  );
sky130_fd_sc_hd__tap_1 TAP_7732 (  );
sky130_fd_sc_hd__tap_1 TAP_7733 (  );
sky130_fd_sc_hd__tap_1 TAP_7734 (  );
sky130_fd_sc_hd__tap_1 TAP_7735 (  );
sky130_fd_sc_hd__tap_1 TAP_7736 (  );
sky130_fd_sc_hd__tap_1 TAP_7737 (  );
sky130_fd_sc_hd__tap_1 TAP_7738 (  );
sky130_fd_sc_hd__tap_1 TAP_7739 (  );
sky130_fd_sc_hd__tap_1 TAP_774 (  );
sky130_fd_sc_hd__tap_1 TAP_7740 (  );
sky130_fd_sc_hd__tap_1 TAP_7741 (  );
sky130_fd_sc_hd__tap_1 TAP_7742 (  );
sky130_fd_sc_hd__tap_1 TAP_7743 (  );
sky130_fd_sc_hd__tap_1 TAP_7744 (  );
sky130_fd_sc_hd__tap_1 TAP_7745 (  );
sky130_fd_sc_hd__tap_1 TAP_7746 (  );
sky130_fd_sc_hd__tap_1 TAP_7747 (  );
sky130_fd_sc_hd__tap_1 TAP_7748 (  );
sky130_fd_sc_hd__tap_1 TAP_7749 (  );
sky130_fd_sc_hd__tap_1 TAP_775 (  );
sky130_fd_sc_hd__tap_1 TAP_7750 (  );
sky130_fd_sc_hd__tap_1 TAP_7751 (  );
sky130_fd_sc_hd__tap_1 TAP_7752 (  );
sky130_fd_sc_hd__tap_1 TAP_7753 (  );
sky130_fd_sc_hd__tap_1 TAP_7754 (  );
sky130_fd_sc_hd__tap_1 TAP_7755 (  );
sky130_fd_sc_hd__tap_1 TAP_7756 (  );
sky130_fd_sc_hd__tap_1 TAP_7757 (  );
sky130_fd_sc_hd__tap_1 TAP_7758 (  );
sky130_fd_sc_hd__tap_1 TAP_7759 (  );
sky130_fd_sc_hd__tap_1 TAP_776 (  );
sky130_fd_sc_hd__tap_1 TAP_7760 (  );
sky130_fd_sc_hd__tap_1 TAP_7761 (  );
sky130_fd_sc_hd__tap_1 TAP_7762 (  );
sky130_fd_sc_hd__tap_1 TAP_7763 (  );
sky130_fd_sc_hd__tap_1 TAP_7764 (  );
sky130_fd_sc_hd__tap_1 TAP_7765 (  );
sky130_fd_sc_hd__tap_1 TAP_7766 (  );
sky130_fd_sc_hd__tap_1 TAP_7767 (  );
sky130_fd_sc_hd__tap_1 TAP_7768 (  );
sky130_fd_sc_hd__tap_1 TAP_7769 (  );
sky130_fd_sc_hd__tap_1 TAP_777 (  );
sky130_fd_sc_hd__tap_1 TAP_7770 (  );
sky130_fd_sc_hd__tap_1 TAP_7771 (  );
sky130_fd_sc_hd__tap_1 TAP_7772 (  );
sky130_fd_sc_hd__tap_1 TAP_7773 (  );
sky130_fd_sc_hd__tap_1 TAP_7774 (  );
sky130_fd_sc_hd__tap_1 TAP_7775 (  );
sky130_fd_sc_hd__tap_1 TAP_7776 (  );
sky130_fd_sc_hd__tap_1 TAP_7777 (  );
sky130_fd_sc_hd__tap_1 TAP_7778 (  );
sky130_fd_sc_hd__tap_1 TAP_7779 (  );
sky130_fd_sc_hd__tap_1 TAP_778 (  );
sky130_fd_sc_hd__tap_1 TAP_7780 (  );
sky130_fd_sc_hd__tap_1 TAP_7781 (  );
sky130_fd_sc_hd__tap_1 TAP_7782 (  );
sky130_fd_sc_hd__tap_1 TAP_7783 (  );
sky130_fd_sc_hd__tap_1 TAP_7784 (  );
sky130_fd_sc_hd__tap_1 TAP_7785 (  );
sky130_fd_sc_hd__tap_1 TAP_7786 (  );
sky130_fd_sc_hd__tap_1 TAP_7787 (  );
sky130_fd_sc_hd__tap_1 TAP_7788 (  );
sky130_fd_sc_hd__tap_1 TAP_7789 (  );
sky130_fd_sc_hd__tap_1 TAP_779 (  );
sky130_fd_sc_hd__tap_1 TAP_7790 (  );
sky130_fd_sc_hd__tap_1 TAP_7791 (  );
sky130_fd_sc_hd__tap_1 TAP_7792 (  );
sky130_fd_sc_hd__tap_1 TAP_7793 (  );
sky130_fd_sc_hd__tap_1 TAP_7794 (  );
sky130_fd_sc_hd__tap_1 TAP_7795 (  );
sky130_fd_sc_hd__tap_1 TAP_7796 (  );
sky130_fd_sc_hd__tap_1 TAP_7797 (  );
sky130_fd_sc_hd__tap_1 TAP_7798 (  );
sky130_fd_sc_hd__tap_1 TAP_7799 (  );
sky130_fd_sc_hd__tap_1 TAP_780 (  );
sky130_fd_sc_hd__tap_1 TAP_7800 (  );
sky130_fd_sc_hd__tap_1 TAP_7801 (  );
sky130_fd_sc_hd__tap_1 TAP_7802 (  );
sky130_fd_sc_hd__tap_1 TAP_7803 (  );
sky130_fd_sc_hd__tap_1 TAP_7804 (  );
sky130_fd_sc_hd__tap_1 TAP_7805 (  );
sky130_fd_sc_hd__tap_1 TAP_7806 (  );
sky130_fd_sc_hd__tap_1 TAP_7807 (  );
sky130_fd_sc_hd__tap_1 TAP_7808 (  );
sky130_fd_sc_hd__tap_1 TAP_7809 (  );
sky130_fd_sc_hd__tap_1 TAP_781 (  );
sky130_fd_sc_hd__tap_1 TAP_7810 (  );
sky130_fd_sc_hd__tap_1 TAP_7811 (  );
sky130_fd_sc_hd__tap_1 TAP_7812 (  );
sky130_fd_sc_hd__tap_1 TAP_7813 (  );
sky130_fd_sc_hd__tap_1 TAP_7814 (  );
sky130_fd_sc_hd__tap_1 TAP_7815 (  );
sky130_fd_sc_hd__tap_1 TAP_7816 (  );
sky130_fd_sc_hd__tap_1 TAP_7817 (  );
sky130_fd_sc_hd__tap_1 TAP_7818 (  );
sky130_fd_sc_hd__tap_1 TAP_7819 (  );
sky130_fd_sc_hd__tap_1 TAP_782 (  );
sky130_fd_sc_hd__tap_1 TAP_7820 (  );
sky130_fd_sc_hd__tap_1 TAP_7821 (  );
sky130_fd_sc_hd__tap_1 TAP_7822 (  );
sky130_fd_sc_hd__tap_1 TAP_7823 (  );
sky130_fd_sc_hd__tap_1 TAP_7824 (  );
sky130_fd_sc_hd__tap_1 TAP_7825 (  );
sky130_fd_sc_hd__tap_1 TAP_7826 (  );
sky130_fd_sc_hd__tap_1 TAP_7827 (  );
sky130_fd_sc_hd__tap_1 TAP_7828 (  );
sky130_fd_sc_hd__tap_1 TAP_7829 (  );
sky130_fd_sc_hd__tap_1 TAP_783 (  );
sky130_fd_sc_hd__tap_1 TAP_7830 (  );
sky130_fd_sc_hd__tap_1 TAP_7831 (  );
sky130_fd_sc_hd__tap_1 TAP_7832 (  );
sky130_fd_sc_hd__tap_1 TAP_7833 (  );
sky130_fd_sc_hd__tap_1 TAP_7834 (  );
sky130_fd_sc_hd__tap_1 TAP_7835 (  );
sky130_fd_sc_hd__tap_1 TAP_7836 (  );
sky130_fd_sc_hd__tap_1 TAP_7837 (  );
sky130_fd_sc_hd__tap_1 TAP_7838 (  );
sky130_fd_sc_hd__tap_1 TAP_7839 (  );
sky130_fd_sc_hd__tap_1 TAP_784 (  );
sky130_fd_sc_hd__tap_1 TAP_7840 (  );
sky130_fd_sc_hd__tap_1 TAP_7841 (  );
sky130_fd_sc_hd__tap_1 TAP_7842 (  );
sky130_fd_sc_hd__tap_1 TAP_7843 (  );
sky130_fd_sc_hd__tap_1 TAP_7844 (  );
sky130_fd_sc_hd__tap_1 TAP_7845 (  );
sky130_fd_sc_hd__tap_1 TAP_7846 (  );
sky130_fd_sc_hd__tap_1 TAP_7847 (  );
sky130_fd_sc_hd__tap_1 TAP_7848 (  );
sky130_fd_sc_hd__tap_1 TAP_7849 (  );
sky130_fd_sc_hd__tap_1 TAP_785 (  );
sky130_fd_sc_hd__tap_1 TAP_7850 (  );
sky130_fd_sc_hd__tap_1 TAP_7851 (  );
sky130_fd_sc_hd__tap_1 TAP_7852 (  );
sky130_fd_sc_hd__tap_1 TAP_7853 (  );
sky130_fd_sc_hd__tap_1 TAP_7854 (  );
sky130_fd_sc_hd__tap_1 TAP_7855 (  );
sky130_fd_sc_hd__tap_1 TAP_7856 (  );
sky130_fd_sc_hd__tap_1 TAP_7857 (  );
sky130_fd_sc_hd__tap_1 TAP_7858 (  );
sky130_fd_sc_hd__tap_1 TAP_7859 (  );
sky130_fd_sc_hd__tap_1 TAP_786 (  );
sky130_fd_sc_hd__tap_1 TAP_7860 (  );
sky130_fd_sc_hd__tap_1 TAP_7861 (  );
sky130_fd_sc_hd__tap_1 TAP_7862 (  );
sky130_fd_sc_hd__tap_1 TAP_7863 (  );
sky130_fd_sc_hd__tap_1 TAP_7864 (  );
sky130_fd_sc_hd__tap_1 TAP_7865 (  );
sky130_fd_sc_hd__tap_1 TAP_7866 (  );
sky130_fd_sc_hd__tap_1 TAP_7867 (  );
sky130_fd_sc_hd__tap_1 TAP_7868 (  );
sky130_fd_sc_hd__tap_1 TAP_7869 (  );
sky130_fd_sc_hd__tap_1 TAP_787 (  );
sky130_fd_sc_hd__tap_1 TAP_7870 (  );
sky130_fd_sc_hd__tap_1 TAP_7871 (  );
sky130_fd_sc_hd__tap_1 TAP_7872 (  );
sky130_fd_sc_hd__tap_1 TAP_7873 (  );
sky130_fd_sc_hd__tap_1 TAP_7874 (  );
sky130_fd_sc_hd__tap_1 TAP_7875 (  );
sky130_fd_sc_hd__tap_1 TAP_7876 (  );
sky130_fd_sc_hd__tap_1 TAP_7877 (  );
sky130_fd_sc_hd__tap_1 TAP_7878 (  );
sky130_fd_sc_hd__tap_1 TAP_7879 (  );
sky130_fd_sc_hd__tap_1 TAP_788 (  );
sky130_fd_sc_hd__tap_1 TAP_7880 (  );
sky130_fd_sc_hd__tap_1 TAP_7881 (  );
sky130_fd_sc_hd__tap_1 TAP_7882 (  );
sky130_fd_sc_hd__tap_1 TAP_7883 (  );
sky130_fd_sc_hd__tap_1 TAP_7884 (  );
sky130_fd_sc_hd__tap_1 TAP_7885 (  );
sky130_fd_sc_hd__tap_1 TAP_7886 (  );
sky130_fd_sc_hd__tap_1 TAP_7887 (  );
sky130_fd_sc_hd__tap_1 TAP_7888 (  );
sky130_fd_sc_hd__tap_1 TAP_7889 (  );
sky130_fd_sc_hd__tap_1 TAP_789 (  );
sky130_fd_sc_hd__tap_1 TAP_7890 (  );
sky130_fd_sc_hd__tap_1 TAP_7891 (  );
sky130_fd_sc_hd__tap_1 TAP_7892 (  );
sky130_fd_sc_hd__tap_1 TAP_7893 (  );
sky130_fd_sc_hd__tap_1 TAP_7894 (  );
sky130_fd_sc_hd__tap_1 TAP_7895 (  );
sky130_fd_sc_hd__tap_1 TAP_7896 (  );
sky130_fd_sc_hd__tap_1 TAP_7897 (  );
sky130_fd_sc_hd__tap_1 TAP_7898 (  );
sky130_fd_sc_hd__tap_1 TAP_7899 (  );
sky130_fd_sc_hd__tap_1 TAP_790 (  );
sky130_fd_sc_hd__tap_1 TAP_7900 (  );
sky130_fd_sc_hd__tap_1 TAP_7901 (  );
sky130_fd_sc_hd__tap_1 TAP_7902 (  );
sky130_fd_sc_hd__tap_1 TAP_7903 (  );
sky130_fd_sc_hd__tap_1 TAP_7904 (  );
sky130_fd_sc_hd__tap_1 TAP_7905 (  );
sky130_fd_sc_hd__tap_1 TAP_7906 (  );
sky130_fd_sc_hd__tap_1 TAP_7907 (  );
sky130_fd_sc_hd__tap_1 TAP_7908 (  );
sky130_fd_sc_hd__tap_1 TAP_7909 (  );
sky130_fd_sc_hd__tap_1 TAP_791 (  );
sky130_fd_sc_hd__tap_1 TAP_7910 (  );
sky130_fd_sc_hd__tap_1 TAP_7911 (  );
sky130_fd_sc_hd__tap_1 TAP_7912 (  );
sky130_fd_sc_hd__tap_1 TAP_7913 (  );
sky130_fd_sc_hd__tap_1 TAP_7914 (  );
sky130_fd_sc_hd__tap_1 TAP_7915 (  );
sky130_fd_sc_hd__tap_1 TAP_7916 (  );
sky130_fd_sc_hd__tap_1 TAP_7917 (  );
sky130_fd_sc_hd__tap_1 TAP_7918 (  );
sky130_fd_sc_hd__tap_1 TAP_7919 (  );
sky130_fd_sc_hd__tap_1 TAP_792 (  );
sky130_fd_sc_hd__tap_1 TAP_7920 (  );
sky130_fd_sc_hd__tap_1 TAP_7921 (  );
sky130_fd_sc_hd__tap_1 TAP_7922 (  );
sky130_fd_sc_hd__tap_1 TAP_7923 (  );
sky130_fd_sc_hd__tap_1 TAP_7924 (  );
sky130_fd_sc_hd__tap_1 TAP_7925 (  );
sky130_fd_sc_hd__tap_1 TAP_7926 (  );
sky130_fd_sc_hd__tap_1 TAP_7927 (  );
sky130_fd_sc_hd__tap_1 TAP_7928 (  );
sky130_fd_sc_hd__tap_1 TAP_7929 (  );
sky130_fd_sc_hd__tap_1 TAP_793 (  );
sky130_fd_sc_hd__tap_1 TAP_7930 (  );
sky130_fd_sc_hd__tap_1 TAP_7931 (  );
sky130_fd_sc_hd__tap_1 TAP_7932 (  );
sky130_fd_sc_hd__tap_1 TAP_7933 (  );
sky130_fd_sc_hd__tap_1 TAP_7934 (  );
sky130_fd_sc_hd__tap_1 TAP_7935 (  );
sky130_fd_sc_hd__tap_1 TAP_7936 (  );
sky130_fd_sc_hd__tap_1 TAP_7937 (  );
sky130_fd_sc_hd__tap_1 TAP_7938 (  );
sky130_fd_sc_hd__tap_1 TAP_7939 (  );
sky130_fd_sc_hd__tap_1 TAP_794 (  );
sky130_fd_sc_hd__tap_1 TAP_7940 (  );
sky130_fd_sc_hd__tap_1 TAP_7941 (  );
sky130_fd_sc_hd__tap_1 TAP_7942 (  );
sky130_fd_sc_hd__tap_1 TAP_7943 (  );
sky130_fd_sc_hd__tap_1 TAP_7944 (  );
sky130_fd_sc_hd__tap_1 TAP_7945 (  );
sky130_fd_sc_hd__tap_1 TAP_7946 (  );
sky130_fd_sc_hd__tap_1 TAP_7947 (  );
sky130_fd_sc_hd__tap_1 TAP_7948 (  );
sky130_fd_sc_hd__tap_1 TAP_7949 (  );
sky130_fd_sc_hd__tap_1 TAP_795 (  );
sky130_fd_sc_hd__tap_1 TAP_7950 (  );
sky130_fd_sc_hd__tap_1 TAP_7951 (  );
sky130_fd_sc_hd__tap_1 TAP_7952 (  );
sky130_fd_sc_hd__tap_1 TAP_7953 (  );
sky130_fd_sc_hd__tap_1 TAP_7954 (  );
sky130_fd_sc_hd__tap_1 TAP_7955 (  );
sky130_fd_sc_hd__tap_1 TAP_7956 (  );
sky130_fd_sc_hd__tap_1 TAP_7957 (  );
sky130_fd_sc_hd__tap_1 TAP_7958 (  );
sky130_fd_sc_hd__tap_1 TAP_7959 (  );
sky130_fd_sc_hd__tap_1 TAP_796 (  );
sky130_fd_sc_hd__tap_1 TAP_7960 (  );
sky130_fd_sc_hd__tap_1 TAP_7961 (  );
sky130_fd_sc_hd__tap_1 TAP_7962 (  );
sky130_fd_sc_hd__tap_1 TAP_7963 (  );
sky130_fd_sc_hd__tap_1 TAP_7964 (  );
sky130_fd_sc_hd__tap_1 TAP_7965 (  );
sky130_fd_sc_hd__tap_1 TAP_7966 (  );
sky130_fd_sc_hd__tap_1 TAP_7967 (  );
sky130_fd_sc_hd__tap_1 TAP_7968 (  );
sky130_fd_sc_hd__tap_1 TAP_7969 (  );
sky130_fd_sc_hd__tap_1 TAP_797 (  );
sky130_fd_sc_hd__tap_1 TAP_7970 (  );
sky130_fd_sc_hd__tap_1 TAP_7971 (  );
sky130_fd_sc_hd__tap_1 TAP_7972 (  );
sky130_fd_sc_hd__tap_1 TAP_7973 (  );
sky130_fd_sc_hd__tap_1 TAP_7974 (  );
sky130_fd_sc_hd__tap_1 TAP_7975 (  );
sky130_fd_sc_hd__tap_1 TAP_7976 (  );
sky130_fd_sc_hd__tap_1 TAP_7977 (  );
sky130_fd_sc_hd__tap_1 TAP_7978 (  );
sky130_fd_sc_hd__tap_1 TAP_7979 (  );
sky130_fd_sc_hd__tap_1 TAP_798 (  );
sky130_fd_sc_hd__tap_1 TAP_7980 (  );
sky130_fd_sc_hd__tap_1 TAP_7981 (  );
sky130_fd_sc_hd__tap_1 TAP_7982 (  );
sky130_fd_sc_hd__tap_1 TAP_7983 (  );
sky130_fd_sc_hd__tap_1 TAP_7984 (  );
sky130_fd_sc_hd__tap_1 TAP_7985 (  );
sky130_fd_sc_hd__tap_1 TAP_7986 (  );
sky130_fd_sc_hd__tap_1 TAP_7987 (  );
sky130_fd_sc_hd__tap_1 TAP_7988 (  );
sky130_fd_sc_hd__tap_1 TAP_7989 (  );
sky130_fd_sc_hd__tap_1 TAP_799 (  );
sky130_fd_sc_hd__tap_1 TAP_7990 (  );
sky130_fd_sc_hd__tap_1 TAP_7991 (  );
sky130_fd_sc_hd__tap_1 TAP_7992 (  );
sky130_fd_sc_hd__tap_1 TAP_7993 (  );
sky130_fd_sc_hd__tap_1 TAP_7994 (  );
sky130_fd_sc_hd__tap_1 TAP_7995 (  );
sky130_fd_sc_hd__tap_1 TAP_7996 (  );
sky130_fd_sc_hd__tap_1 TAP_7997 (  );
sky130_fd_sc_hd__tap_1 TAP_7998 (  );
sky130_fd_sc_hd__tap_1 TAP_7999 (  );
sky130_fd_sc_hd__tap_1 TAP_800 (  );
sky130_fd_sc_hd__tap_1 TAP_8000 (  );
sky130_fd_sc_hd__tap_1 TAP_8001 (  );
sky130_fd_sc_hd__tap_1 TAP_8002 (  );
sky130_fd_sc_hd__tap_1 TAP_8003 (  );
sky130_fd_sc_hd__tap_1 TAP_8004 (  );
sky130_fd_sc_hd__tap_1 TAP_8005 (  );
sky130_fd_sc_hd__tap_1 TAP_8006 (  );
sky130_fd_sc_hd__tap_1 TAP_8007 (  );
sky130_fd_sc_hd__tap_1 TAP_8008 (  );
sky130_fd_sc_hd__tap_1 TAP_8009 (  );
sky130_fd_sc_hd__tap_1 TAP_801 (  );
sky130_fd_sc_hd__tap_1 TAP_8010 (  );
sky130_fd_sc_hd__tap_1 TAP_8011 (  );
sky130_fd_sc_hd__tap_1 TAP_8012 (  );
sky130_fd_sc_hd__tap_1 TAP_8013 (  );
sky130_fd_sc_hd__tap_1 TAP_8014 (  );
sky130_fd_sc_hd__tap_1 TAP_8015 (  );
sky130_fd_sc_hd__tap_1 TAP_8016 (  );
sky130_fd_sc_hd__tap_1 TAP_8017 (  );
sky130_fd_sc_hd__tap_1 TAP_8018 (  );
sky130_fd_sc_hd__tap_1 TAP_8019 (  );
sky130_fd_sc_hd__tap_1 TAP_802 (  );
sky130_fd_sc_hd__tap_1 TAP_8020 (  );
sky130_fd_sc_hd__tap_1 TAP_8021 (  );
sky130_fd_sc_hd__tap_1 TAP_8022 (  );
sky130_fd_sc_hd__tap_1 TAP_8023 (  );
sky130_fd_sc_hd__tap_1 TAP_8024 (  );
sky130_fd_sc_hd__tap_1 TAP_8025 (  );
sky130_fd_sc_hd__tap_1 TAP_8026 (  );
sky130_fd_sc_hd__tap_1 TAP_8027 (  );
sky130_fd_sc_hd__tap_1 TAP_8028 (  );
sky130_fd_sc_hd__tap_1 TAP_8029 (  );
sky130_fd_sc_hd__tap_1 TAP_803 (  );
sky130_fd_sc_hd__tap_1 TAP_8030 (  );
sky130_fd_sc_hd__tap_1 TAP_8031 (  );
sky130_fd_sc_hd__tap_1 TAP_8032 (  );
sky130_fd_sc_hd__tap_1 TAP_8033 (  );
sky130_fd_sc_hd__tap_1 TAP_8034 (  );
sky130_fd_sc_hd__tap_1 TAP_8035 (  );
sky130_fd_sc_hd__tap_1 TAP_8036 (  );
sky130_fd_sc_hd__tap_1 TAP_8037 (  );
sky130_fd_sc_hd__tap_1 TAP_8038 (  );
sky130_fd_sc_hd__tap_1 TAP_8039 (  );
sky130_fd_sc_hd__tap_1 TAP_804 (  );
sky130_fd_sc_hd__tap_1 TAP_8040 (  );
sky130_fd_sc_hd__tap_1 TAP_8041 (  );
sky130_fd_sc_hd__tap_1 TAP_8042 (  );
sky130_fd_sc_hd__tap_1 TAP_8043 (  );
sky130_fd_sc_hd__tap_1 TAP_8044 (  );
sky130_fd_sc_hd__tap_1 TAP_8045 (  );
sky130_fd_sc_hd__tap_1 TAP_8046 (  );
sky130_fd_sc_hd__tap_1 TAP_8047 (  );
sky130_fd_sc_hd__tap_1 TAP_8048 (  );
sky130_fd_sc_hd__tap_1 TAP_8049 (  );
sky130_fd_sc_hd__tap_1 TAP_805 (  );
sky130_fd_sc_hd__tap_1 TAP_8050 (  );
sky130_fd_sc_hd__tap_1 TAP_8051 (  );
sky130_fd_sc_hd__tap_1 TAP_8052 (  );
sky130_fd_sc_hd__tap_1 TAP_8053 (  );
sky130_fd_sc_hd__tap_1 TAP_8054 (  );
sky130_fd_sc_hd__tap_1 TAP_8055 (  );
sky130_fd_sc_hd__tap_1 TAP_8056 (  );
sky130_fd_sc_hd__tap_1 TAP_8057 (  );
sky130_fd_sc_hd__tap_1 TAP_8058 (  );
sky130_fd_sc_hd__tap_1 TAP_8059 (  );
sky130_fd_sc_hd__tap_1 TAP_806 (  );
sky130_fd_sc_hd__tap_1 TAP_8060 (  );
sky130_fd_sc_hd__tap_1 TAP_8061 (  );
sky130_fd_sc_hd__tap_1 TAP_8062 (  );
sky130_fd_sc_hd__tap_1 TAP_8063 (  );
sky130_fd_sc_hd__tap_1 TAP_8064 (  );
sky130_fd_sc_hd__tap_1 TAP_8065 (  );
sky130_fd_sc_hd__tap_1 TAP_8066 (  );
sky130_fd_sc_hd__tap_1 TAP_8067 (  );
sky130_fd_sc_hd__tap_1 TAP_8068 (  );
sky130_fd_sc_hd__tap_1 TAP_8069 (  );
sky130_fd_sc_hd__tap_1 TAP_807 (  );
sky130_fd_sc_hd__tap_1 TAP_8070 (  );
sky130_fd_sc_hd__tap_1 TAP_8071 (  );
sky130_fd_sc_hd__tap_1 TAP_8072 (  );
sky130_fd_sc_hd__tap_1 TAP_8073 (  );
sky130_fd_sc_hd__tap_1 TAP_8074 (  );
sky130_fd_sc_hd__tap_1 TAP_8075 (  );
sky130_fd_sc_hd__tap_1 TAP_8076 (  );
sky130_fd_sc_hd__tap_1 TAP_8077 (  );
sky130_fd_sc_hd__tap_1 TAP_8078 (  );
sky130_fd_sc_hd__tap_1 TAP_8079 (  );
sky130_fd_sc_hd__tap_1 TAP_808 (  );
sky130_fd_sc_hd__tap_1 TAP_8080 (  );
sky130_fd_sc_hd__tap_1 TAP_8081 (  );
sky130_fd_sc_hd__tap_1 TAP_8082 (  );
sky130_fd_sc_hd__tap_1 TAP_8083 (  );
sky130_fd_sc_hd__tap_1 TAP_8084 (  );
sky130_fd_sc_hd__tap_1 TAP_8085 (  );
sky130_fd_sc_hd__tap_1 TAP_8086 (  );
sky130_fd_sc_hd__tap_1 TAP_8087 (  );
sky130_fd_sc_hd__tap_1 TAP_8088 (  );
sky130_fd_sc_hd__tap_1 TAP_8089 (  );
sky130_fd_sc_hd__tap_1 TAP_809 (  );
sky130_fd_sc_hd__tap_1 TAP_8090 (  );
sky130_fd_sc_hd__tap_1 TAP_8091 (  );
sky130_fd_sc_hd__tap_1 TAP_8092 (  );
sky130_fd_sc_hd__tap_1 TAP_8093 (  );
sky130_fd_sc_hd__tap_1 TAP_8094 (  );
sky130_fd_sc_hd__tap_1 TAP_8095 (  );
sky130_fd_sc_hd__tap_1 TAP_8096 (  );
sky130_fd_sc_hd__tap_1 TAP_8097 (  );
sky130_fd_sc_hd__tap_1 TAP_8098 (  );
sky130_fd_sc_hd__tap_1 TAP_8099 (  );
sky130_fd_sc_hd__tap_1 TAP_810 (  );
sky130_fd_sc_hd__tap_1 TAP_8100 (  );
sky130_fd_sc_hd__tap_1 TAP_8101 (  );
sky130_fd_sc_hd__tap_1 TAP_8102 (  );
sky130_fd_sc_hd__tap_1 TAP_8103 (  );
sky130_fd_sc_hd__tap_1 TAP_8104 (  );
sky130_fd_sc_hd__tap_1 TAP_8105 (  );
sky130_fd_sc_hd__tap_1 TAP_8106 (  );
sky130_fd_sc_hd__tap_1 TAP_8107 (  );
sky130_fd_sc_hd__tap_1 TAP_8108 (  );
sky130_fd_sc_hd__tap_1 TAP_8109 (  );
sky130_fd_sc_hd__tap_1 TAP_811 (  );
sky130_fd_sc_hd__tap_1 TAP_8110 (  );
sky130_fd_sc_hd__tap_1 TAP_8111 (  );
sky130_fd_sc_hd__tap_1 TAP_8112 (  );
sky130_fd_sc_hd__tap_1 TAP_8113 (  );
sky130_fd_sc_hd__tap_1 TAP_8114 (  );
sky130_fd_sc_hd__tap_1 TAP_8115 (  );
sky130_fd_sc_hd__tap_1 TAP_8116 (  );
sky130_fd_sc_hd__tap_1 TAP_8117 (  );
sky130_fd_sc_hd__tap_1 TAP_8118 (  );
sky130_fd_sc_hd__tap_1 TAP_8119 (  );
sky130_fd_sc_hd__tap_1 TAP_812 (  );
sky130_fd_sc_hd__tap_1 TAP_8120 (  );
sky130_fd_sc_hd__tap_1 TAP_8121 (  );
sky130_fd_sc_hd__tap_1 TAP_8122 (  );
sky130_fd_sc_hd__tap_1 TAP_8123 (  );
sky130_fd_sc_hd__tap_1 TAP_8124 (  );
sky130_fd_sc_hd__tap_1 TAP_8125 (  );
sky130_fd_sc_hd__tap_1 TAP_8126 (  );
sky130_fd_sc_hd__tap_1 TAP_8127 (  );
sky130_fd_sc_hd__tap_1 TAP_8128 (  );
sky130_fd_sc_hd__tap_1 TAP_8129 (  );
sky130_fd_sc_hd__tap_1 TAP_813 (  );
sky130_fd_sc_hd__tap_1 TAP_8130 (  );
sky130_fd_sc_hd__tap_1 TAP_8131 (  );
sky130_fd_sc_hd__tap_1 TAP_8132 (  );
sky130_fd_sc_hd__tap_1 TAP_8133 (  );
sky130_fd_sc_hd__tap_1 TAP_8134 (  );
sky130_fd_sc_hd__tap_1 TAP_8135 (  );
sky130_fd_sc_hd__tap_1 TAP_8136 (  );
sky130_fd_sc_hd__tap_1 TAP_8137 (  );
sky130_fd_sc_hd__tap_1 TAP_8138 (  );
sky130_fd_sc_hd__tap_1 TAP_8139 (  );
sky130_fd_sc_hd__tap_1 TAP_814 (  );
sky130_fd_sc_hd__tap_1 TAP_8140 (  );
sky130_fd_sc_hd__tap_1 TAP_8141 (  );
sky130_fd_sc_hd__tap_1 TAP_8142 (  );
sky130_fd_sc_hd__tap_1 TAP_8143 (  );
sky130_fd_sc_hd__tap_1 TAP_8144 (  );
sky130_fd_sc_hd__tap_1 TAP_8145 (  );
sky130_fd_sc_hd__tap_1 TAP_8146 (  );
sky130_fd_sc_hd__tap_1 TAP_8147 (  );
sky130_fd_sc_hd__tap_1 TAP_8148 (  );
sky130_fd_sc_hd__tap_1 TAP_8149 (  );
sky130_fd_sc_hd__tap_1 TAP_815 (  );
sky130_fd_sc_hd__tap_1 TAP_8150 (  );
sky130_fd_sc_hd__tap_1 TAP_8151 (  );
sky130_fd_sc_hd__tap_1 TAP_8152 (  );
sky130_fd_sc_hd__tap_1 TAP_8153 (  );
sky130_fd_sc_hd__tap_1 TAP_8154 (  );
sky130_fd_sc_hd__tap_1 TAP_8155 (  );
sky130_fd_sc_hd__tap_1 TAP_8156 (  );
sky130_fd_sc_hd__tap_1 TAP_8157 (  );
sky130_fd_sc_hd__tap_1 TAP_8158 (  );
sky130_fd_sc_hd__tap_1 TAP_8159 (  );
sky130_fd_sc_hd__tap_1 TAP_816 (  );
sky130_fd_sc_hd__tap_1 TAP_8160 (  );
sky130_fd_sc_hd__tap_1 TAP_8161 (  );
sky130_fd_sc_hd__tap_1 TAP_8162 (  );
sky130_fd_sc_hd__tap_1 TAP_8163 (  );
sky130_fd_sc_hd__tap_1 TAP_8164 (  );
sky130_fd_sc_hd__tap_1 TAP_8165 (  );
sky130_fd_sc_hd__tap_1 TAP_8166 (  );
sky130_fd_sc_hd__tap_1 TAP_8167 (  );
sky130_fd_sc_hd__tap_1 TAP_8168 (  );
sky130_fd_sc_hd__tap_1 TAP_8169 (  );
sky130_fd_sc_hd__tap_1 TAP_817 (  );
sky130_fd_sc_hd__tap_1 TAP_8170 (  );
sky130_fd_sc_hd__tap_1 TAP_8171 (  );
sky130_fd_sc_hd__tap_1 TAP_8172 (  );
sky130_fd_sc_hd__tap_1 TAP_8173 (  );
sky130_fd_sc_hd__tap_1 TAP_8174 (  );
sky130_fd_sc_hd__tap_1 TAP_8175 (  );
sky130_fd_sc_hd__tap_1 TAP_8176 (  );
sky130_fd_sc_hd__tap_1 TAP_8177 (  );
sky130_fd_sc_hd__tap_1 TAP_8178 (  );
sky130_fd_sc_hd__tap_1 TAP_8179 (  );
sky130_fd_sc_hd__tap_1 TAP_818 (  );
sky130_fd_sc_hd__tap_1 TAP_8180 (  );
sky130_fd_sc_hd__tap_1 TAP_8181 (  );
sky130_fd_sc_hd__tap_1 TAP_8182 (  );
sky130_fd_sc_hd__tap_1 TAP_8183 (  );
sky130_fd_sc_hd__tap_1 TAP_8184 (  );
sky130_fd_sc_hd__tap_1 TAP_8185 (  );
sky130_fd_sc_hd__tap_1 TAP_8186 (  );
sky130_fd_sc_hd__tap_1 TAP_8187 (  );
sky130_fd_sc_hd__tap_1 TAP_8188 (  );
sky130_fd_sc_hd__tap_1 TAP_8189 (  );
sky130_fd_sc_hd__tap_1 TAP_819 (  );
sky130_fd_sc_hd__tap_1 TAP_8190 (  );
sky130_fd_sc_hd__tap_1 TAP_8191 (  );
sky130_fd_sc_hd__tap_1 TAP_8192 (  );
sky130_fd_sc_hd__tap_1 TAP_8193 (  );
sky130_fd_sc_hd__tap_1 TAP_8194 (  );
sky130_fd_sc_hd__tap_1 TAP_8195 (  );
sky130_fd_sc_hd__tap_1 TAP_8196 (  );
sky130_fd_sc_hd__tap_1 TAP_8197 (  );
sky130_fd_sc_hd__tap_1 TAP_8198 (  );
sky130_fd_sc_hd__tap_1 TAP_8199 (  );
sky130_fd_sc_hd__tap_1 TAP_820 (  );
sky130_fd_sc_hd__tap_1 TAP_8200 (  );
sky130_fd_sc_hd__tap_1 TAP_8201 (  );
sky130_fd_sc_hd__tap_1 TAP_8202 (  );
sky130_fd_sc_hd__tap_1 TAP_8203 (  );
sky130_fd_sc_hd__tap_1 TAP_8204 (  );
sky130_fd_sc_hd__tap_1 TAP_8205 (  );
sky130_fd_sc_hd__tap_1 TAP_8206 (  );
sky130_fd_sc_hd__tap_1 TAP_8207 (  );
sky130_fd_sc_hd__tap_1 TAP_8208 (  );
sky130_fd_sc_hd__tap_1 TAP_8209 (  );
sky130_fd_sc_hd__tap_1 TAP_821 (  );
sky130_fd_sc_hd__tap_1 TAP_8210 (  );
sky130_fd_sc_hd__tap_1 TAP_8211 (  );
sky130_fd_sc_hd__tap_1 TAP_8212 (  );
sky130_fd_sc_hd__tap_1 TAP_8213 (  );
sky130_fd_sc_hd__tap_1 TAP_8214 (  );
sky130_fd_sc_hd__tap_1 TAP_8215 (  );
sky130_fd_sc_hd__tap_1 TAP_8216 (  );
sky130_fd_sc_hd__tap_1 TAP_8217 (  );
sky130_fd_sc_hd__tap_1 TAP_8218 (  );
sky130_fd_sc_hd__tap_1 TAP_8219 (  );
sky130_fd_sc_hd__tap_1 TAP_822 (  );
sky130_fd_sc_hd__tap_1 TAP_8220 (  );
sky130_fd_sc_hd__tap_1 TAP_8221 (  );
sky130_fd_sc_hd__tap_1 TAP_8222 (  );
sky130_fd_sc_hd__tap_1 TAP_8223 (  );
sky130_fd_sc_hd__tap_1 TAP_8224 (  );
sky130_fd_sc_hd__tap_1 TAP_8225 (  );
sky130_fd_sc_hd__tap_1 TAP_8226 (  );
sky130_fd_sc_hd__tap_1 TAP_8227 (  );
sky130_fd_sc_hd__tap_1 TAP_8228 (  );
sky130_fd_sc_hd__tap_1 TAP_8229 (  );
sky130_fd_sc_hd__tap_1 TAP_823 (  );
sky130_fd_sc_hd__tap_1 TAP_8230 (  );
sky130_fd_sc_hd__tap_1 TAP_8231 (  );
sky130_fd_sc_hd__tap_1 TAP_8232 (  );
sky130_fd_sc_hd__tap_1 TAP_8233 (  );
sky130_fd_sc_hd__tap_1 TAP_8234 (  );
sky130_fd_sc_hd__tap_1 TAP_8235 (  );
sky130_fd_sc_hd__tap_1 TAP_8236 (  );
sky130_fd_sc_hd__tap_1 TAP_8237 (  );
sky130_fd_sc_hd__tap_1 TAP_8238 (  );
sky130_fd_sc_hd__tap_1 TAP_8239 (  );
sky130_fd_sc_hd__tap_1 TAP_824 (  );
sky130_fd_sc_hd__tap_1 TAP_8240 (  );
sky130_fd_sc_hd__tap_1 TAP_8241 (  );
sky130_fd_sc_hd__tap_1 TAP_8242 (  );
sky130_fd_sc_hd__tap_1 TAP_8243 (  );
sky130_fd_sc_hd__tap_1 TAP_8244 (  );
sky130_fd_sc_hd__tap_1 TAP_8245 (  );
sky130_fd_sc_hd__tap_1 TAP_8246 (  );
sky130_fd_sc_hd__tap_1 TAP_8247 (  );
sky130_fd_sc_hd__tap_1 TAP_8248 (  );
sky130_fd_sc_hd__tap_1 TAP_8249 (  );
sky130_fd_sc_hd__tap_1 TAP_825 (  );
sky130_fd_sc_hd__tap_1 TAP_8250 (  );
sky130_fd_sc_hd__tap_1 TAP_8251 (  );
sky130_fd_sc_hd__tap_1 TAP_8252 (  );
sky130_fd_sc_hd__tap_1 TAP_8253 (  );
sky130_fd_sc_hd__tap_1 TAP_8254 (  );
sky130_fd_sc_hd__tap_1 TAP_8255 (  );
sky130_fd_sc_hd__tap_1 TAP_8256 (  );
sky130_fd_sc_hd__tap_1 TAP_8257 (  );
sky130_fd_sc_hd__tap_1 TAP_8258 (  );
sky130_fd_sc_hd__tap_1 TAP_8259 (  );
sky130_fd_sc_hd__tap_1 TAP_826 (  );
sky130_fd_sc_hd__tap_1 TAP_8260 (  );
sky130_fd_sc_hd__tap_1 TAP_8261 (  );
sky130_fd_sc_hd__tap_1 TAP_8262 (  );
sky130_fd_sc_hd__tap_1 TAP_8263 (  );
sky130_fd_sc_hd__tap_1 TAP_8264 (  );
sky130_fd_sc_hd__tap_1 TAP_8265 (  );
sky130_fd_sc_hd__tap_1 TAP_8266 (  );
sky130_fd_sc_hd__tap_1 TAP_8267 (  );
sky130_fd_sc_hd__tap_1 TAP_8268 (  );
sky130_fd_sc_hd__tap_1 TAP_8269 (  );
sky130_fd_sc_hd__tap_1 TAP_827 (  );
sky130_fd_sc_hd__tap_1 TAP_8270 (  );
sky130_fd_sc_hd__tap_1 TAP_8271 (  );
sky130_fd_sc_hd__tap_1 TAP_8272 (  );
sky130_fd_sc_hd__tap_1 TAP_8273 (  );
sky130_fd_sc_hd__tap_1 TAP_8274 (  );
sky130_fd_sc_hd__tap_1 TAP_8275 (  );
sky130_fd_sc_hd__tap_1 TAP_8276 (  );
sky130_fd_sc_hd__tap_1 TAP_8277 (  );
sky130_fd_sc_hd__tap_1 TAP_8278 (  );
sky130_fd_sc_hd__tap_1 TAP_8279 (  );
sky130_fd_sc_hd__tap_1 TAP_828 (  );
sky130_fd_sc_hd__tap_1 TAP_8280 (  );
sky130_fd_sc_hd__tap_1 TAP_8281 (  );
sky130_fd_sc_hd__tap_1 TAP_8282 (  );
sky130_fd_sc_hd__tap_1 TAP_8283 (  );
sky130_fd_sc_hd__tap_1 TAP_8284 (  );
sky130_fd_sc_hd__tap_1 TAP_8285 (  );
sky130_fd_sc_hd__tap_1 TAP_8286 (  );
sky130_fd_sc_hd__tap_1 TAP_8287 (  );
sky130_fd_sc_hd__tap_1 TAP_8288 (  );
sky130_fd_sc_hd__tap_1 TAP_8289 (  );
sky130_fd_sc_hd__tap_1 TAP_829 (  );
sky130_fd_sc_hd__tap_1 TAP_8290 (  );
sky130_fd_sc_hd__tap_1 TAP_8291 (  );
sky130_fd_sc_hd__tap_1 TAP_8292 (  );
sky130_fd_sc_hd__tap_1 TAP_8293 (  );
sky130_fd_sc_hd__tap_1 TAP_8294 (  );
sky130_fd_sc_hd__tap_1 TAP_8295 (  );
sky130_fd_sc_hd__tap_1 TAP_8296 (  );
sky130_fd_sc_hd__tap_1 TAP_8297 (  );
sky130_fd_sc_hd__tap_1 TAP_8298 (  );
sky130_fd_sc_hd__tap_1 TAP_8299 (  );
sky130_fd_sc_hd__tap_1 TAP_830 (  );
sky130_fd_sc_hd__tap_1 TAP_8300 (  );
sky130_fd_sc_hd__tap_1 TAP_8301 (  );
sky130_fd_sc_hd__tap_1 TAP_8302 (  );
sky130_fd_sc_hd__tap_1 TAP_8303 (  );
sky130_fd_sc_hd__tap_1 TAP_8304 (  );
sky130_fd_sc_hd__tap_1 TAP_8305 (  );
sky130_fd_sc_hd__tap_1 TAP_8306 (  );
sky130_fd_sc_hd__tap_1 TAP_8307 (  );
sky130_fd_sc_hd__tap_1 TAP_8308 (  );
sky130_fd_sc_hd__tap_1 TAP_8309 (  );
sky130_fd_sc_hd__tap_1 TAP_831 (  );
sky130_fd_sc_hd__tap_1 TAP_8310 (  );
sky130_fd_sc_hd__tap_1 TAP_8311 (  );
sky130_fd_sc_hd__tap_1 TAP_8312 (  );
sky130_fd_sc_hd__tap_1 TAP_8313 (  );
sky130_fd_sc_hd__tap_1 TAP_8314 (  );
sky130_fd_sc_hd__tap_1 TAP_8315 (  );
sky130_fd_sc_hd__tap_1 TAP_8316 (  );
sky130_fd_sc_hd__tap_1 TAP_8317 (  );
sky130_fd_sc_hd__tap_1 TAP_8318 (  );
sky130_fd_sc_hd__tap_1 TAP_8319 (  );
sky130_fd_sc_hd__tap_1 TAP_832 (  );
sky130_fd_sc_hd__tap_1 TAP_8320 (  );
sky130_fd_sc_hd__tap_1 TAP_8321 (  );
sky130_fd_sc_hd__tap_1 TAP_8322 (  );
sky130_fd_sc_hd__tap_1 TAP_8323 (  );
sky130_fd_sc_hd__tap_1 TAP_8324 (  );
sky130_fd_sc_hd__tap_1 TAP_8325 (  );
sky130_fd_sc_hd__tap_1 TAP_8326 (  );
sky130_fd_sc_hd__tap_1 TAP_8327 (  );
sky130_fd_sc_hd__tap_1 TAP_8328 (  );
sky130_fd_sc_hd__tap_1 TAP_8329 (  );
sky130_fd_sc_hd__tap_1 TAP_833 (  );
sky130_fd_sc_hd__tap_1 TAP_8330 (  );
sky130_fd_sc_hd__tap_1 TAP_8331 (  );
sky130_fd_sc_hd__tap_1 TAP_8332 (  );
sky130_fd_sc_hd__tap_1 TAP_8333 (  );
sky130_fd_sc_hd__tap_1 TAP_8334 (  );
sky130_fd_sc_hd__tap_1 TAP_8335 (  );
sky130_fd_sc_hd__tap_1 TAP_8336 (  );
sky130_fd_sc_hd__tap_1 TAP_8337 (  );
sky130_fd_sc_hd__tap_1 TAP_8338 (  );
sky130_fd_sc_hd__tap_1 TAP_8339 (  );
sky130_fd_sc_hd__tap_1 TAP_834 (  );
sky130_fd_sc_hd__tap_1 TAP_8340 (  );
sky130_fd_sc_hd__tap_1 TAP_8341 (  );
sky130_fd_sc_hd__tap_1 TAP_8342 (  );
sky130_fd_sc_hd__tap_1 TAP_8343 (  );
sky130_fd_sc_hd__tap_1 TAP_8344 (  );
sky130_fd_sc_hd__tap_1 TAP_8345 (  );
sky130_fd_sc_hd__tap_1 TAP_8346 (  );
sky130_fd_sc_hd__tap_1 TAP_8347 (  );
sky130_fd_sc_hd__tap_1 TAP_8348 (  );
sky130_fd_sc_hd__tap_1 TAP_8349 (  );
sky130_fd_sc_hd__tap_1 TAP_835 (  );
sky130_fd_sc_hd__tap_1 TAP_8350 (  );
sky130_fd_sc_hd__tap_1 TAP_8351 (  );
sky130_fd_sc_hd__tap_1 TAP_8352 (  );
sky130_fd_sc_hd__tap_1 TAP_8353 (  );
sky130_fd_sc_hd__tap_1 TAP_8354 (  );
sky130_fd_sc_hd__tap_1 TAP_8355 (  );
sky130_fd_sc_hd__tap_1 TAP_8356 (  );
sky130_fd_sc_hd__tap_1 TAP_8357 (  );
sky130_fd_sc_hd__tap_1 TAP_8358 (  );
sky130_fd_sc_hd__tap_1 TAP_8359 (  );
sky130_fd_sc_hd__tap_1 TAP_836 (  );
sky130_fd_sc_hd__tap_1 TAP_8360 (  );
sky130_fd_sc_hd__tap_1 TAP_8361 (  );
sky130_fd_sc_hd__tap_1 TAP_8362 (  );
sky130_fd_sc_hd__tap_1 TAP_8363 (  );
sky130_fd_sc_hd__tap_1 TAP_8364 (  );
sky130_fd_sc_hd__tap_1 TAP_8365 (  );
sky130_fd_sc_hd__tap_1 TAP_8366 (  );
sky130_fd_sc_hd__tap_1 TAP_8367 (  );
sky130_fd_sc_hd__tap_1 TAP_8368 (  );
sky130_fd_sc_hd__tap_1 TAP_8369 (  );
sky130_fd_sc_hd__tap_1 TAP_837 (  );
sky130_fd_sc_hd__tap_1 TAP_8370 (  );
sky130_fd_sc_hd__tap_1 TAP_8371 (  );
sky130_fd_sc_hd__tap_1 TAP_8372 (  );
sky130_fd_sc_hd__tap_1 TAP_8373 (  );
sky130_fd_sc_hd__tap_1 TAP_8374 (  );
sky130_fd_sc_hd__tap_1 TAP_8375 (  );
sky130_fd_sc_hd__tap_1 TAP_8376 (  );
sky130_fd_sc_hd__tap_1 TAP_8377 (  );
sky130_fd_sc_hd__tap_1 TAP_8378 (  );
sky130_fd_sc_hd__tap_1 TAP_8379 (  );
sky130_fd_sc_hd__tap_1 TAP_838 (  );
sky130_fd_sc_hd__tap_1 TAP_8380 (  );
sky130_fd_sc_hd__tap_1 TAP_8381 (  );
sky130_fd_sc_hd__tap_1 TAP_8382 (  );
sky130_fd_sc_hd__tap_1 TAP_8383 (  );
sky130_fd_sc_hd__tap_1 TAP_8384 (  );
sky130_fd_sc_hd__tap_1 TAP_8385 (  );
sky130_fd_sc_hd__tap_1 TAP_8386 (  );
sky130_fd_sc_hd__tap_1 TAP_8387 (  );
sky130_fd_sc_hd__tap_1 TAP_8388 (  );
sky130_fd_sc_hd__tap_1 TAP_8389 (  );
sky130_fd_sc_hd__tap_1 TAP_839 (  );
sky130_fd_sc_hd__tap_1 TAP_8390 (  );
sky130_fd_sc_hd__tap_1 TAP_8391 (  );
sky130_fd_sc_hd__tap_1 TAP_8392 (  );
sky130_fd_sc_hd__tap_1 TAP_8393 (  );
sky130_fd_sc_hd__tap_1 TAP_8394 (  );
sky130_fd_sc_hd__tap_1 TAP_8395 (  );
sky130_fd_sc_hd__tap_1 TAP_8396 (  );
sky130_fd_sc_hd__tap_1 TAP_8397 (  );
sky130_fd_sc_hd__tap_1 TAP_8398 (  );
sky130_fd_sc_hd__tap_1 TAP_8399 (  );
sky130_fd_sc_hd__tap_1 TAP_840 (  );
sky130_fd_sc_hd__tap_1 TAP_8400 (  );
sky130_fd_sc_hd__tap_1 TAP_8401 (  );
sky130_fd_sc_hd__tap_1 TAP_8402 (  );
sky130_fd_sc_hd__tap_1 TAP_8403 (  );
sky130_fd_sc_hd__tap_1 TAP_8404 (  );
sky130_fd_sc_hd__tap_1 TAP_8405 (  );
sky130_fd_sc_hd__tap_1 TAP_8406 (  );
sky130_fd_sc_hd__tap_1 TAP_8407 (  );
sky130_fd_sc_hd__tap_1 TAP_8408 (  );
sky130_fd_sc_hd__tap_1 TAP_8409 (  );
sky130_fd_sc_hd__tap_1 TAP_841 (  );
sky130_fd_sc_hd__tap_1 TAP_8410 (  );
sky130_fd_sc_hd__tap_1 TAP_8411 (  );
sky130_fd_sc_hd__tap_1 TAP_8412 (  );
sky130_fd_sc_hd__tap_1 TAP_8413 (  );
sky130_fd_sc_hd__tap_1 TAP_8414 (  );
sky130_fd_sc_hd__tap_1 TAP_8415 (  );
sky130_fd_sc_hd__tap_1 TAP_8416 (  );
sky130_fd_sc_hd__tap_1 TAP_8417 (  );
sky130_fd_sc_hd__tap_1 TAP_8418 (  );
sky130_fd_sc_hd__tap_1 TAP_8419 (  );
sky130_fd_sc_hd__tap_1 TAP_842 (  );
sky130_fd_sc_hd__tap_1 TAP_8420 (  );
sky130_fd_sc_hd__tap_1 TAP_8421 (  );
sky130_fd_sc_hd__tap_1 TAP_8422 (  );
sky130_fd_sc_hd__tap_1 TAP_8423 (  );
sky130_fd_sc_hd__tap_1 TAP_8424 (  );
sky130_fd_sc_hd__tap_1 TAP_8425 (  );
sky130_fd_sc_hd__tap_1 TAP_8426 (  );
sky130_fd_sc_hd__tap_1 TAP_8427 (  );
sky130_fd_sc_hd__tap_1 TAP_8428 (  );
sky130_fd_sc_hd__tap_1 TAP_8429 (  );
sky130_fd_sc_hd__tap_1 TAP_843 (  );
sky130_fd_sc_hd__tap_1 TAP_8430 (  );
sky130_fd_sc_hd__tap_1 TAP_8431 (  );
sky130_fd_sc_hd__tap_1 TAP_8432 (  );
sky130_fd_sc_hd__tap_1 TAP_8433 (  );
sky130_fd_sc_hd__tap_1 TAP_8434 (  );
sky130_fd_sc_hd__tap_1 TAP_8435 (  );
sky130_fd_sc_hd__tap_1 TAP_8436 (  );
sky130_fd_sc_hd__tap_1 TAP_8437 (  );
sky130_fd_sc_hd__tap_1 TAP_8438 (  );
sky130_fd_sc_hd__tap_1 TAP_8439 (  );
sky130_fd_sc_hd__tap_1 TAP_844 (  );
sky130_fd_sc_hd__tap_1 TAP_8440 (  );
sky130_fd_sc_hd__tap_1 TAP_8441 (  );
sky130_fd_sc_hd__tap_1 TAP_8442 (  );
sky130_fd_sc_hd__tap_1 TAP_8443 (  );
sky130_fd_sc_hd__tap_1 TAP_8444 (  );
sky130_fd_sc_hd__tap_1 TAP_8445 (  );
sky130_fd_sc_hd__tap_1 TAP_8446 (  );
sky130_fd_sc_hd__tap_1 TAP_8447 (  );
sky130_fd_sc_hd__tap_1 TAP_8448 (  );
sky130_fd_sc_hd__tap_1 TAP_8449 (  );
sky130_fd_sc_hd__tap_1 TAP_845 (  );
sky130_fd_sc_hd__tap_1 TAP_8450 (  );
sky130_fd_sc_hd__tap_1 TAP_8451 (  );
sky130_fd_sc_hd__tap_1 TAP_8452 (  );
sky130_fd_sc_hd__tap_1 TAP_8453 (  );
sky130_fd_sc_hd__tap_1 TAP_8454 (  );
sky130_fd_sc_hd__tap_1 TAP_8455 (  );
sky130_fd_sc_hd__tap_1 TAP_8456 (  );
sky130_fd_sc_hd__tap_1 TAP_8457 (  );
sky130_fd_sc_hd__tap_1 TAP_8458 (  );
sky130_fd_sc_hd__tap_1 TAP_8459 (  );
sky130_fd_sc_hd__tap_1 TAP_846 (  );
sky130_fd_sc_hd__tap_1 TAP_8460 (  );
sky130_fd_sc_hd__tap_1 TAP_8461 (  );
sky130_fd_sc_hd__tap_1 TAP_8462 (  );
sky130_fd_sc_hd__tap_1 TAP_8463 (  );
sky130_fd_sc_hd__tap_1 TAP_8464 (  );
sky130_fd_sc_hd__tap_1 TAP_8465 (  );
sky130_fd_sc_hd__tap_1 TAP_8466 (  );
sky130_fd_sc_hd__tap_1 TAP_8467 (  );
sky130_fd_sc_hd__tap_1 TAP_8468 (  );
sky130_fd_sc_hd__tap_1 TAP_8469 (  );
sky130_fd_sc_hd__tap_1 TAP_847 (  );
sky130_fd_sc_hd__tap_1 TAP_8470 (  );
sky130_fd_sc_hd__tap_1 TAP_8471 (  );
sky130_fd_sc_hd__tap_1 TAP_8472 (  );
sky130_fd_sc_hd__tap_1 TAP_8473 (  );
sky130_fd_sc_hd__tap_1 TAP_8474 (  );
sky130_fd_sc_hd__tap_1 TAP_8475 (  );
sky130_fd_sc_hd__tap_1 TAP_8476 (  );
sky130_fd_sc_hd__tap_1 TAP_8477 (  );
sky130_fd_sc_hd__tap_1 TAP_8478 (  );
sky130_fd_sc_hd__tap_1 TAP_8479 (  );
sky130_fd_sc_hd__tap_1 TAP_848 (  );
sky130_fd_sc_hd__tap_1 TAP_8480 (  );
sky130_fd_sc_hd__tap_1 TAP_8481 (  );
sky130_fd_sc_hd__tap_1 TAP_8482 (  );
sky130_fd_sc_hd__tap_1 TAP_8483 (  );
sky130_fd_sc_hd__tap_1 TAP_8484 (  );
sky130_fd_sc_hd__tap_1 TAP_8485 (  );
sky130_fd_sc_hd__tap_1 TAP_8486 (  );
sky130_fd_sc_hd__tap_1 TAP_8487 (  );
sky130_fd_sc_hd__tap_1 TAP_8488 (  );
sky130_fd_sc_hd__tap_1 TAP_8489 (  );
sky130_fd_sc_hd__tap_1 TAP_849 (  );
sky130_fd_sc_hd__tap_1 TAP_8490 (  );
sky130_fd_sc_hd__tap_1 TAP_8491 (  );
sky130_fd_sc_hd__tap_1 TAP_8492 (  );
sky130_fd_sc_hd__tap_1 TAP_8493 (  );
sky130_fd_sc_hd__tap_1 TAP_8494 (  );
sky130_fd_sc_hd__tap_1 TAP_8495 (  );
sky130_fd_sc_hd__tap_1 TAP_8496 (  );
sky130_fd_sc_hd__tap_1 TAP_8497 (  );
sky130_fd_sc_hd__tap_1 TAP_8498 (  );
sky130_fd_sc_hd__tap_1 TAP_8499 (  );
sky130_fd_sc_hd__tap_1 TAP_850 (  );
sky130_fd_sc_hd__tap_1 TAP_8500 (  );
sky130_fd_sc_hd__tap_1 TAP_8501 (  );
sky130_fd_sc_hd__tap_1 TAP_8502 (  );
sky130_fd_sc_hd__tap_1 TAP_8503 (  );
sky130_fd_sc_hd__tap_1 TAP_8504 (  );
sky130_fd_sc_hd__tap_1 TAP_8505 (  );
sky130_fd_sc_hd__tap_1 TAP_8506 (  );
sky130_fd_sc_hd__tap_1 TAP_8507 (  );
sky130_fd_sc_hd__tap_1 TAP_8508 (  );
sky130_fd_sc_hd__tap_1 TAP_8509 (  );
sky130_fd_sc_hd__tap_1 TAP_851 (  );
sky130_fd_sc_hd__tap_1 TAP_8510 (  );
sky130_fd_sc_hd__tap_1 TAP_8511 (  );
sky130_fd_sc_hd__tap_1 TAP_8512 (  );
sky130_fd_sc_hd__tap_1 TAP_8513 (  );
sky130_fd_sc_hd__tap_1 TAP_8514 (  );
sky130_fd_sc_hd__tap_1 TAP_8515 (  );
sky130_fd_sc_hd__tap_1 TAP_8516 (  );
sky130_fd_sc_hd__tap_1 TAP_8517 (  );
sky130_fd_sc_hd__tap_1 TAP_8518 (  );
sky130_fd_sc_hd__tap_1 TAP_8519 (  );
sky130_fd_sc_hd__tap_1 TAP_852 (  );
sky130_fd_sc_hd__tap_1 TAP_8520 (  );
sky130_fd_sc_hd__tap_1 TAP_8521 (  );
sky130_fd_sc_hd__tap_1 TAP_8522 (  );
sky130_fd_sc_hd__tap_1 TAP_8523 (  );
sky130_fd_sc_hd__tap_1 TAP_8524 (  );
sky130_fd_sc_hd__tap_1 TAP_8525 (  );
sky130_fd_sc_hd__tap_1 TAP_8526 (  );
sky130_fd_sc_hd__tap_1 TAP_8527 (  );
sky130_fd_sc_hd__tap_1 TAP_8528 (  );
sky130_fd_sc_hd__tap_1 TAP_8529 (  );
sky130_fd_sc_hd__tap_1 TAP_853 (  );
sky130_fd_sc_hd__tap_1 TAP_8530 (  );
sky130_fd_sc_hd__tap_1 TAP_8531 (  );
sky130_fd_sc_hd__tap_1 TAP_8532 (  );
sky130_fd_sc_hd__tap_1 TAP_8533 (  );
sky130_fd_sc_hd__tap_1 TAP_8534 (  );
sky130_fd_sc_hd__tap_1 TAP_8535 (  );
sky130_fd_sc_hd__tap_1 TAP_8536 (  );
sky130_fd_sc_hd__tap_1 TAP_8537 (  );
sky130_fd_sc_hd__tap_1 TAP_8538 (  );
sky130_fd_sc_hd__tap_1 TAP_8539 (  );
sky130_fd_sc_hd__tap_1 TAP_854 (  );
sky130_fd_sc_hd__tap_1 TAP_8540 (  );
sky130_fd_sc_hd__tap_1 TAP_8541 (  );
sky130_fd_sc_hd__tap_1 TAP_8542 (  );
sky130_fd_sc_hd__tap_1 TAP_8543 (  );
sky130_fd_sc_hd__tap_1 TAP_8544 (  );
sky130_fd_sc_hd__tap_1 TAP_8545 (  );
sky130_fd_sc_hd__tap_1 TAP_8546 (  );
sky130_fd_sc_hd__tap_1 TAP_8547 (  );
sky130_fd_sc_hd__tap_1 TAP_8548 (  );
sky130_fd_sc_hd__tap_1 TAP_8549 (  );
sky130_fd_sc_hd__tap_1 TAP_855 (  );
sky130_fd_sc_hd__tap_1 TAP_8550 (  );
sky130_fd_sc_hd__tap_1 TAP_8551 (  );
sky130_fd_sc_hd__tap_1 TAP_8552 (  );
sky130_fd_sc_hd__tap_1 TAP_8553 (  );
sky130_fd_sc_hd__tap_1 TAP_8554 (  );
sky130_fd_sc_hd__tap_1 TAP_8555 (  );
sky130_fd_sc_hd__tap_1 TAP_8556 (  );
sky130_fd_sc_hd__tap_1 TAP_8557 (  );
sky130_fd_sc_hd__tap_1 TAP_8558 (  );
sky130_fd_sc_hd__tap_1 TAP_8559 (  );
sky130_fd_sc_hd__tap_1 TAP_856 (  );
sky130_fd_sc_hd__tap_1 TAP_8560 (  );
sky130_fd_sc_hd__tap_1 TAP_8561 (  );
sky130_fd_sc_hd__tap_1 TAP_8562 (  );
sky130_fd_sc_hd__tap_1 TAP_8563 (  );
sky130_fd_sc_hd__tap_1 TAP_8564 (  );
sky130_fd_sc_hd__tap_1 TAP_8565 (  );
sky130_fd_sc_hd__tap_1 TAP_8566 (  );
sky130_fd_sc_hd__tap_1 TAP_8567 (  );
sky130_fd_sc_hd__tap_1 TAP_8568 (  );
sky130_fd_sc_hd__tap_1 TAP_8569 (  );
sky130_fd_sc_hd__tap_1 TAP_857 (  );
sky130_fd_sc_hd__tap_1 TAP_8570 (  );
sky130_fd_sc_hd__tap_1 TAP_8571 (  );
sky130_fd_sc_hd__tap_1 TAP_8572 (  );
sky130_fd_sc_hd__tap_1 TAP_8573 (  );
sky130_fd_sc_hd__tap_1 TAP_8574 (  );
sky130_fd_sc_hd__tap_1 TAP_8575 (  );
sky130_fd_sc_hd__tap_1 TAP_8576 (  );
sky130_fd_sc_hd__tap_1 TAP_8577 (  );
sky130_fd_sc_hd__tap_1 TAP_8578 (  );
sky130_fd_sc_hd__tap_1 TAP_8579 (  );
sky130_fd_sc_hd__tap_1 TAP_858 (  );
sky130_fd_sc_hd__tap_1 TAP_8580 (  );
sky130_fd_sc_hd__tap_1 TAP_8581 (  );
sky130_fd_sc_hd__tap_1 TAP_8582 (  );
sky130_fd_sc_hd__tap_1 TAP_8583 (  );
sky130_fd_sc_hd__tap_1 TAP_8584 (  );
sky130_fd_sc_hd__tap_1 TAP_8585 (  );
sky130_fd_sc_hd__tap_1 TAP_8586 (  );
sky130_fd_sc_hd__tap_1 TAP_8587 (  );
sky130_fd_sc_hd__tap_1 TAP_8588 (  );
sky130_fd_sc_hd__tap_1 TAP_8589 (  );
sky130_fd_sc_hd__tap_1 TAP_859 (  );
sky130_fd_sc_hd__tap_1 TAP_8590 (  );
sky130_fd_sc_hd__tap_1 TAP_8591 (  );
sky130_fd_sc_hd__tap_1 TAP_8592 (  );
sky130_fd_sc_hd__tap_1 TAP_8593 (  );
sky130_fd_sc_hd__tap_1 TAP_8594 (  );
sky130_fd_sc_hd__tap_1 TAP_8595 (  );
sky130_fd_sc_hd__tap_1 TAP_8596 (  );
sky130_fd_sc_hd__tap_1 TAP_8597 (  );
sky130_fd_sc_hd__tap_1 TAP_8598 (  );
sky130_fd_sc_hd__tap_1 TAP_8599 (  );
sky130_fd_sc_hd__tap_1 TAP_860 (  );
sky130_fd_sc_hd__tap_1 TAP_8600 (  );
sky130_fd_sc_hd__tap_1 TAP_8601 (  );
sky130_fd_sc_hd__tap_1 TAP_8602 (  );
sky130_fd_sc_hd__tap_1 TAP_8603 (  );
sky130_fd_sc_hd__tap_1 TAP_8604 (  );
sky130_fd_sc_hd__tap_1 TAP_8605 (  );
sky130_fd_sc_hd__tap_1 TAP_8606 (  );
sky130_fd_sc_hd__tap_1 TAP_8607 (  );
sky130_fd_sc_hd__tap_1 TAP_8608 (  );
sky130_fd_sc_hd__tap_1 TAP_8609 (  );
sky130_fd_sc_hd__tap_1 TAP_861 (  );
sky130_fd_sc_hd__tap_1 TAP_8610 (  );
sky130_fd_sc_hd__tap_1 TAP_8611 (  );
sky130_fd_sc_hd__tap_1 TAP_8612 (  );
sky130_fd_sc_hd__tap_1 TAP_8613 (  );
sky130_fd_sc_hd__tap_1 TAP_8614 (  );
sky130_fd_sc_hd__tap_1 TAP_8615 (  );
sky130_fd_sc_hd__tap_1 TAP_8616 (  );
sky130_fd_sc_hd__tap_1 TAP_8617 (  );
sky130_fd_sc_hd__tap_1 TAP_8618 (  );
sky130_fd_sc_hd__tap_1 TAP_8619 (  );
sky130_fd_sc_hd__tap_1 TAP_862 (  );
sky130_fd_sc_hd__tap_1 TAP_8620 (  );
sky130_fd_sc_hd__tap_1 TAP_8621 (  );
sky130_fd_sc_hd__tap_1 TAP_8622 (  );
sky130_fd_sc_hd__tap_1 TAP_8623 (  );
sky130_fd_sc_hd__tap_1 TAP_8624 (  );
sky130_fd_sc_hd__tap_1 TAP_8625 (  );
sky130_fd_sc_hd__tap_1 TAP_8626 (  );
sky130_fd_sc_hd__tap_1 TAP_8627 (  );
sky130_fd_sc_hd__tap_1 TAP_8628 (  );
sky130_fd_sc_hd__tap_1 TAP_8629 (  );
sky130_fd_sc_hd__tap_1 TAP_863 (  );
sky130_fd_sc_hd__tap_1 TAP_8630 (  );
sky130_fd_sc_hd__tap_1 TAP_8631 (  );
sky130_fd_sc_hd__tap_1 TAP_8632 (  );
sky130_fd_sc_hd__tap_1 TAP_8633 (  );
sky130_fd_sc_hd__tap_1 TAP_8634 (  );
sky130_fd_sc_hd__tap_1 TAP_8635 (  );
sky130_fd_sc_hd__tap_1 TAP_8636 (  );
sky130_fd_sc_hd__tap_1 TAP_8637 (  );
sky130_fd_sc_hd__tap_1 TAP_8638 (  );
sky130_fd_sc_hd__tap_1 TAP_8639 (  );
sky130_fd_sc_hd__tap_1 TAP_864 (  );
sky130_fd_sc_hd__tap_1 TAP_8640 (  );
sky130_fd_sc_hd__tap_1 TAP_8641 (  );
sky130_fd_sc_hd__tap_1 TAP_8642 (  );
sky130_fd_sc_hd__tap_1 TAP_8643 (  );
sky130_fd_sc_hd__tap_1 TAP_8644 (  );
sky130_fd_sc_hd__tap_1 TAP_8645 (  );
sky130_fd_sc_hd__tap_1 TAP_8646 (  );
sky130_fd_sc_hd__tap_1 TAP_8647 (  );
sky130_fd_sc_hd__tap_1 TAP_8648 (  );
sky130_fd_sc_hd__tap_1 TAP_8649 (  );
sky130_fd_sc_hd__tap_1 TAP_865 (  );
sky130_fd_sc_hd__tap_1 TAP_8650 (  );
sky130_fd_sc_hd__tap_1 TAP_8651 (  );
sky130_fd_sc_hd__tap_1 TAP_8652 (  );
sky130_fd_sc_hd__tap_1 TAP_8653 (  );
sky130_fd_sc_hd__tap_1 TAP_8654 (  );
sky130_fd_sc_hd__tap_1 TAP_8655 (  );
sky130_fd_sc_hd__tap_1 TAP_8656 (  );
sky130_fd_sc_hd__tap_1 TAP_8657 (  );
sky130_fd_sc_hd__tap_1 TAP_8658 (  );
sky130_fd_sc_hd__tap_1 TAP_8659 (  );
sky130_fd_sc_hd__tap_1 TAP_866 (  );
sky130_fd_sc_hd__tap_1 TAP_8660 (  );
sky130_fd_sc_hd__tap_1 TAP_8661 (  );
sky130_fd_sc_hd__tap_1 TAP_8662 (  );
sky130_fd_sc_hd__tap_1 TAP_8663 (  );
sky130_fd_sc_hd__tap_1 TAP_8664 (  );
sky130_fd_sc_hd__tap_1 TAP_8665 (  );
sky130_fd_sc_hd__tap_1 TAP_8666 (  );
sky130_fd_sc_hd__tap_1 TAP_8667 (  );
sky130_fd_sc_hd__tap_1 TAP_8668 (  );
sky130_fd_sc_hd__tap_1 TAP_8669 (  );
sky130_fd_sc_hd__tap_1 TAP_867 (  );
sky130_fd_sc_hd__tap_1 TAP_8670 (  );
sky130_fd_sc_hd__tap_1 TAP_8671 (  );
sky130_fd_sc_hd__tap_1 TAP_8672 (  );
sky130_fd_sc_hd__tap_1 TAP_8673 (  );
sky130_fd_sc_hd__tap_1 TAP_8674 (  );
sky130_fd_sc_hd__tap_1 TAP_8675 (  );
sky130_fd_sc_hd__tap_1 TAP_8676 (  );
sky130_fd_sc_hd__tap_1 TAP_8677 (  );
sky130_fd_sc_hd__tap_1 TAP_8678 (  );
sky130_fd_sc_hd__tap_1 TAP_8679 (  );
sky130_fd_sc_hd__tap_1 TAP_868 (  );
sky130_fd_sc_hd__tap_1 TAP_8680 (  );
sky130_fd_sc_hd__tap_1 TAP_8681 (  );
sky130_fd_sc_hd__tap_1 TAP_8682 (  );
sky130_fd_sc_hd__tap_1 TAP_8683 (  );
sky130_fd_sc_hd__tap_1 TAP_8684 (  );
sky130_fd_sc_hd__tap_1 TAP_8685 (  );
sky130_fd_sc_hd__tap_1 TAP_8686 (  );
sky130_fd_sc_hd__tap_1 TAP_8687 (  );
sky130_fd_sc_hd__tap_1 TAP_8688 (  );
sky130_fd_sc_hd__tap_1 TAP_8689 (  );
sky130_fd_sc_hd__tap_1 TAP_869 (  );
sky130_fd_sc_hd__tap_1 TAP_8690 (  );
sky130_fd_sc_hd__tap_1 TAP_8691 (  );
sky130_fd_sc_hd__tap_1 TAP_8692 (  );
sky130_fd_sc_hd__tap_1 TAP_8693 (  );
sky130_fd_sc_hd__tap_1 TAP_8694 (  );
sky130_fd_sc_hd__tap_1 TAP_8695 (  );
sky130_fd_sc_hd__tap_1 TAP_8696 (  );
sky130_fd_sc_hd__tap_1 TAP_8697 (  );
sky130_fd_sc_hd__tap_1 TAP_8698 (  );
sky130_fd_sc_hd__tap_1 TAP_8699 (  );
sky130_fd_sc_hd__tap_1 TAP_870 (  );
sky130_fd_sc_hd__tap_1 TAP_8700 (  );
sky130_fd_sc_hd__tap_1 TAP_8701 (  );
sky130_fd_sc_hd__tap_1 TAP_8702 (  );
sky130_fd_sc_hd__tap_1 TAP_8703 (  );
sky130_fd_sc_hd__tap_1 TAP_8704 (  );
sky130_fd_sc_hd__tap_1 TAP_8705 (  );
sky130_fd_sc_hd__tap_1 TAP_8706 (  );
sky130_fd_sc_hd__tap_1 TAP_8707 (  );
sky130_fd_sc_hd__tap_1 TAP_8708 (  );
sky130_fd_sc_hd__tap_1 TAP_8709 (  );
sky130_fd_sc_hd__tap_1 TAP_871 (  );
sky130_fd_sc_hd__tap_1 TAP_8710 (  );
sky130_fd_sc_hd__tap_1 TAP_8711 (  );
sky130_fd_sc_hd__tap_1 TAP_8712 (  );
sky130_fd_sc_hd__tap_1 TAP_8713 (  );
sky130_fd_sc_hd__tap_1 TAP_8714 (  );
sky130_fd_sc_hd__tap_1 TAP_8715 (  );
sky130_fd_sc_hd__tap_1 TAP_8716 (  );
sky130_fd_sc_hd__tap_1 TAP_8717 (  );
sky130_fd_sc_hd__tap_1 TAP_8718 (  );
sky130_fd_sc_hd__tap_1 TAP_8719 (  );
sky130_fd_sc_hd__tap_1 TAP_872 (  );
sky130_fd_sc_hd__tap_1 TAP_8720 (  );
sky130_fd_sc_hd__tap_1 TAP_8721 (  );
sky130_fd_sc_hd__tap_1 TAP_8722 (  );
sky130_fd_sc_hd__tap_1 TAP_8723 (  );
sky130_fd_sc_hd__tap_1 TAP_8724 (  );
sky130_fd_sc_hd__tap_1 TAP_8725 (  );
sky130_fd_sc_hd__tap_1 TAP_8726 (  );
sky130_fd_sc_hd__tap_1 TAP_8727 (  );
sky130_fd_sc_hd__tap_1 TAP_8728 (  );
sky130_fd_sc_hd__tap_1 TAP_8729 (  );
sky130_fd_sc_hd__tap_1 TAP_873 (  );
sky130_fd_sc_hd__tap_1 TAP_8730 (  );
sky130_fd_sc_hd__tap_1 TAP_8731 (  );
sky130_fd_sc_hd__tap_1 TAP_8732 (  );
sky130_fd_sc_hd__tap_1 TAP_8733 (  );
sky130_fd_sc_hd__tap_1 TAP_8734 (  );
sky130_fd_sc_hd__tap_1 TAP_8735 (  );
sky130_fd_sc_hd__tap_1 TAP_8736 (  );
sky130_fd_sc_hd__tap_1 TAP_8737 (  );
sky130_fd_sc_hd__tap_1 TAP_8738 (  );
sky130_fd_sc_hd__tap_1 TAP_8739 (  );
sky130_fd_sc_hd__tap_1 TAP_874 (  );
sky130_fd_sc_hd__tap_1 TAP_8740 (  );
sky130_fd_sc_hd__tap_1 TAP_8741 (  );
sky130_fd_sc_hd__tap_1 TAP_8742 (  );
sky130_fd_sc_hd__tap_1 TAP_8743 (  );
sky130_fd_sc_hd__tap_1 TAP_8744 (  );
sky130_fd_sc_hd__tap_1 TAP_8745 (  );
sky130_fd_sc_hd__tap_1 TAP_8746 (  );
sky130_fd_sc_hd__tap_1 TAP_8747 (  );
sky130_fd_sc_hd__tap_1 TAP_8748 (  );
sky130_fd_sc_hd__tap_1 TAP_8749 (  );
sky130_fd_sc_hd__tap_1 TAP_875 (  );
sky130_fd_sc_hd__tap_1 TAP_8750 (  );
sky130_fd_sc_hd__tap_1 TAP_8751 (  );
sky130_fd_sc_hd__tap_1 TAP_8752 (  );
sky130_fd_sc_hd__tap_1 TAP_8753 (  );
sky130_fd_sc_hd__tap_1 TAP_8754 (  );
sky130_fd_sc_hd__tap_1 TAP_8755 (  );
sky130_fd_sc_hd__tap_1 TAP_8756 (  );
sky130_fd_sc_hd__tap_1 TAP_8757 (  );
sky130_fd_sc_hd__tap_1 TAP_8758 (  );
sky130_fd_sc_hd__tap_1 TAP_8759 (  );
sky130_fd_sc_hd__tap_1 TAP_876 (  );
sky130_fd_sc_hd__tap_1 TAP_8760 (  );
sky130_fd_sc_hd__tap_1 TAP_8761 (  );
sky130_fd_sc_hd__tap_1 TAP_8762 (  );
sky130_fd_sc_hd__tap_1 TAP_8763 (  );
sky130_fd_sc_hd__tap_1 TAP_8764 (  );
sky130_fd_sc_hd__tap_1 TAP_8765 (  );
sky130_fd_sc_hd__tap_1 TAP_8766 (  );
sky130_fd_sc_hd__tap_1 TAP_8767 (  );
sky130_fd_sc_hd__tap_1 TAP_8768 (  );
sky130_fd_sc_hd__tap_1 TAP_8769 (  );
sky130_fd_sc_hd__tap_1 TAP_877 (  );
sky130_fd_sc_hd__tap_1 TAP_8770 (  );
sky130_fd_sc_hd__tap_1 TAP_8771 (  );
sky130_fd_sc_hd__tap_1 TAP_8772 (  );
sky130_fd_sc_hd__tap_1 TAP_8773 (  );
sky130_fd_sc_hd__tap_1 TAP_8774 (  );
sky130_fd_sc_hd__tap_1 TAP_8775 (  );
sky130_fd_sc_hd__tap_1 TAP_8776 (  );
sky130_fd_sc_hd__tap_1 TAP_8777 (  );
sky130_fd_sc_hd__tap_1 TAP_8778 (  );
sky130_fd_sc_hd__tap_1 TAP_8779 (  );
sky130_fd_sc_hd__tap_1 TAP_878 (  );
sky130_fd_sc_hd__tap_1 TAP_8780 (  );
sky130_fd_sc_hd__tap_1 TAP_8781 (  );
sky130_fd_sc_hd__tap_1 TAP_8782 (  );
sky130_fd_sc_hd__tap_1 TAP_8783 (  );
sky130_fd_sc_hd__tap_1 TAP_8784 (  );
sky130_fd_sc_hd__tap_1 TAP_8785 (  );
sky130_fd_sc_hd__tap_1 TAP_8786 (  );
sky130_fd_sc_hd__tap_1 TAP_8787 (  );
sky130_fd_sc_hd__tap_1 TAP_8788 (  );
sky130_fd_sc_hd__tap_1 TAP_8789 (  );
sky130_fd_sc_hd__tap_1 TAP_879 (  );
sky130_fd_sc_hd__tap_1 TAP_8790 (  );
sky130_fd_sc_hd__tap_1 TAP_8791 (  );
sky130_fd_sc_hd__tap_1 TAP_8792 (  );
sky130_fd_sc_hd__tap_1 TAP_8793 (  );
sky130_fd_sc_hd__tap_1 TAP_8794 (  );
sky130_fd_sc_hd__tap_1 TAP_8795 (  );
sky130_fd_sc_hd__tap_1 TAP_8796 (  );
sky130_fd_sc_hd__tap_1 TAP_8797 (  );
sky130_fd_sc_hd__tap_1 TAP_8798 (  );
sky130_fd_sc_hd__tap_1 TAP_8799 (  );
sky130_fd_sc_hd__tap_1 TAP_880 (  );
sky130_fd_sc_hd__tap_1 TAP_8800 (  );
sky130_fd_sc_hd__tap_1 TAP_8801 (  );
sky130_fd_sc_hd__tap_1 TAP_8802 (  );
sky130_fd_sc_hd__tap_1 TAP_8803 (  );
sky130_fd_sc_hd__tap_1 TAP_8804 (  );
sky130_fd_sc_hd__tap_1 TAP_8805 (  );
sky130_fd_sc_hd__tap_1 TAP_8806 (  );
sky130_fd_sc_hd__tap_1 TAP_8807 (  );
sky130_fd_sc_hd__tap_1 TAP_8808 (  );
sky130_fd_sc_hd__tap_1 TAP_8809 (  );
sky130_fd_sc_hd__tap_1 TAP_881 (  );
sky130_fd_sc_hd__tap_1 TAP_8810 (  );
sky130_fd_sc_hd__tap_1 TAP_8811 (  );
sky130_fd_sc_hd__tap_1 TAP_8812 (  );
sky130_fd_sc_hd__tap_1 TAP_8813 (  );
sky130_fd_sc_hd__tap_1 TAP_8814 (  );
sky130_fd_sc_hd__tap_1 TAP_8815 (  );
sky130_fd_sc_hd__tap_1 TAP_8816 (  );
sky130_fd_sc_hd__tap_1 TAP_8817 (  );
sky130_fd_sc_hd__tap_1 TAP_8818 (  );
sky130_fd_sc_hd__tap_1 TAP_8819 (  );
sky130_fd_sc_hd__tap_1 TAP_882 (  );
sky130_fd_sc_hd__tap_1 TAP_8820 (  );
sky130_fd_sc_hd__tap_1 TAP_8821 (  );
sky130_fd_sc_hd__tap_1 TAP_8822 (  );
sky130_fd_sc_hd__tap_1 TAP_8823 (  );
sky130_fd_sc_hd__tap_1 TAP_8824 (  );
sky130_fd_sc_hd__tap_1 TAP_8825 (  );
sky130_fd_sc_hd__tap_1 TAP_8826 (  );
sky130_fd_sc_hd__tap_1 TAP_8827 (  );
sky130_fd_sc_hd__tap_1 TAP_8828 (  );
sky130_fd_sc_hd__tap_1 TAP_8829 (  );
sky130_fd_sc_hd__tap_1 TAP_883 (  );
sky130_fd_sc_hd__tap_1 TAP_8830 (  );
sky130_fd_sc_hd__tap_1 TAP_8831 (  );
sky130_fd_sc_hd__tap_1 TAP_8832 (  );
sky130_fd_sc_hd__tap_1 TAP_8833 (  );
sky130_fd_sc_hd__tap_1 TAP_8834 (  );
sky130_fd_sc_hd__tap_1 TAP_8835 (  );
sky130_fd_sc_hd__tap_1 TAP_8836 (  );
sky130_fd_sc_hd__tap_1 TAP_8837 (  );
sky130_fd_sc_hd__tap_1 TAP_8838 (  );
sky130_fd_sc_hd__tap_1 TAP_8839 (  );
sky130_fd_sc_hd__tap_1 TAP_884 (  );
sky130_fd_sc_hd__tap_1 TAP_8840 (  );
sky130_fd_sc_hd__tap_1 TAP_8841 (  );
sky130_fd_sc_hd__tap_1 TAP_8842 (  );
sky130_fd_sc_hd__tap_1 TAP_8843 (  );
sky130_fd_sc_hd__tap_1 TAP_8844 (  );
sky130_fd_sc_hd__tap_1 TAP_8845 (  );
sky130_fd_sc_hd__tap_1 TAP_8846 (  );
sky130_fd_sc_hd__tap_1 TAP_8847 (  );
sky130_fd_sc_hd__tap_1 TAP_8848 (  );
sky130_fd_sc_hd__tap_1 TAP_8849 (  );
sky130_fd_sc_hd__tap_1 TAP_885 (  );
sky130_fd_sc_hd__tap_1 TAP_8850 (  );
sky130_fd_sc_hd__tap_1 TAP_8851 (  );
sky130_fd_sc_hd__tap_1 TAP_8852 (  );
sky130_fd_sc_hd__tap_1 TAP_8853 (  );
sky130_fd_sc_hd__tap_1 TAP_8854 (  );
sky130_fd_sc_hd__tap_1 TAP_8855 (  );
sky130_fd_sc_hd__tap_1 TAP_8856 (  );
sky130_fd_sc_hd__tap_1 TAP_8857 (  );
sky130_fd_sc_hd__tap_1 TAP_8858 (  );
sky130_fd_sc_hd__tap_1 TAP_8859 (  );
sky130_fd_sc_hd__tap_1 TAP_886 (  );
sky130_fd_sc_hd__tap_1 TAP_8860 (  );
sky130_fd_sc_hd__tap_1 TAP_8861 (  );
sky130_fd_sc_hd__tap_1 TAP_8862 (  );
sky130_fd_sc_hd__tap_1 TAP_8863 (  );
sky130_fd_sc_hd__tap_1 TAP_8864 (  );
sky130_fd_sc_hd__tap_1 TAP_8865 (  );
sky130_fd_sc_hd__tap_1 TAP_8866 (  );
sky130_fd_sc_hd__tap_1 TAP_8867 (  );
sky130_fd_sc_hd__tap_1 TAP_8868 (  );
sky130_fd_sc_hd__tap_1 TAP_8869 (  );
sky130_fd_sc_hd__tap_1 TAP_887 (  );
sky130_fd_sc_hd__tap_1 TAP_8870 (  );
sky130_fd_sc_hd__tap_1 TAP_8871 (  );
sky130_fd_sc_hd__tap_1 TAP_8872 (  );
sky130_fd_sc_hd__tap_1 TAP_8873 (  );
sky130_fd_sc_hd__tap_1 TAP_8874 (  );
sky130_fd_sc_hd__tap_1 TAP_8875 (  );
sky130_fd_sc_hd__tap_1 TAP_8876 (  );
sky130_fd_sc_hd__tap_1 TAP_8877 (  );
sky130_fd_sc_hd__tap_1 TAP_8878 (  );
sky130_fd_sc_hd__tap_1 TAP_8879 (  );
sky130_fd_sc_hd__tap_1 TAP_888 (  );
sky130_fd_sc_hd__tap_1 TAP_8880 (  );
sky130_fd_sc_hd__tap_1 TAP_8881 (  );
sky130_fd_sc_hd__tap_1 TAP_8882 (  );
sky130_fd_sc_hd__tap_1 TAP_8883 (  );
sky130_fd_sc_hd__tap_1 TAP_8884 (  );
sky130_fd_sc_hd__tap_1 TAP_8885 (  );
sky130_fd_sc_hd__tap_1 TAP_8886 (  );
sky130_fd_sc_hd__tap_1 TAP_8887 (  );
sky130_fd_sc_hd__tap_1 TAP_8888 (  );
sky130_fd_sc_hd__tap_1 TAP_8889 (  );
sky130_fd_sc_hd__tap_1 TAP_889 (  );
sky130_fd_sc_hd__tap_1 TAP_8890 (  );
sky130_fd_sc_hd__tap_1 TAP_8891 (  );
sky130_fd_sc_hd__tap_1 TAP_8892 (  );
sky130_fd_sc_hd__tap_1 TAP_8893 (  );
sky130_fd_sc_hd__tap_1 TAP_8894 (  );
sky130_fd_sc_hd__tap_1 TAP_8895 (  );
sky130_fd_sc_hd__tap_1 TAP_8896 (  );
sky130_fd_sc_hd__tap_1 TAP_8897 (  );
sky130_fd_sc_hd__tap_1 TAP_8898 (  );
sky130_fd_sc_hd__tap_1 TAP_8899 (  );
sky130_fd_sc_hd__tap_1 TAP_890 (  );
sky130_fd_sc_hd__tap_1 TAP_8900 (  );
sky130_fd_sc_hd__tap_1 TAP_8901 (  );
sky130_fd_sc_hd__tap_1 TAP_8902 (  );
sky130_fd_sc_hd__tap_1 TAP_8903 (  );
sky130_fd_sc_hd__tap_1 TAP_8904 (  );
sky130_fd_sc_hd__tap_1 TAP_8905 (  );
sky130_fd_sc_hd__tap_1 TAP_8906 (  );
sky130_fd_sc_hd__tap_1 TAP_8907 (  );
sky130_fd_sc_hd__tap_1 TAP_8908 (  );
sky130_fd_sc_hd__tap_1 TAP_8909 (  );
sky130_fd_sc_hd__tap_1 TAP_891 (  );
sky130_fd_sc_hd__tap_1 TAP_8910 (  );
sky130_fd_sc_hd__tap_1 TAP_8911 (  );
sky130_fd_sc_hd__tap_1 TAP_8912 (  );
sky130_fd_sc_hd__tap_1 TAP_8913 (  );
sky130_fd_sc_hd__tap_1 TAP_8914 (  );
sky130_fd_sc_hd__tap_1 TAP_8915 (  );
sky130_fd_sc_hd__tap_1 TAP_8916 (  );
sky130_fd_sc_hd__tap_1 TAP_8917 (  );
sky130_fd_sc_hd__tap_1 TAP_8918 (  );
sky130_fd_sc_hd__tap_1 TAP_8919 (  );
sky130_fd_sc_hd__tap_1 TAP_892 (  );
sky130_fd_sc_hd__tap_1 TAP_8920 (  );
sky130_fd_sc_hd__tap_1 TAP_8921 (  );
sky130_fd_sc_hd__tap_1 TAP_8922 (  );
sky130_fd_sc_hd__tap_1 TAP_8923 (  );
sky130_fd_sc_hd__tap_1 TAP_8924 (  );
sky130_fd_sc_hd__tap_1 TAP_8925 (  );
sky130_fd_sc_hd__tap_1 TAP_8926 (  );
sky130_fd_sc_hd__tap_1 TAP_8927 (  );
sky130_fd_sc_hd__tap_1 TAP_8928 (  );
sky130_fd_sc_hd__tap_1 TAP_8929 (  );
sky130_fd_sc_hd__tap_1 TAP_893 (  );
sky130_fd_sc_hd__tap_1 TAP_8930 (  );
sky130_fd_sc_hd__tap_1 TAP_8931 (  );
sky130_fd_sc_hd__tap_1 TAP_8932 (  );
sky130_fd_sc_hd__tap_1 TAP_8933 (  );
sky130_fd_sc_hd__tap_1 TAP_8934 (  );
sky130_fd_sc_hd__tap_1 TAP_8935 (  );
sky130_fd_sc_hd__tap_1 TAP_8936 (  );
sky130_fd_sc_hd__tap_1 TAP_8937 (  );
sky130_fd_sc_hd__tap_1 TAP_8938 (  );
sky130_fd_sc_hd__tap_1 TAP_8939 (  );
sky130_fd_sc_hd__tap_1 TAP_894 (  );
sky130_fd_sc_hd__tap_1 TAP_8940 (  );
sky130_fd_sc_hd__tap_1 TAP_8941 (  );
sky130_fd_sc_hd__tap_1 TAP_8942 (  );
sky130_fd_sc_hd__tap_1 TAP_8943 (  );
sky130_fd_sc_hd__tap_1 TAP_8944 (  );
sky130_fd_sc_hd__tap_1 TAP_8945 (  );
sky130_fd_sc_hd__tap_1 TAP_8946 (  );
sky130_fd_sc_hd__tap_1 TAP_8947 (  );
sky130_fd_sc_hd__tap_1 TAP_8948 (  );
sky130_fd_sc_hd__tap_1 TAP_8949 (  );
sky130_fd_sc_hd__tap_1 TAP_895 (  );
sky130_fd_sc_hd__tap_1 TAP_8950 (  );
sky130_fd_sc_hd__tap_1 TAP_8951 (  );
sky130_fd_sc_hd__tap_1 TAP_8952 (  );
sky130_fd_sc_hd__tap_1 TAP_8953 (  );
sky130_fd_sc_hd__tap_1 TAP_8954 (  );
sky130_fd_sc_hd__tap_1 TAP_8955 (  );
sky130_fd_sc_hd__tap_1 TAP_8956 (  );
sky130_fd_sc_hd__tap_1 TAP_8957 (  );
sky130_fd_sc_hd__tap_1 TAP_8958 (  );
sky130_fd_sc_hd__tap_1 TAP_8959 (  );
sky130_fd_sc_hd__tap_1 TAP_896 (  );
sky130_fd_sc_hd__tap_1 TAP_8960 (  );
sky130_fd_sc_hd__tap_1 TAP_8961 (  );
sky130_fd_sc_hd__tap_1 TAP_8962 (  );
sky130_fd_sc_hd__tap_1 TAP_8963 (  );
sky130_fd_sc_hd__tap_1 TAP_8964 (  );
sky130_fd_sc_hd__tap_1 TAP_8965 (  );
sky130_fd_sc_hd__tap_1 TAP_8966 (  );
sky130_fd_sc_hd__tap_1 TAP_8967 (  );
sky130_fd_sc_hd__tap_1 TAP_8968 (  );
sky130_fd_sc_hd__tap_1 TAP_8969 (  );
sky130_fd_sc_hd__tap_1 TAP_897 (  );
sky130_fd_sc_hd__tap_1 TAP_8970 (  );
sky130_fd_sc_hd__tap_1 TAP_8971 (  );
sky130_fd_sc_hd__tap_1 TAP_8972 (  );
sky130_fd_sc_hd__tap_1 TAP_8973 (  );
sky130_fd_sc_hd__tap_1 TAP_8974 (  );
sky130_fd_sc_hd__tap_1 TAP_8975 (  );
sky130_fd_sc_hd__tap_1 TAP_8976 (  );
sky130_fd_sc_hd__tap_1 TAP_8977 (  );
sky130_fd_sc_hd__tap_1 TAP_8978 (  );
sky130_fd_sc_hd__tap_1 TAP_8979 (  );
sky130_fd_sc_hd__tap_1 TAP_898 (  );
sky130_fd_sc_hd__tap_1 TAP_8980 (  );
sky130_fd_sc_hd__tap_1 TAP_8981 (  );
sky130_fd_sc_hd__tap_1 TAP_8982 (  );
sky130_fd_sc_hd__tap_1 TAP_8983 (  );
sky130_fd_sc_hd__tap_1 TAP_8984 (  );
sky130_fd_sc_hd__tap_1 TAP_8985 (  );
sky130_fd_sc_hd__tap_1 TAP_8986 (  );
sky130_fd_sc_hd__tap_1 TAP_8987 (  );
sky130_fd_sc_hd__tap_1 TAP_8988 (  );
sky130_fd_sc_hd__tap_1 TAP_8989 (  );
sky130_fd_sc_hd__tap_1 TAP_899 (  );
sky130_fd_sc_hd__tap_1 TAP_8990 (  );
sky130_fd_sc_hd__tap_1 TAP_8991 (  );
sky130_fd_sc_hd__tap_1 TAP_8992 (  );
sky130_fd_sc_hd__tap_1 TAP_8993 (  );
sky130_fd_sc_hd__tap_1 TAP_8994 (  );
sky130_fd_sc_hd__tap_1 TAP_8995 (  );
sky130_fd_sc_hd__tap_1 TAP_8996 (  );
sky130_fd_sc_hd__tap_1 TAP_8997 (  );
sky130_fd_sc_hd__tap_1 TAP_8998 (  );
sky130_fd_sc_hd__tap_1 TAP_8999 (  );
sky130_fd_sc_hd__tap_1 TAP_900 (  );
sky130_fd_sc_hd__tap_1 TAP_9000 (  );
sky130_fd_sc_hd__tap_1 TAP_9001 (  );
sky130_fd_sc_hd__tap_1 TAP_9002 (  );
sky130_fd_sc_hd__tap_1 TAP_9003 (  );
sky130_fd_sc_hd__tap_1 TAP_9004 (  );
sky130_fd_sc_hd__tap_1 TAP_9005 (  );
sky130_fd_sc_hd__tap_1 TAP_9006 (  );
sky130_fd_sc_hd__tap_1 TAP_9007 (  );
sky130_fd_sc_hd__tap_1 TAP_9008 (  );
sky130_fd_sc_hd__tap_1 TAP_9009 (  );
sky130_fd_sc_hd__tap_1 TAP_901 (  );
sky130_fd_sc_hd__tap_1 TAP_9010 (  );
sky130_fd_sc_hd__tap_1 TAP_9011 (  );
sky130_fd_sc_hd__tap_1 TAP_9012 (  );
sky130_fd_sc_hd__tap_1 TAP_9013 (  );
sky130_fd_sc_hd__tap_1 TAP_9014 (  );
sky130_fd_sc_hd__tap_1 TAP_9015 (  );
sky130_fd_sc_hd__tap_1 TAP_9016 (  );
sky130_fd_sc_hd__tap_1 TAP_9017 (  );
sky130_fd_sc_hd__tap_1 TAP_9018 (  );
sky130_fd_sc_hd__tap_1 TAP_9019 (  );
sky130_fd_sc_hd__tap_1 TAP_902 (  );
sky130_fd_sc_hd__tap_1 TAP_9020 (  );
sky130_fd_sc_hd__tap_1 TAP_9021 (  );
sky130_fd_sc_hd__tap_1 TAP_9022 (  );
sky130_fd_sc_hd__tap_1 TAP_9023 (  );
sky130_fd_sc_hd__tap_1 TAP_9024 (  );
sky130_fd_sc_hd__tap_1 TAP_9025 (  );
sky130_fd_sc_hd__tap_1 TAP_9026 (  );
sky130_fd_sc_hd__tap_1 TAP_9027 (  );
sky130_fd_sc_hd__tap_1 TAP_9028 (  );
sky130_fd_sc_hd__tap_1 TAP_9029 (  );
sky130_fd_sc_hd__tap_1 TAP_903 (  );
sky130_fd_sc_hd__tap_1 TAP_9030 (  );
sky130_fd_sc_hd__tap_1 TAP_9031 (  );
sky130_fd_sc_hd__tap_1 TAP_9032 (  );
sky130_fd_sc_hd__tap_1 TAP_9033 (  );
sky130_fd_sc_hd__tap_1 TAP_9034 (  );
sky130_fd_sc_hd__tap_1 TAP_9035 (  );
sky130_fd_sc_hd__tap_1 TAP_9036 (  );
sky130_fd_sc_hd__tap_1 TAP_9037 (  );
sky130_fd_sc_hd__tap_1 TAP_9038 (  );
sky130_fd_sc_hd__tap_1 TAP_9039 (  );
sky130_fd_sc_hd__tap_1 TAP_904 (  );
sky130_fd_sc_hd__tap_1 TAP_9040 (  );
sky130_fd_sc_hd__tap_1 TAP_9041 (  );
sky130_fd_sc_hd__tap_1 TAP_9042 (  );
sky130_fd_sc_hd__tap_1 TAP_9043 (  );
sky130_fd_sc_hd__tap_1 TAP_9044 (  );
sky130_fd_sc_hd__tap_1 TAP_9045 (  );
sky130_fd_sc_hd__tap_1 TAP_9046 (  );
sky130_fd_sc_hd__tap_1 TAP_9047 (  );
sky130_fd_sc_hd__tap_1 TAP_9048 (  );
sky130_fd_sc_hd__tap_1 TAP_9049 (  );
sky130_fd_sc_hd__tap_1 TAP_905 (  );
sky130_fd_sc_hd__tap_1 TAP_9050 (  );
sky130_fd_sc_hd__tap_1 TAP_9051 (  );
sky130_fd_sc_hd__tap_1 TAP_9052 (  );
sky130_fd_sc_hd__tap_1 TAP_9053 (  );
sky130_fd_sc_hd__tap_1 TAP_9054 (  );
sky130_fd_sc_hd__tap_1 TAP_9055 (  );
sky130_fd_sc_hd__tap_1 TAP_9056 (  );
sky130_fd_sc_hd__tap_1 TAP_9057 (  );
sky130_fd_sc_hd__tap_1 TAP_9058 (  );
sky130_fd_sc_hd__tap_1 TAP_9059 (  );
sky130_fd_sc_hd__tap_1 TAP_906 (  );
sky130_fd_sc_hd__tap_1 TAP_9060 (  );
sky130_fd_sc_hd__tap_1 TAP_9061 (  );
sky130_fd_sc_hd__tap_1 TAP_9062 (  );
sky130_fd_sc_hd__tap_1 TAP_9063 (  );
sky130_fd_sc_hd__tap_1 TAP_9064 (  );
sky130_fd_sc_hd__tap_1 TAP_9065 (  );
sky130_fd_sc_hd__tap_1 TAP_9066 (  );
sky130_fd_sc_hd__tap_1 TAP_9067 (  );
sky130_fd_sc_hd__tap_1 TAP_9068 (  );
sky130_fd_sc_hd__tap_1 TAP_9069 (  );
sky130_fd_sc_hd__tap_1 TAP_907 (  );
sky130_fd_sc_hd__tap_1 TAP_9070 (  );
sky130_fd_sc_hd__tap_1 TAP_9071 (  );
sky130_fd_sc_hd__tap_1 TAP_9072 (  );
sky130_fd_sc_hd__tap_1 TAP_9073 (  );
sky130_fd_sc_hd__tap_1 TAP_9074 (  );
sky130_fd_sc_hd__tap_1 TAP_9075 (  );
sky130_fd_sc_hd__tap_1 TAP_9076 (  );
sky130_fd_sc_hd__tap_1 TAP_9077 (  );
sky130_fd_sc_hd__tap_1 TAP_9078 (  );
sky130_fd_sc_hd__tap_1 TAP_9079 (  );
sky130_fd_sc_hd__tap_1 TAP_908 (  );
sky130_fd_sc_hd__tap_1 TAP_9080 (  );
sky130_fd_sc_hd__tap_1 TAP_9081 (  );
sky130_fd_sc_hd__tap_1 TAP_9082 (  );
sky130_fd_sc_hd__tap_1 TAP_9083 (  );
sky130_fd_sc_hd__tap_1 TAP_9084 (  );
sky130_fd_sc_hd__tap_1 TAP_9085 (  );
sky130_fd_sc_hd__tap_1 TAP_9086 (  );
sky130_fd_sc_hd__tap_1 TAP_9087 (  );
sky130_fd_sc_hd__tap_1 TAP_9088 (  );
sky130_fd_sc_hd__tap_1 TAP_9089 (  );
sky130_fd_sc_hd__tap_1 TAP_909 (  );
sky130_fd_sc_hd__tap_1 TAP_9090 (  );
sky130_fd_sc_hd__tap_1 TAP_9091 (  );
sky130_fd_sc_hd__tap_1 TAP_9092 (  );
sky130_fd_sc_hd__tap_1 TAP_9093 (  );
sky130_fd_sc_hd__tap_1 TAP_9094 (  );
sky130_fd_sc_hd__tap_1 TAP_9095 (  );
sky130_fd_sc_hd__tap_1 TAP_9096 (  );
sky130_fd_sc_hd__tap_1 TAP_9097 (  );
sky130_fd_sc_hd__tap_1 TAP_9098 (  );
sky130_fd_sc_hd__tap_1 TAP_9099 (  );
sky130_fd_sc_hd__tap_1 TAP_910 (  );
sky130_fd_sc_hd__tap_1 TAP_9100 (  );
sky130_fd_sc_hd__tap_1 TAP_9101 (  );
sky130_fd_sc_hd__tap_1 TAP_9102 (  );
sky130_fd_sc_hd__tap_1 TAP_9103 (  );
sky130_fd_sc_hd__tap_1 TAP_9104 (  );
sky130_fd_sc_hd__tap_1 TAP_9105 (  );
sky130_fd_sc_hd__tap_1 TAP_9106 (  );
sky130_fd_sc_hd__tap_1 TAP_9107 (  );
sky130_fd_sc_hd__tap_1 TAP_9108 (  );
sky130_fd_sc_hd__tap_1 TAP_9109 (  );
sky130_fd_sc_hd__tap_1 TAP_911 (  );
sky130_fd_sc_hd__tap_1 TAP_9110 (  );
sky130_fd_sc_hd__tap_1 TAP_9111 (  );
sky130_fd_sc_hd__tap_1 TAP_9112 (  );
sky130_fd_sc_hd__tap_1 TAP_9113 (  );
sky130_fd_sc_hd__tap_1 TAP_9114 (  );
sky130_fd_sc_hd__tap_1 TAP_9115 (  );
sky130_fd_sc_hd__tap_1 TAP_9116 (  );
sky130_fd_sc_hd__tap_1 TAP_9117 (  );
sky130_fd_sc_hd__tap_1 TAP_9118 (  );
sky130_fd_sc_hd__tap_1 TAP_9119 (  );
sky130_fd_sc_hd__tap_1 TAP_912 (  );
sky130_fd_sc_hd__tap_1 TAP_9120 (  );
sky130_fd_sc_hd__tap_1 TAP_9121 (  );
sky130_fd_sc_hd__tap_1 TAP_9122 (  );
sky130_fd_sc_hd__tap_1 TAP_9123 (  );
sky130_fd_sc_hd__tap_1 TAP_9124 (  );
sky130_fd_sc_hd__tap_1 TAP_9125 (  );
sky130_fd_sc_hd__tap_1 TAP_9126 (  );
sky130_fd_sc_hd__tap_1 TAP_9127 (  );
sky130_fd_sc_hd__tap_1 TAP_9128 (  );
sky130_fd_sc_hd__tap_1 TAP_9129 (  );
sky130_fd_sc_hd__tap_1 TAP_913 (  );
sky130_fd_sc_hd__tap_1 TAP_9130 (  );
sky130_fd_sc_hd__tap_1 TAP_9131 (  );
sky130_fd_sc_hd__tap_1 TAP_9132 (  );
sky130_fd_sc_hd__tap_1 TAP_9133 (  );
sky130_fd_sc_hd__tap_1 TAP_9134 (  );
sky130_fd_sc_hd__tap_1 TAP_9135 (  );
sky130_fd_sc_hd__tap_1 TAP_9136 (  );
sky130_fd_sc_hd__tap_1 TAP_9137 (  );
sky130_fd_sc_hd__tap_1 TAP_9138 (  );
sky130_fd_sc_hd__tap_1 TAP_9139 (  );
sky130_fd_sc_hd__tap_1 TAP_914 (  );
sky130_fd_sc_hd__tap_1 TAP_9140 (  );
sky130_fd_sc_hd__tap_1 TAP_9141 (  );
sky130_fd_sc_hd__tap_1 TAP_9142 (  );
sky130_fd_sc_hd__tap_1 TAP_9143 (  );
sky130_fd_sc_hd__tap_1 TAP_9144 (  );
sky130_fd_sc_hd__tap_1 TAP_9145 (  );
sky130_fd_sc_hd__tap_1 TAP_9146 (  );
sky130_fd_sc_hd__tap_1 TAP_9147 (  );
sky130_fd_sc_hd__tap_1 TAP_9148 (  );
sky130_fd_sc_hd__tap_1 TAP_9149 (  );
sky130_fd_sc_hd__tap_1 TAP_915 (  );
sky130_fd_sc_hd__tap_1 TAP_9150 (  );
sky130_fd_sc_hd__tap_1 TAP_9151 (  );
sky130_fd_sc_hd__tap_1 TAP_9152 (  );
sky130_fd_sc_hd__tap_1 TAP_9153 (  );
sky130_fd_sc_hd__tap_1 TAP_9154 (  );
sky130_fd_sc_hd__tap_1 TAP_9155 (  );
sky130_fd_sc_hd__tap_1 TAP_9156 (  );
sky130_fd_sc_hd__tap_1 TAP_9157 (  );
sky130_fd_sc_hd__tap_1 TAP_9158 (  );
sky130_fd_sc_hd__tap_1 TAP_9159 (  );
sky130_fd_sc_hd__tap_1 TAP_916 (  );
sky130_fd_sc_hd__tap_1 TAP_9160 (  );
sky130_fd_sc_hd__tap_1 TAP_9161 (  );
sky130_fd_sc_hd__tap_1 TAP_9162 (  );
sky130_fd_sc_hd__tap_1 TAP_9163 (  );
sky130_fd_sc_hd__tap_1 TAP_9164 (  );
sky130_fd_sc_hd__tap_1 TAP_9165 (  );
sky130_fd_sc_hd__tap_1 TAP_9166 (  );
sky130_fd_sc_hd__tap_1 TAP_9167 (  );
sky130_fd_sc_hd__tap_1 TAP_9168 (  );
sky130_fd_sc_hd__tap_1 TAP_9169 (  );
sky130_fd_sc_hd__tap_1 TAP_917 (  );
sky130_fd_sc_hd__tap_1 TAP_9170 (  );
sky130_fd_sc_hd__tap_1 TAP_9171 (  );
sky130_fd_sc_hd__tap_1 TAP_9172 (  );
sky130_fd_sc_hd__tap_1 TAP_9173 (  );
sky130_fd_sc_hd__tap_1 TAP_9174 (  );
sky130_fd_sc_hd__tap_1 TAP_9175 (  );
sky130_fd_sc_hd__tap_1 TAP_9176 (  );
sky130_fd_sc_hd__tap_1 TAP_9177 (  );
sky130_fd_sc_hd__tap_1 TAP_9178 (  );
sky130_fd_sc_hd__tap_1 TAP_9179 (  );
sky130_fd_sc_hd__tap_1 TAP_918 (  );
sky130_fd_sc_hd__tap_1 TAP_9180 (  );
sky130_fd_sc_hd__tap_1 TAP_9181 (  );
sky130_fd_sc_hd__tap_1 TAP_9182 (  );
sky130_fd_sc_hd__tap_1 TAP_9183 (  );
sky130_fd_sc_hd__tap_1 TAP_9184 (  );
sky130_fd_sc_hd__tap_1 TAP_9185 (  );
sky130_fd_sc_hd__tap_1 TAP_9186 (  );
sky130_fd_sc_hd__tap_1 TAP_9187 (  );
sky130_fd_sc_hd__tap_1 TAP_9188 (  );
sky130_fd_sc_hd__tap_1 TAP_9189 (  );
sky130_fd_sc_hd__tap_1 TAP_919 (  );
sky130_fd_sc_hd__tap_1 TAP_9190 (  );
sky130_fd_sc_hd__tap_1 TAP_9191 (  );
sky130_fd_sc_hd__tap_1 TAP_9192 (  );
sky130_fd_sc_hd__tap_1 TAP_9193 (  );
sky130_fd_sc_hd__tap_1 TAP_9194 (  );
sky130_fd_sc_hd__tap_1 TAP_9195 (  );
sky130_fd_sc_hd__tap_1 TAP_9196 (  );
sky130_fd_sc_hd__tap_1 TAP_9197 (  );
sky130_fd_sc_hd__tap_1 TAP_9198 (  );
sky130_fd_sc_hd__tap_1 TAP_9199 (  );
sky130_fd_sc_hd__tap_1 TAP_920 (  );
sky130_fd_sc_hd__tap_1 TAP_9200 (  );
sky130_fd_sc_hd__tap_1 TAP_9201 (  );
sky130_fd_sc_hd__tap_1 TAP_9202 (  );
sky130_fd_sc_hd__tap_1 TAP_9203 (  );
sky130_fd_sc_hd__tap_1 TAP_9204 (  );
sky130_fd_sc_hd__tap_1 TAP_9205 (  );
sky130_fd_sc_hd__tap_1 TAP_9206 (  );
sky130_fd_sc_hd__tap_1 TAP_9207 (  );
sky130_fd_sc_hd__tap_1 TAP_9208 (  );
sky130_fd_sc_hd__tap_1 TAP_9209 (  );
sky130_fd_sc_hd__tap_1 TAP_921 (  );
sky130_fd_sc_hd__tap_1 TAP_9210 (  );
sky130_fd_sc_hd__tap_1 TAP_9211 (  );
sky130_fd_sc_hd__tap_1 TAP_9212 (  );
sky130_fd_sc_hd__tap_1 TAP_9213 (  );
sky130_fd_sc_hd__tap_1 TAP_9214 (  );
sky130_fd_sc_hd__tap_1 TAP_9215 (  );
sky130_fd_sc_hd__tap_1 TAP_9216 (  );
sky130_fd_sc_hd__tap_1 TAP_9217 (  );
sky130_fd_sc_hd__tap_1 TAP_9218 (  );
sky130_fd_sc_hd__tap_1 TAP_9219 (  );
sky130_fd_sc_hd__tap_1 TAP_922 (  );
sky130_fd_sc_hd__tap_1 TAP_9220 (  );
sky130_fd_sc_hd__tap_1 TAP_9221 (  );
sky130_fd_sc_hd__tap_1 TAP_9222 (  );
sky130_fd_sc_hd__tap_1 TAP_9223 (  );
sky130_fd_sc_hd__tap_1 TAP_9224 (  );
sky130_fd_sc_hd__tap_1 TAP_9225 (  );
sky130_fd_sc_hd__tap_1 TAP_9226 (  );
sky130_fd_sc_hd__tap_1 TAP_9227 (  );
sky130_fd_sc_hd__tap_1 TAP_9228 (  );
sky130_fd_sc_hd__tap_1 TAP_9229 (  );
sky130_fd_sc_hd__tap_1 TAP_923 (  );
sky130_fd_sc_hd__tap_1 TAP_9230 (  );
sky130_fd_sc_hd__tap_1 TAP_9231 (  );
sky130_fd_sc_hd__tap_1 TAP_9232 (  );
sky130_fd_sc_hd__tap_1 TAP_9233 (  );
sky130_fd_sc_hd__tap_1 TAP_9234 (  );
sky130_fd_sc_hd__tap_1 TAP_9235 (  );
sky130_fd_sc_hd__tap_1 TAP_9236 (  );
sky130_fd_sc_hd__tap_1 TAP_9237 (  );
sky130_fd_sc_hd__tap_1 TAP_9238 (  );
sky130_fd_sc_hd__tap_1 TAP_9239 (  );
sky130_fd_sc_hd__tap_1 TAP_924 (  );
sky130_fd_sc_hd__tap_1 TAP_9240 (  );
sky130_fd_sc_hd__tap_1 TAP_9241 (  );
sky130_fd_sc_hd__tap_1 TAP_9242 (  );
sky130_fd_sc_hd__tap_1 TAP_9243 (  );
sky130_fd_sc_hd__tap_1 TAP_9244 (  );
sky130_fd_sc_hd__tap_1 TAP_9245 (  );
sky130_fd_sc_hd__tap_1 TAP_9246 (  );
sky130_fd_sc_hd__tap_1 TAP_9247 (  );
sky130_fd_sc_hd__tap_1 TAP_9248 (  );
sky130_fd_sc_hd__tap_1 TAP_9249 (  );
sky130_fd_sc_hd__tap_1 TAP_925 (  );
sky130_fd_sc_hd__tap_1 TAP_9250 (  );
sky130_fd_sc_hd__tap_1 TAP_9251 (  );
sky130_fd_sc_hd__tap_1 TAP_9252 (  );
sky130_fd_sc_hd__tap_1 TAP_9253 (  );
sky130_fd_sc_hd__tap_1 TAP_9254 (  );
sky130_fd_sc_hd__tap_1 TAP_9255 (  );
sky130_fd_sc_hd__tap_1 TAP_9256 (  );
sky130_fd_sc_hd__tap_1 TAP_9257 (  );
sky130_fd_sc_hd__tap_1 TAP_9258 (  );
sky130_fd_sc_hd__tap_1 TAP_9259 (  );
sky130_fd_sc_hd__tap_1 TAP_926 (  );
sky130_fd_sc_hd__tap_1 TAP_9260 (  );
sky130_fd_sc_hd__tap_1 TAP_9261 (  );
sky130_fd_sc_hd__tap_1 TAP_9262 (  );
sky130_fd_sc_hd__tap_1 TAP_9263 (  );
sky130_fd_sc_hd__tap_1 TAP_9264 (  );
sky130_fd_sc_hd__tap_1 TAP_9265 (  );
sky130_fd_sc_hd__tap_1 TAP_9266 (  );
sky130_fd_sc_hd__tap_1 TAP_9267 (  );
sky130_fd_sc_hd__tap_1 TAP_9268 (  );
sky130_fd_sc_hd__tap_1 TAP_9269 (  );
sky130_fd_sc_hd__tap_1 TAP_927 (  );
sky130_fd_sc_hd__tap_1 TAP_9270 (  );
sky130_fd_sc_hd__tap_1 TAP_9271 (  );
sky130_fd_sc_hd__tap_1 TAP_9272 (  );
sky130_fd_sc_hd__tap_1 TAP_9273 (  );
sky130_fd_sc_hd__tap_1 TAP_9274 (  );
sky130_fd_sc_hd__tap_1 TAP_9275 (  );
sky130_fd_sc_hd__tap_1 TAP_9276 (  );
sky130_fd_sc_hd__tap_1 TAP_9277 (  );
sky130_fd_sc_hd__tap_1 TAP_9278 (  );
sky130_fd_sc_hd__tap_1 TAP_9279 (  );
sky130_fd_sc_hd__tap_1 TAP_928 (  );
sky130_fd_sc_hd__tap_1 TAP_9280 (  );
sky130_fd_sc_hd__tap_1 TAP_9281 (  );
sky130_fd_sc_hd__tap_1 TAP_9282 (  );
sky130_fd_sc_hd__tap_1 TAP_9283 (  );
sky130_fd_sc_hd__tap_1 TAP_9284 (  );
sky130_fd_sc_hd__tap_1 TAP_9285 (  );
sky130_fd_sc_hd__tap_1 TAP_9286 (  );
sky130_fd_sc_hd__tap_1 TAP_9287 (  );
sky130_fd_sc_hd__tap_1 TAP_9288 (  );
sky130_fd_sc_hd__tap_1 TAP_9289 (  );
sky130_fd_sc_hd__tap_1 TAP_929 (  );
sky130_fd_sc_hd__tap_1 TAP_9290 (  );
sky130_fd_sc_hd__tap_1 TAP_9291 (  );
sky130_fd_sc_hd__tap_1 TAP_9292 (  );
sky130_fd_sc_hd__tap_1 TAP_9293 (  );
sky130_fd_sc_hd__tap_1 TAP_9294 (  );
sky130_fd_sc_hd__tap_1 TAP_9295 (  );
sky130_fd_sc_hd__tap_1 TAP_9296 (  );
sky130_fd_sc_hd__tap_1 TAP_9297 (  );
sky130_fd_sc_hd__tap_1 TAP_9298 (  );
sky130_fd_sc_hd__tap_1 TAP_9299 (  );
sky130_fd_sc_hd__tap_1 TAP_930 (  );
sky130_fd_sc_hd__tap_1 TAP_9300 (  );
sky130_fd_sc_hd__tap_1 TAP_9301 (  );
sky130_fd_sc_hd__tap_1 TAP_9302 (  );
sky130_fd_sc_hd__tap_1 TAP_9303 (  );
sky130_fd_sc_hd__tap_1 TAP_9304 (  );
sky130_fd_sc_hd__tap_1 TAP_9305 (  );
sky130_fd_sc_hd__tap_1 TAP_9306 (  );
sky130_fd_sc_hd__tap_1 TAP_9307 (  );
sky130_fd_sc_hd__tap_1 TAP_9308 (  );
sky130_fd_sc_hd__tap_1 TAP_9309 (  );
sky130_fd_sc_hd__tap_1 TAP_931 (  );
sky130_fd_sc_hd__tap_1 TAP_9310 (  );
sky130_fd_sc_hd__tap_1 TAP_9311 (  );
sky130_fd_sc_hd__tap_1 TAP_9312 (  );
sky130_fd_sc_hd__tap_1 TAP_9313 (  );
sky130_fd_sc_hd__tap_1 TAP_9314 (  );
sky130_fd_sc_hd__tap_1 TAP_9315 (  );
sky130_fd_sc_hd__tap_1 TAP_9316 (  );
sky130_fd_sc_hd__tap_1 TAP_9317 (  );
sky130_fd_sc_hd__tap_1 TAP_9318 (  );
sky130_fd_sc_hd__tap_1 TAP_9319 (  );
sky130_fd_sc_hd__tap_1 TAP_932 (  );
sky130_fd_sc_hd__tap_1 TAP_9320 (  );
sky130_fd_sc_hd__tap_1 TAP_9321 (  );
sky130_fd_sc_hd__tap_1 TAP_9322 (  );
sky130_fd_sc_hd__tap_1 TAP_9323 (  );
sky130_fd_sc_hd__tap_1 TAP_9324 (  );
sky130_fd_sc_hd__tap_1 TAP_9325 (  );
sky130_fd_sc_hd__tap_1 TAP_9326 (  );
sky130_fd_sc_hd__tap_1 TAP_9327 (  );
sky130_fd_sc_hd__tap_1 TAP_9328 (  );
sky130_fd_sc_hd__tap_1 TAP_9329 (  );
sky130_fd_sc_hd__tap_1 TAP_933 (  );
sky130_fd_sc_hd__tap_1 TAP_9330 (  );
sky130_fd_sc_hd__tap_1 TAP_9331 (  );
sky130_fd_sc_hd__tap_1 TAP_9332 (  );
sky130_fd_sc_hd__tap_1 TAP_9333 (  );
sky130_fd_sc_hd__tap_1 TAP_9334 (  );
sky130_fd_sc_hd__tap_1 TAP_9335 (  );
sky130_fd_sc_hd__tap_1 TAP_9336 (  );
sky130_fd_sc_hd__tap_1 TAP_9337 (  );
sky130_fd_sc_hd__tap_1 TAP_9338 (  );
sky130_fd_sc_hd__tap_1 TAP_9339 (  );
sky130_fd_sc_hd__tap_1 TAP_934 (  );
sky130_fd_sc_hd__tap_1 TAP_9340 (  );
sky130_fd_sc_hd__tap_1 TAP_9341 (  );
sky130_fd_sc_hd__tap_1 TAP_9342 (  );
sky130_fd_sc_hd__tap_1 TAP_9343 (  );
sky130_fd_sc_hd__tap_1 TAP_9344 (  );
sky130_fd_sc_hd__tap_1 TAP_9345 (  );
sky130_fd_sc_hd__tap_1 TAP_9346 (  );
sky130_fd_sc_hd__tap_1 TAP_9347 (  );
sky130_fd_sc_hd__tap_1 TAP_9348 (  );
sky130_fd_sc_hd__tap_1 TAP_9349 (  );
sky130_fd_sc_hd__tap_1 TAP_935 (  );
sky130_fd_sc_hd__tap_1 TAP_9350 (  );
sky130_fd_sc_hd__tap_1 TAP_9351 (  );
sky130_fd_sc_hd__tap_1 TAP_9352 (  );
sky130_fd_sc_hd__tap_1 TAP_9353 (  );
sky130_fd_sc_hd__tap_1 TAP_9354 (  );
sky130_fd_sc_hd__tap_1 TAP_9355 (  );
sky130_fd_sc_hd__tap_1 TAP_9356 (  );
sky130_fd_sc_hd__tap_1 TAP_9357 (  );
sky130_fd_sc_hd__tap_1 TAP_9358 (  );
sky130_fd_sc_hd__tap_1 TAP_9359 (  );
sky130_fd_sc_hd__tap_1 TAP_936 (  );
sky130_fd_sc_hd__tap_1 TAP_9360 (  );
sky130_fd_sc_hd__tap_1 TAP_9361 (  );
sky130_fd_sc_hd__tap_1 TAP_9362 (  );
sky130_fd_sc_hd__tap_1 TAP_9363 (  );
sky130_fd_sc_hd__tap_1 TAP_9364 (  );
sky130_fd_sc_hd__tap_1 TAP_9365 (  );
sky130_fd_sc_hd__tap_1 TAP_9366 (  );
sky130_fd_sc_hd__tap_1 TAP_9367 (  );
sky130_fd_sc_hd__tap_1 TAP_9368 (  );
sky130_fd_sc_hd__tap_1 TAP_9369 (  );
sky130_fd_sc_hd__tap_1 TAP_937 (  );
sky130_fd_sc_hd__tap_1 TAP_9370 (  );
sky130_fd_sc_hd__tap_1 TAP_9371 (  );
sky130_fd_sc_hd__tap_1 TAP_9372 (  );
sky130_fd_sc_hd__tap_1 TAP_9373 (  );
sky130_fd_sc_hd__tap_1 TAP_9374 (  );
sky130_fd_sc_hd__tap_1 TAP_9375 (  );
sky130_fd_sc_hd__tap_1 TAP_9376 (  );
sky130_fd_sc_hd__tap_1 TAP_9377 (  );
sky130_fd_sc_hd__tap_1 TAP_9378 (  );
sky130_fd_sc_hd__tap_1 TAP_9379 (  );
sky130_fd_sc_hd__tap_1 TAP_938 (  );
sky130_fd_sc_hd__tap_1 TAP_9380 (  );
sky130_fd_sc_hd__tap_1 TAP_9381 (  );
sky130_fd_sc_hd__tap_1 TAP_9382 (  );
sky130_fd_sc_hd__tap_1 TAP_9383 (  );
sky130_fd_sc_hd__tap_1 TAP_9384 (  );
sky130_fd_sc_hd__tap_1 TAP_9385 (  );
sky130_fd_sc_hd__tap_1 TAP_9386 (  );
sky130_fd_sc_hd__tap_1 TAP_9387 (  );
sky130_fd_sc_hd__tap_1 TAP_9388 (  );
sky130_fd_sc_hd__tap_1 TAP_9389 (  );
sky130_fd_sc_hd__tap_1 TAP_939 (  );
sky130_fd_sc_hd__tap_1 TAP_9390 (  );
sky130_fd_sc_hd__tap_1 TAP_9391 (  );
sky130_fd_sc_hd__tap_1 TAP_9392 (  );
sky130_fd_sc_hd__tap_1 TAP_9393 (  );
sky130_fd_sc_hd__tap_1 TAP_9394 (  );
sky130_fd_sc_hd__tap_1 TAP_9395 (  );
sky130_fd_sc_hd__tap_1 TAP_9396 (  );
sky130_fd_sc_hd__tap_1 TAP_9397 (  );
sky130_fd_sc_hd__tap_1 TAP_9398 (  );
sky130_fd_sc_hd__tap_1 TAP_9399 (  );
sky130_fd_sc_hd__tap_1 TAP_940 (  );
sky130_fd_sc_hd__tap_1 TAP_9400 (  );
sky130_fd_sc_hd__tap_1 TAP_9401 (  );
sky130_fd_sc_hd__tap_1 TAP_9402 (  );
sky130_fd_sc_hd__tap_1 TAP_9403 (  );
sky130_fd_sc_hd__tap_1 TAP_9404 (  );
sky130_fd_sc_hd__tap_1 TAP_9405 (  );
sky130_fd_sc_hd__tap_1 TAP_9406 (  );
sky130_fd_sc_hd__tap_1 TAP_9407 (  );
sky130_fd_sc_hd__tap_1 TAP_9408 (  );
sky130_fd_sc_hd__tap_1 TAP_9409 (  );
sky130_fd_sc_hd__tap_1 TAP_941 (  );
sky130_fd_sc_hd__tap_1 TAP_9410 (  );
sky130_fd_sc_hd__tap_1 TAP_9411 (  );
sky130_fd_sc_hd__tap_1 TAP_9412 (  );
sky130_fd_sc_hd__tap_1 TAP_9413 (  );
sky130_fd_sc_hd__tap_1 TAP_9414 (  );
sky130_fd_sc_hd__tap_1 TAP_9415 (  );
sky130_fd_sc_hd__tap_1 TAP_9416 (  );
sky130_fd_sc_hd__tap_1 TAP_9417 (  );
sky130_fd_sc_hd__tap_1 TAP_9418 (  );
sky130_fd_sc_hd__tap_1 TAP_9419 (  );
sky130_fd_sc_hd__tap_1 TAP_942 (  );
sky130_fd_sc_hd__tap_1 TAP_9420 (  );
sky130_fd_sc_hd__tap_1 TAP_9421 (  );
sky130_fd_sc_hd__tap_1 TAP_9422 (  );
sky130_fd_sc_hd__tap_1 TAP_9423 (  );
sky130_fd_sc_hd__tap_1 TAP_9424 (  );
sky130_fd_sc_hd__tap_1 TAP_9425 (  );
sky130_fd_sc_hd__tap_1 TAP_9426 (  );
sky130_fd_sc_hd__tap_1 TAP_9427 (  );
sky130_fd_sc_hd__tap_1 TAP_9428 (  );
sky130_fd_sc_hd__tap_1 TAP_9429 (  );
sky130_fd_sc_hd__tap_1 TAP_943 (  );
sky130_fd_sc_hd__tap_1 TAP_9430 (  );
sky130_fd_sc_hd__tap_1 TAP_9431 (  );
sky130_fd_sc_hd__tap_1 TAP_9432 (  );
sky130_fd_sc_hd__tap_1 TAP_9433 (  );
sky130_fd_sc_hd__tap_1 TAP_9434 (  );
sky130_fd_sc_hd__tap_1 TAP_9435 (  );
sky130_fd_sc_hd__tap_1 TAP_9436 (  );
sky130_fd_sc_hd__tap_1 TAP_9437 (  );
sky130_fd_sc_hd__tap_1 TAP_9438 (  );
sky130_fd_sc_hd__tap_1 TAP_9439 (  );
sky130_fd_sc_hd__tap_1 TAP_944 (  );
sky130_fd_sc_hd__tap_1 TAP_9440 (  );
sky130_fd_sc_hd__tap_1 TAP_9441 (  );
sky130_fd_sc_hd__tap_1 TAP_9442 (  );
sky130_fd_sc_hd__tap_1 TAP_9443 (  );
sky130_fd_sc_hd__tap_1 TAP_9444 (  );
sky130_fd_sc_hd__tap_1 TAP_9445 (  );
sky130_fd_sc_hd__tap_1 TAP_9446 (  );
sky130_fd_sc_hd__tap_1 TAP_9447 (  );
sky130_fd_sc_hd__tap_1 TAP_9448 (  );
sky130_fd_sc_hd__tap_1 TAP_9449 (  );
sky130_fd_sc_hd__tap_1 TAP_945 (  );
sky130_fd_sc_hd__tap_1 TAP_9450 (  );
sky130_fd_sc_hd__tap_1 TAP_9451 (  );
sky130_fd_sc_hd__tap_1 TAP_9452 (  );
sky130_fd_sc_hd__tap_1 TAP_9453 (  );
sky130_fd_sc_hd__tap_1 TAP_9454 (  );
sky130_fd_sc_hd__tap_1 TAP_9455 (  );
sky130_fd_sc_hd__tap_1 TAP_9456 (  );
sky130_fd_sc_hd__tap_1 TAP_9457 (  );
sky130_fd_sc_hd__tap_1 TAP_9458 (  );
sky130_fd_sc_hd__tap_1 TAP_9459 (  );
sky130_fd_sc_hd__tap_1 TAP_946 (  );
sky130_fd_sc_hd__tap_1 TAP_9460 (  );
sky130_fd_sc_hd__tap_1 TAP_9461 (  );
sky130_fd_sc_hd__tap_1 TAP_9462 (  );
sky130_fd_sc_hd__tap_1 TAP_9463 (  );
sky130_fd_sc_hd__tap_1 TAP_9464 (  );
sky130_fd_sc_hd__tap_1 TAP_9465 (  );
sky130_fd_sc_hd__tap_1 TAP_9466 (  );
sky130_fd_sc_hd__tap_1 TAP_9467 (  );
sky130_fd_sc_hd__tap_1 TAP_9468 (  );
sky130_fd_sc_hd__tap_1 TAP_9469 (  );
sky130_fd_sc_hd__tap_1 TAP_947 (  );
sky130_fd_sc_hd__tap_1 TAP_9470 (  );
sky130_fd_sc_hd__tap_1 TAP_9471 (  );
sky130_fd_sc_hd__tap_1 TAP_9472 (  );
sky130_fd_sc_hd__tap_1 TAP_9473 (  );
sky130_fd_sc_hd__tap_1 TAP_9474 (  );
sky130_fd_sc_hd__tap_1 TAP_9475 (  );
sky130_fd_sc_hd__tap_1 TAP_9476 (  );
sky130_fd_sc_hd__tap_1 TAP_9477 (  );
sky130_fd_sc_hd__tap_1 TAP_9478 (  );
sky130_fd_sc_hd__tap_1 TAP_9479 (  );
sky130_fd_sc_hd__tap_1 TAP_948 (  );
sky130_fd_sc_hd__tap_1 TAP_9480 (  );
sky130_fd_sc_hd__tap_1 TAP_9481 (  );
sky130_fd_sc_hd__tap_1 TAP_9482 (  );
sky130_fd_sc_hd__tap_1 TAP_9483 (  );
sky130_fd_sc_hd__tap_1 TAP_9484 (  );
sky130_fd_sc_hd__tap_1 TAP_9485 (  );
sky130_fd_sc_hd__tap_1 TAP_9486 (  );
sky130_fd_sc_hd__tap_1 TAP_9487 (  );
sky130_fd_sc_hd__tap_1 TAP_9488 (  );
sky130_fd_sc_hd__tap_1 TAP_9489 (  );
sky130_fd_sc_hd__tap_1 TAP_949 (  );
sky130_fd_sc_hd__tap_1 TAP_9490 (  );
sky130_fd_sc_hd__tap_1 TAP_9491 (  );
sky130_fd_sc_hd__tap_1 TAP_9492 (  );
sky130_fd_sc_hd__tap_1 TAP_9493 (  );
sky130_fd_sc_hd__tap_1 TAP_9494 (  );
sky130_fd_sc_hd__tap_1 TAP_9495 (  );
sky130_fd_sc_hd__tap_1 TAP_9496 (  );
sky130_fd_sc_hd__tap_1 TAP_9497 (  );
sky130_fd_sc_hd__tap_1 TAP_9498 (  );
sky130_fd_sc_hd__tap_1 TAP_9499 (  );
sky130_fd_sc_hd__tap_1 TAP_950 (  );
sky130_fd_sc_hd__tap_1 TAP_9500 (  );
sky130_fd_sc_hd__tap_1 TAP_9501 (  );
sky130_fd_sc_hd__tap_1 TAP_9502 (  );
sky130_fd_sc_hd__tap_1 TAP_9503 (  );
sky130_fd_sc_hd__tap_1 TAP_9504 (  );
sky130_fd_sc_hd__tap_1 TAP_9505 (  );
sky130_fd_sc_hd__tap_1 TAP_9506 (  );
sky130_fd_sc_hd__tap_1 TAP_9507 (  );
sky130_fd_sc_hd__tap_1 TAP_9508 (  );
sky130_fd_sc_hd__tap_1 TAP_9509 (  );
sky130_fd_sc_hd__tap_1 TAP_951 (  );
sky130_fd_sc_hd__tap_1 TAP_9510 (  );
sky130_fd_sc_hd__tap_1 TAP_9511 (  );
sky130_fd_sc_hd__tap_1 TAP_9512 (  );
sky130_fd_sc_hd__tap_1 TAP_9513 (  );
sky130_fd_sc_hd__tap_1 TAP_9514 (  );
sky130_fd_sc_hd__tap_1 TAP_9515 (  );
sky130_fd_sc_hd__tap_1 TAP_9516 (  );
sky130_fd_sc_hd__tap_1 TAP_9517 (  );
sky130_fd_sc_hd__tap_1 TAP_9518 (  );
sky130_fd_sc_hd__tap_1 TAP_9519 (  );
sky130_fd_sc_hd__tap_1 TAP_952 (  );
sky130_fd_sc_hd__tap_1 TAP_9520 (  );
sky130_fd_sc_hd__tap_1 TAP_9521 (  );
sky130_fd_sc_hd__tap_1 TAP_9522 (  );
sky130_fd_sc_hd__tap_1 TAP_9523 (  );
sky130_fd_sc_hd__tap_1 TAP_9524 (  );
sky130_fd_sc_hd__tap_1 TAP_9525 (  );
sky130_fd_sc_hd__tap_1 TAP_9526 (  );
sky130_fd_sc_hd__tap_1 TAP_9527 (  );
sky130_fd_sc_hd__tap_1 TAP_9528 (  );
sky130_fd_sc_hd__tap_1 TAP_9529 (  );
sky130_fd_sc_hd__tap_1 TAP_953 (  );
sky130_fd_sc_hd__tap_1 TAP_9530 (  );
sky130_fd_sc_hd__tap_1 TAP_9531 (  );
sky130_fd_sc_hd__tap_1 TAP_9532 (  );
sky130_fd_sc_hd__tap_1 TAP_9533 (  );
sky130_fd_sc_hd__tap_1 TAP_9534 (  );
sky130_fd_sc_hd__tap_1 TAP_9535 (  );
sky130_fd_sc_hd__tap_1 TAP_9536 (  );
sky130_fd_sc_hd__tap_1 TAP_9537 (  );
sky130_fd_sc_hd__tap_1 TAP_9538 (  );
sky130_fd_sc_hd__tap_1 TAP_9539 (  );
sky130_fd_sc_hd__tap_1 TAP_954 (  );
sky130_fd_sc_hd__tap_1 TAP_9540 (  );
sky130_fd_sc_hd__tap_1 TAP_9541 (  );
sky130_fd_sc_hd__tap_1 TAP_9542 (  );
sky130_fd_sc_hd__tap_1 TAP_9543 (  );
sky130_fd_sc_hd__tap_1 TAP_9544 (  );
sky130_fd_sc_hd__tap_1 TAP_9545 (  );
sky130_fd_sc_hd__tap_1 TAP_9546 (  );
sky130_fd_sc_hd__tap_1 TAP_9547 (  );
sky130_fd_sc_hd__tap_1 TAP_9548 (  );
sky130_fd_sc_hd__tap_1 TAP_9549 (  );
sky130_fd_sc_hd__tap_1 TAP_955 (  );
sky130_fd_sc_hd__tap_1 TAP_9550 (  );
sky130_fd_sc_hd__tap_1 TAP_9551 (  );
sky130_fd_sc_hd__tap_1 TAP_9552 (  );
sky130_fd_sc_hd__tap_1 TAP_9553 (  );
sky130_fd_sc_hd__tap_1 TAP_9554 (  );
sky130_fd_sc_hd__tap_1 TAP_9555 (  );
sky130_fd_sc_hd__tap_1 TAP_9556 (  );
sky130_fd_sc_hd__tap_1 TAP_9557 (  );
sky130_fd_sc_hd__tap_1 TAP_9558 (  );
sky130_fd_sc_hd__tap_1 TAP_9559 (  );
sky130_fd_sc_hd__tap_1 TAP_956 (  );
sky130_fd_sc_hd__tap_1 TAP_9560 (  );
sky130_fd_sc_hd__tap_1 TAP_9561 (  );
sky130_fd_sc_hd__tap_1 TAP_9562 (  );
sky130_fd_sc_hd__tap_1 TAP_9563 (  );
sky130_fd_sc_hd__tap_1 TAP_9564 (  );
sky130_fd_sc_hd__tap_1 TAP_9565 (  );
sky130_fd_sc_hd__tap_1 TAP_9566 (  );
sky130_fd_sc_hd__tap_1 TAP_9567 (  );
sky130_fd_sc_hd__tap_1 TAP_9568 (  );
sky130_fd_sc_hd__tap_1 TAP_9569 (  );
sky130_fd_sc_hd__tap_1 TAP_957 (  );
sky130_fd_sc_hd__tap_1 TAP_9570 (  );
sky130_fd_sc_hd__tap_1 TAP_9571 (  );
sky130_fd_sc_hd__tap_1 TAP_9572 (  );
sky130_fd_sc_hd__tap_1 TAP_9573 (  );
sky130_fd_sc_hd__tap_1 TAP_9574 (  );
sky130_fd_sc_hd__tap_1 TAP_9575 (  );
sky130_fd_sc_hd__tap_1 TAP_9576 (  );
sky130_fd_sc_hd__tap_1 TAP_9577 (  );
sky130_fd_sc_hd__tap_1 TAP_9578 (  );
sky130_fd_sc_hd__tap_1 TAP_9579 (  );
sky130_fd_sc_hd__tap_1 TAP_958 (  );
sky130_fd_sc_hd__tap_1 TAP_9580 (  );
sky130_fd_sc_hd__tap_1 TAP_9581 (  );
sky130_fd_sc_hd__tap_1 TAP_9582 (  );
sky130_fd_sc_hd__tap_1 TAP_9583 (  );
sky130_fd_sc_hd__tap_1 TAP_9584 (  );
sky130_fd_sc_hd__tap_1 TAP_9585 (  );
sky130_fd_sc_hd__tap_1 TAP_9586 (  );
sky130_fd_sc_hd__tap_1 TAP_9587 (  );
sky130_fd_sc_hd__tap_1 TAP_9588 (  );
sky130_fd_sc_hd__tap_1 TAP_9589 (  );
sky130_fd_sc_hd__tap_1 TAP_959 (  );
sky130_fd_sc_hd__tap_1 TAP_9590 (  );
sky130_fd_sc_hd__tap_1 TAP_9591 (  );
sky130_fd_sc_hd__tap_1 TAP_9592 (  );
sky130_fd_sc_hd__tap_1 TAP_9593 (  );
sky130_fd_sc_hd__tap_1 TAP_9594 (  );
sky130_fd_sc_hd__tap_1 TAP_9595 (  );
sky130_fd_sc_hd__tap_1 TAP_9596 (  );
sky130_fd_sc_hd__tap_1 TAP_9597 (  );
sky130_fd_sc_hd__tap_1 TAP_9598 (  );
sky130_fd_sc_hd__tap_1 TAP_9599 (  );
sky130_fd_sc_hd__tap_1 TAP_960 (  );
sky130_fd_sc_hd__tap_1 TAP_9600 (  );
sky130_fd_sc_hd__tap_1 TAP_9601 (  );
sky130_fd_sc_hd__tap_1 TAP_9602 (  );
sky130_fd_sc_hd__tap_1 TAP_9603 (  );
sky130_fd_sc_hd__tap_1 TAP_9604 (  );
sky130_fd_sc_hd__tap_1 TAP_9605 (  );
sky130_fd_sc_hd__tap_1 TAP_9606 (  );
sky130_fd_sc_hd__tap_1 TAP_9607 (  );
sky130_fd_sc_hd__tap_1 TAP_9608 (  );
sky130_fd_sc_hd__tap_1 TAP_9609 (  );
sky130_fd_sc_hd__tap_1 TAP_961 (  );
sky130_fd_sc_hd__tap_1 TAP_9610 (  );
sky130_fd_sc_hd__tap_1 TAP_9611 (  );
sky130_fd_sc_hd__tap_1 TAP_9612 (  );
sky130_fd_sc_hd__tap_1 TAP_9613 (  );
sky130_fd_sc_hd__tap_1 TAP_9614 (  );
sky130_fd_sc_hd__tap_1 TAP_9615 (  );
sky130_fd_sc_hd__tap_1 TAP_9616 (  );
sky130_fd_sc_hd__tap_1 TAP_9617 (  );
sky130_fd_sc_hd__tap_1 TAP_9618 (  );
sky130_fd_sc_hd__tap_1 TAP_9619 (  );
sky130_fd_sc_hd__tap_1 TAP_962 (  );
sky130_fd_sc_hd__tap_1 TAP_9620 (  );
sky130_fd_sc_hd__tap_1 TAP_9621 (  );
sky130_fd_sc_hd__tap_1 TAP_9622 (  );
sky130_fd_sc_hd__tap_1 TAP_9623 (  );
sky130_fd_sc_hd__tap_1 TAP_9624 (  );
sky130_fd_sc_hd__tap_1 TAP_9625 (  );
sky130_fd_sc_hd__tap_1 TAP_9626 (  );
sky130_fd_sc_hd__tap_1 TAP_9627 (  );
sky130_fd_sc_hd__tap_1 TAP_9628 (  );
sky130_fd_sc_hd__tap_1 TAP_9629 (  );
sky130_fd_sc_hd__tap_1 TAP_963 (  );
sky130_fd_sc_hd__tap_1 TAP_9630 (  );
sky130_fd_sc_hd__tap_1 TAP_9631 (  );
sky130_fd_sc_hd__tap_1 TAP_9632 (  );
sky130_fd_sc_hd__tap_1 TAP_9633 (  );
sky130_fd_sc_hd__tap_1 TAP_9634 (  );
sky130_fd_sc_hd__tap_1 TAP_9635 (  );
sky130_fd_sc_hd__tap_1 TAP_9636 (  );
sky130_fd_sc_hd__tap_1 TAP_9637 (  );
sky130_fd_sc_hd__tap_1 TAP_9638 (  );
sky130_fd_sc_hd__tap_1 TAP_9639 (  );
sky130_fd_sc_hd__tap_1 TAP_964 (  );
sky130_fd_sc_hd__tap_1 TAP_9640 (  );
sky130_fd_sc_hd__tap_1 TAP_9641 (  );
sky130_fd_sc_hd__tap_1 TAP_9642 (  );
sky130_fd_sc_hd__tap_1 TAP_9643 (  );
sky130_fd_sc_hd__tap_1 TAP_9644 (  );
sky130_fd_sc_hd__tap_1 TAP_9645 (  );
sky130_fd_sc_hd__tap_1 TAP_9646 (  );
sky130_fd_sc_hd__tap_1 TAP_9647 (  );
sky130_fd_sc_hd__tap_1 TAP_9648 (  );
sky130_fd_sc_hd__tap_1 TAP_9649 (  );
sky130_fd_sc_hd__tap_1 TAP_965 (  );
sky130_fd_sc_hd__tap_1 TAP_9650 (  );
sky130_fd_sc_hd__tap_1 TAP_9651 (  );
sky130_fd_sc_hd__tap_1 TAP_9652 (  );
sky130_fd_sc_hd__tap_1 TAP_9653 (  );
sky130_fd_sc_hd__tap_1 TAP_9654 (  );
sky130_fd_sc_hd__tap_1 TAP_9655 (  );
sky130_fd_sc_hd__tap_1 TAP_9656 (  );
sky130_fd_sc_hd__tap_1 TAP_9657 (  );
sky130_fd_sc_hd__tap_1 TAP_9658 (  );
sky130_fd_sc_hd__tap_1 TAP_9659 (  );
sky130_fd_sc_hd__tap_1 TAP_966 (  );
sky130_fd_sc_hd__tap_1 TAP_9660 (  );
sky130_fd_sc_hd__tap_1 TAP_9661 (  );
sky130_fd_sc_hd__tap_1 TAP_9662 (  );
sky130_fd_sc_hd__tap_1 TAP_9663 (  );
sky130_fd_sc_hd__tap_1 TAP_9664 (  );
sky130_fd_sc_hd__tap_1 TAP_9665 (  );
sky130_fd_sc_hd__tap_1 TAP_9666 (  );
sky130_fd_sc_hd__tap_1 TAP_9667 (  );
sky130_fd_sc_hd__tap_1 TAP_9668 (  );
sky130_fd_sc_hd__tap_1 TAP_9669 (  );
sky130_fd_sc_hd__tap_1 TAP_967 (  );
sky130_fd_sc_hd__tap_1 TAP_9670 (  );
sky130_fd_sc_hd__tap_1 TAP_9671 (  );
sky130_fd_sc_hd__tap_1 TAP_9672 (  );
sky130_fd_sc_hd__tap_1 TAP_9673 (  );
sky130_fd_sc_hd__tap_1 TAP_9674 (  );
sky130_fd_sc_hd__tap_1 TAP_9675 (  );
sky130_fd_sc_hd__tap_1 TAP_9676 (  );
sky130_fd_sc_hd__tap_1 TAP_9677 (  );
sky130_fd_sc_hd__tap_1 TAP_9678 (  );
sky130_fd_sc_hd__tap_1 TAP_9679 (  );
sky130_fd_sc_hd__tap_1 TAP_968 (  );
sky130_fd_sc_hd__tap_1 TAP_9680 (  );
sky130_fd_sc_hd__tap_1 TAP_9681 (  );
sky130_fd_sc_hd__tap_1 TAP_9682 (  );
sky130_fd_sc_hd__tap_1 TAP_9683 (  );
sky130_fd_sc_hd__tap_1 TAP_9684 (  );
sky130_fd_sc_hd__tap_1 TAP_9685 (  );
sky130_fd_sc_hd__tap_1 TAP_9686 (  );
sky130_fd_sc_hd__tap_1 TAP_9687 (  );
sky130_fd_sc_hd__tap_1 TAP_9688 (  );
sky130_fd_sc_hd__tap_1 TAP_9689 (  );
sky130_fd_sc_hd__tap_1 TAP_969 (  );
sky130_fd_sc_hd__tap_1 TAP_9690 (  );
sky130_fd_sc_hd__tap_1 TAP_9691 (  );
sky130_fd_sc_hd__tap_1 TAP_9692 (  );
sky130_fd_sc_hd__tap_1 TAP_9693 (  );
sky130_fd_sc_hd__tap_1 TAP_9694 (  );
sky130_fd_sc_hd__tap_1 TAP_9695 (  );
sky130_fd_sc_hd__tap_1 TAP_9696 (  );
sky130_fd_sc_hd__tap_1 TAP_9697 (  );
sky130_fd_sc_hd__tap_1 TAP_9698 (  );
sky130_fd_sc_hd__tap_1 TAP_9699 (  );
sky130_fd_sc_hd__tap_1 TAP_970 (  );
sky130_fd_sc_hd__tap_1 TAP_9700 (  );
sky130_fd_sc_hd__tap_1 TAP_9701 (  );
sky130_fd_sc_hd__tap_1 TAP_9702 (  );
sky130_fd_sc_hd__tap_1 TAP_9703 (  );
sky130_fd_sc_hd__tap_1 TAP_9704 (  );
sky130_fd_sc_hd__tap_1 TAP_9705 (  );
sky130_fd_sc_hd__tap_1 TAP_9706 (  );
sky130_fd_sc_hd__tap_1 TAP_9707 (  );
sky130_fd_sc_hd__tap_1 TAP_9708 (  );
sky130_fd_sc_hd__tap_1 TAP_9709 (  );
sky130_fd_sc_hd__tap_1 TAP_971 (  );
sky130_fd_sc_hd__tap_1 TAP_9710 (  );
sky130_fd_sc_hd__tap_1 TAP_9711 (  );
sky130_fd_sc_hd__tap_1 TAP_9712 (  );
sky130_fd_sc_hd__tap_1 TAP_9713 (  );
sky130_fd_sc_hd__tap_1 TAP_9714 (  );
sky130_fd_sc_hd__tap_1 TAP_9715 (  );
sky130_fd_sc_hd__tap_1 TAP_9716 (  );
sky130_fd_sc_hd__tap_1 TAP_9717 (  );
sky130_fd_sc_hd__tap_1 TAP_9718 (  );
sky130_fd_sc_hd__tap_1 TAP_9719 (  );
sky130_fd_sc_hd__tap_1 TAP_972 (  );
sky130_fd_sc_hd__tap_1 TAP_9720 (  );
sky130_fd_sc_hd__tap_1 TAP_9721 (  );
sky130_fd_sc_hd__tap_1 TAP_9722 (  );
sky130_fd_sc_hd__tap_1 TAP_9723 (  );
sky130_fd_sc_hd__tap_1 TAP_9724 (  );
sky130_fd_sc_hd__tap_1 TAP_9725 (  );
sky130_fd_sc_hd__tap_1 TAP_9726 (  );
sky130_fd_sc_hd__tap_1 TAP_9727 (  );
sky130_fd_sc_hd__tap_1 TAP_9728 (  );
sky130_fd_sc_hd__tap_1 TAP_9729 (  );
sky130_fd_sc_hd__tap_1 TAP_973 (  );
sky130_fd_sc_hd__tap_1 TAP_9730 (  );
sky130_fd_sc_hd__tap_1 TAP_9731 (  );
sky130_fd_sc_hd__tap_1 TAP_9732 (  );
sky130_fd_sc_hd__tap_1 TAP_9733 (  );
sky130_fd_sc_hd__tap_1 TAP_9734 (  );
sky130_fd_sc_hd__tap_1 TAP_9735 (  );
sky130_fd_sc_hd__tap_1 TAP_9736 (  );
sky130_fd_sc_hd__tap_1 TAP_9737 (  );
sky130_fd_sc_hd__tap_1 TAP_9738 (  );
sky130_fd_sc_hd__tap_1 TAP_9739 (  );
sky130_fd_sc_hd__tap_1 TAP_974 (  );
sky130_fd_sc_hd__tap_1 TAP_9740 (  );
sky130_fd_sc_hd__tap_1 TAP_9741 (  );
sky130_fd_sc_hd__tap_1 TAP_9742 (  );
sky130_fd_sc_hd__tap_1 TAP_9743 (  );
sky130_fd_sc_hd__tap_1 TAP_9744 (  );
sky130_fd_sc_hd__tap_1 TAP_9745 (  );
sky130_fd_sc_hd__tap_1 TAP_9746 (  );
sky130_fd_sc_hd__tap_1 TAP_9747 (  );
sky130_fd_sc_hd__tap_1 TAP_9748 (  );
sky130_fd_sc_hd__tap_1 TAP_9749 (  );
sky130_fd_sc_hd__tap_1 TAP_975 (  );
sky130_fd_sc_hd__tap_1 TAP_9750 (  );
sky130_fd_sc_hd__tap_1 TAP_9751 (  );
sky130_fd_sc_hd__tap_1 TAP_9752 (  );
sky130_fd_sc_hd__tap_1 TAP_9753 (  );
sky130_fd_sc_hd__tap_1 TAP_9754 (  );
sky130_fd_sc_hd__tap_1 TAP_9755 (  );
sky130_fd_sc_hd__tap_1 TAP_9756 (  );
sky130_fd_sc_hd__tap_1 TAP_9757 (  );
sky130_fd_sc_hd__tap_1 TAP_9758 (  );
sky130_fd_sc_hd__tap_1 TAP_9759 (  );
sky130_fd_sc_hd__tap_1 TAP_976 (  );
sky130_fd_sc_hd__tap_1 TAP_9760 (  );
sky130_fd_sc_hd__tap_1 TAP_9761 (  );
sky130_fd_sc_hd__tap_1 TAP_9762 (  );
sky130_fd_sc_hd__tap_1 TAP_9763 (  );
sky130_fd_sc_hd__tap_1 TAP_9764 (  );
sky130_fd_sc_hd__tap_1 TAP_9765 (  );
sky130_fd_sc_hd__tap_1 TAP_9766 (  );
sky130_fd_sc_hd__tap_1 TAP_9767 (  );
sky130_fd_sc_hd__tap_1 TAP_9768 (  );
sky130_fd_sc_hd__tap_1 TAP_9769 (  );
sky130_fd_sc_hd__tap_1 TAP_977 (  );
sky130_fd_sc_hd__tap_1 TAP_9770 (  );
sky130_fd_sc_hd__tap_1 TAP_9771 (  );
sky130_fd_sc_hd__tap_1 TAP_9772 (  );
sky130_fd_sc_hd__tap_1 TAP_9773 (  );
sky130_fd_sc_hd__tap_1 TAP_9774 (  );
sky130_fd_sc_hd__tap_1 TAP_9775 (  );
sky130_fd_sc_hd__tap_1 TAP_9776 (  );
sky130_fd_sc_hd__tap_1 TAP_9777 (  );
sky130_fd_sc_hd__tap_1 TAP_9778 (  );
sky130_fd_sc_hd__tap_1 TAP_9779 (  );
sky130_fd_sc_hd__tap_1 TAP_978 (  );
sky130_fd_sc_hd__tap_1 TAP_9780 (  );
sky130_fd_sc_hd__tap_1 TAP_9781 (  );
sky130_fd_sc_hd__tap_1 TAP_9782 (  );
sky130_fd_sc_hd__tap_1 TAP_9783 (  );
sky130_fd_sc_hd__tap_1 TAP_9784 (  );
sky130_fd_sc_hd__tap_1 TAP_9785 (  );
sky130_fd_sc_hd__tap_1 TAP_9786 (  );
sky130_fd_sc_hd__tap_1 TAP_9787 (  );
sky130_fd_sc_hd__tap_1 TAP_9788 (  );
sky130_fd_sc_hd__tap_1 TAP_9789 (  );
sky130_fd_sc_hd__tap_1 TAP_979 (  );
sky130_fd_sc_hd__tap_1 TAP_9790 (  );
sky130_fd_sc_hd__tap_1 TAP_9791 (  );
sky130_fd_sc_hd__tap_1 TAP_9792 (  );
sky130_fd_sc_hd__tap_1 TAP_9793 (  );
sky130_fd_sc_hd__tap_1 TAP_9794 (  );
sky130_fd_sc_hd__tap_1 TAP_9795 (  );
sky130_fd_sc_hd__tap_1 TAP_9796 (  );
sky130_fd_sc_hd__tap_1 TAP_9797 (  );
sky130_fd_sc_hd__tap_1 TAP_9798 (  );
sky130_fd_sc_hd__tap_1 TAP_9799 (  );
sky130_fd_sc_hd__tap_1 TAP_980 (  );
sky130_fd_sc_hd__tap_1 TAP_9800 (  );
sky130_fd_sc_hd__tap_1 TAP_9801 (  );
sky130_fd_sc_hd__tap_1 TAP_9802 (  );
sky130_fd_sc_hd__tap_1 TAP_9803 (  );
sky130_fd_sc_hd__tap_1 TAP_9804 (  );
sky130_fd_sc_hd__tap_1 TAP_9805 (  );
sky130_fd_sc_hd__tap_1 TAP_9806 (  );
sky130_fd_sc_hd__tap_1 TAP_9807 (  );
sky130_fd_sc_hd__tap_1 TAP_9808 (  );
sky130_fd_sc_hd__tap_1 TAP_9809 (  );
sky130_fd_sc_hd__tap_1 TAP_981 (  );
sky130_fd_sc_hd__tap_1 TAP_9810 (  );
sky130_fd_sc_hd__tap_1 TAP_9811 (  );
sky130_fd_sc_hd__tap_1 TAP_9812 (  );
sky130_fd_sc_hd__tap_1 TAP_9813 (  );
sky130_fd_sc_hd__tap_1 TAP_9814 (  );
sky130_fd_sc_hd__tap_1 TAP_9815 (  );
sky130_fd_sc_hd__tap_1 TAP_9816 (  );
sky130_fd_sc_hd__tap_1 TAP_9817 (  );
sky130_fd_sc_hd__tap_1 TAP_9818 (  );
sky130_fd_sc_hd__tap_1 TAP_9819 (  );
sky130_fd_sc_hd__tap_1 TAP_982 (  );
sky130_fd_sc_hd__tap_1 TAP_9820 (  );
sky130_fd_sc_hd__tap_1 TAP_9821 (  );
sky130_fd_sc_hd__tap_1 TAP_9822 (  );
sky130_fd_sc_hd__tap_1 TAP_9823 (  );
sky130_fd_sc_hd__tap_1 TAP_9824 (  );
sky130_fd_sc_hd__tap_1 TAP_9825 (  );
sky130_fd_sc_hd__tap_1 TAP_9826 (  );
sky130_fd_sc_hd__tap_1 TAP_9827 (  );
sky130_fd_sc_hd__tap_1 TAP_9828 (  );
sky130_fd_sc_hd__tap_1 TAP_9829 (  );
sky130_fd_sc_hd__tap_1 TAP_983 (  );
sky130_fd_sc_hd__tap_1 TAP_9830 (  );
sky130_fd_sc_hd__tap_1 TAP_9831 (  );
sky130_fd_sc_hd__tap_1 TAP_9832 (  );
sky130_fd_sc_hd__tap_1 TAP_9833 (  );
sky130_fd_sc_hd__tap_1 TAP_9834 (  );
sky130_fd_sc_hd__tap_1 TAP_9835 (  );
sky130_fd_sc_hd__tap_1 TAP_9836 (  );
sky130_fd_sc_hd__tap_1 TAP_9837 (  );
sky130_fd_sc_hd__tap_1 TAP_9838 (  );
sky130_fd_sc_hd__tap_1 TAP_9839 (  );
sky130_fd_sc_hd__tap_1 TAP_984 (  );
sky130_fd_sc_hd__tap_1 TAP_9840 (  );
sky130_fd_sc_hd__tap_1 TAP_9841 (  );
sky130_fd_sc_hd__tap_1 TAP_9842 (  );
sky130_fd_sc_hd__tap_1 TAP_9843 (  );
sky130_fd_sc_hd__tap_1 TAP_9844 (  );
sky130_fd_sc_hd__tap_1 TAP_9845 (  );
sky130_fd_sc_hd__tap_1 TAP_9846 (  );
sky130_fd_sc_hd__tap_1 TAP_9847 (  );
sky130_fd_sc_hd__tap_1 TAP_9848 (  );
sky130_fd_sc_hd__tap_1 TAP_9849 (  );
sky130_fd_sc_hd__tap_1 TAP_985 (  );
sky130_fd_sc_hd__tap_1 TAP_9850 (  );
sky130_fd_sc_hd__tap_1 TAP_9851 (  );
sky130_fd_sc_hd__tap_1 TAP_9852 (  );
sky130_fd_sc_hd__tap_1 TAP_9853 (  );
sky130_fd_sc_hd__tap_1 TAP_9854 (  );
sky130_fd_sc_hd__tap_1 TAP_9855 (  );
sky130_fd_sc_hd__tap_1 TAP_9856 (  );
sky130_fd_sc_hd__tap_1 TAP_9857 (  );
sky130_fd_sc_hd__tap_1 TAP_9858 (  );
sky130_fd_sc_hd__tap_1 TAP_9859 (  );
sky130_fd_sc_hd__tap_1 TAP_986 (  );
sky130_fd_sc_hd__tap_1 TAP_9860 (  );
sky130_fd_sc_hd__tap_1 TAP_9861 (  );
sky130_fd_sc_hd__tap_1 TAP_9862 (  );
sky130_fd_sc_hd__tap_1 TAP_9863 (  );
sky130_fd_sc_hd__tap_1 TAP_9864 (  );
sky130_fd_sc_hd__tap_1 TAP_9865 (  );
sky130_fd_sc_hd__tap_1 TAP_9866 (  );
sky130_fd_sc_hd__tap_1 TAP_9867 (  );
sky130_fd_sc_hd__tap_1 TAP_9868 (  );
sky130_fd_sc_hd__tap_1 TAP_9869 (  );
sky130_fd_sc_hd__tap_1 TAP_987 (  );
sky130_fd_sc_hd__tap_1 TAP_9870 (  );
sky130_fd_sc_hd__tap_1 TAP_9871 (  );
sky130_fd_sc_hd__tap_1 TAP_9872 (  );
sky130_fd_sc_hd__tap_1 TAP_9873 (  );
sky130_fd_sc_hd__tap_1 TAP_9874 (  );
sky130_fd_sc_hd__tap_1 TAP_9875 (  );
sky130_fd_sc_hd__tap_1 TAP_9876 (  );
sky130_fd_sc_hd__tap_1 TAP_9877 (  );
sky130_fd_sc_hd__tap_1 TAP_9878 (  );
sky130_fd_sc_hd__tap_1 TAP_9879 (  );
sky130_fd_sc_hd__tap_1 TAP_988 (  );
sky130_fd_sc_hd__tap_1 TAP_9880 (  );
sky130_fd_sc_hd__tap_1 TAP_9881 (  );
sky130_fd_sc_hd__tap_1 TAP_9882 (  );
sky130_fd_sc_hd__tap_1 TAP_9883 (  );
sky130_fd_sc_hd__tap_1 TAP_9884 (  );
sky130_fd_sc_hd__tap_1 TAP_9885 (  );
sky130_fd_sc_hd__tap_1 TAP_9886 (  );
sky130_fd_sc_hd__tap_1 TAP_9887 (  );
sky130_fd_sc_hd__tap_1 TAP_9888 (  );
sky130_fd_sc_hd__tap_1 TAP_9889 (  );
sky130_fd_sc_hd__tap_1 TAP_989 (  );
sky130_fd_sc_hd__tap_1 TAP_9890 (  );
sky130_fd_sc_hd__tap_1 TAP_9891 (  );
sky130_fd_sc_hd__tap_1 TAP_9892 (  );
sky130_fd_sc_hd__tap_1 TAP_9893 (  );
sky130_fd_sc_hd__tap_1 TAP_9894 (  );
sky130_fd_sc_hd__tap_1 TAP_9895 (  );
sky130_fd_sc_hd__tap_1 TAP_9896 (  );
sky130_fd_sc_hd__tap_1 TAP_9897 (  );
sky130_fd_sc_hd__tap_1 TAP_9898 (  );
sky130_fd_sc_hd__tap_1 TAP_9899 (  );
sky130_fd_sc_hd__tap_1 TAP_990 (  );
sky130_fd_sc_hd__tap_1 TAP_9900 (  );
sky130_fd_sc_hd__tap_1 TAP_9901 (  );
sky130_fd_sc_hd__tap_1 TAP_9902 (  );
sky130_fd_sc_hd__tap_1 TAP_9903 (  );
sky130_fd_sc_hd__tap_1 TAP_9904 (  );
sky130_fd_sc_hd__tap_1 TAP_9905 (  );
sky130_fd_sc_hd__tap_1 TAP_9906 (  );
sky130_fd_sc_hd__tap_1 TAP_9907 (  );
sky130_fd_sc_hd__tap_1 TAP_9908 (  );
sky130_fd_sc_hd__tap_1 TAP_9909 (  );
sky130_fd_sc_hd__tap_1 TAP_991 (  );
sky130_fd_sc_hd__tap_1 TAP_9910 (  );
sky130_fd_sc_hd__tap_1 TAP_9911 (  );
sky130_fd_sc_hd__tap_1 TAP_9912 (  );
sky130_fd_sc_hd__tap_1 TAP_9913 (  );
sky130_fd_sc_hd__tap_1 TAP_9914 (  );
sky130_fd_sc_hd__tap_1 TAP_9915 (  );
sky130_fd_sc_hd__tap_1 TAP_9916 (  );
sky130_fd_sc_hd__tap_1 TAP_9917 (  );
sky130_fd_sc_hd__tap_1 TAP_9918 (  );
sky130_fd_sc_hd__tap_1 TAP_9919 (  );
sky130_fd_sc_hd__tap_1 TAP_992 (  );
sky130_fd_sc_hd__tap_1 TAP_9920 (  );
sky130_fd_sc_hd__tap_1 TAP_9921 (  );
sky130_fd_sc_hd__tap_1 TAP_9922 (  );
sky130_fd_sc_hd__tap_1 TAP_9923 (  );
sky130_fd_sc_hd__tap_1 TAP_9924 (  );
sky130_fd_sc_hd__tap_1 TAP_9925 (  );
sky130_fd_sc_hd__tap_1 TAP_9926 (  );
sky130_fd_sc_hd__tap_1 TAP_9927 (  );
sky130_fd_sc_hd__tap_1 TAP_9928 (  );
sky130_fd_sc_hd__tap_1 TAP_9929 (  );
sky130_fd_sc_hd__tap_1 TAP_993 (  );
sky130_fd_sc_hd__tap_1 TAP_9930 (  );
sky130_fd_sc_hd__tap_1 TAP_9931 (  );
sky130_fd_sc_hd__tap_1 TAP_9932 (  );
sky130_fd_sc_hd__tap_1 TAP_9933 (  );
sky130_fd_sc_hd__tap_1 TAP_9934 (  );
sky130_fd_sc_hd__tap_1 TAP_9935 (  );
sky130_fd_sc_hd__tap_1 TAP_9936 (  );
sky130_fd_sc_hd__tap_1 TAP_9937 (  );
sky130_fd_sc_hd__tap_1 TAP_9938 (  );
sky130_fd_sc_hd__tap_1 TAP_9939 (  );
sky130_fd_sc_hd__tap_1 TAP_994 (  );
sky130_fd_sc_hd__tap_1 TAP_9940 (  );
sky130_fd_sc_hd__tap_1 TAP_9941 (  );
sky130_fd_sc_hd__tap_1 TAP_9942 (  );
sky130_fd_sc_hd__tap_1 TAP_9943 (  );
sky130_fd_sc_hd__tap_1 TAP_9944 (  );
sky130_fd_sc_hd__tap_1 TAP_9945 (  );
sky130_fd_sc_hd__tap_1 TAP_9946 (  );
sky130_fd_sc_hd__tap_1 TAP_9947 (  );
sky130_fd_sc_hd__tap_1 TAP_9948 (  );
sky130_fd_sc_hd__tap_1 TAP_9949 (  );
sky130_fd_sc_hd__tap_1 TAP_995 (  );
sky130_fd_sc_hd__tap_1 TAP_9950 (  );
sky130_fd_sc_hd__tap_1 TAP_9951 (  );
sky130_fd_sc_hd__tap_1 TAP_9952 (  );
sky130_fd_sc_hd__tap_1 TAP_9953 (  );
sky130_fd_sc_hd__tap_1 TAP_9954 (  );
sky130_fd_sc_hd__tap_1 TAP_9955 (  );
sky130_fd_sc_hd__tap_1 TAP_9956 (  );
sky130_fd_sc_hd__tap_1 TAP_9957 (  );
sky130_fd_sc_hd__tap_1 TAP_9958 (  );
sky130_fd_sc_hd__tap_1 TAP_9959 (  );
sky130_fd_sc_hd__tap_1 TAP_996 (  );
sky130_fd_sc_hd__tap_1 TAP_9960 (  );
sky130_fd_sc_hd__tap_1 TAP_9961 (  );
sky130_fd_sc_hd__tap_1 TAP_9962 (  );
sky130_fd_sc_hd__tap_1 TAP_9963 (  );
sky130_fd_sc_hd__tap_1 TAP_9964 (  );
sky130_fd_sc_hd__tap_1 TAP_9965 (  );
sky130_fd_sc_hd__tap_1 TAP_9966 (  );
sky130_fd_sc_hd__tap_1 TAP_9967 (  );
sky130_fd_sc_hd__tap_1 TAP_9968 (  );
sky130_fd_sc_hd__tap_1 TAP_9969 (  );
sky130_fd_sc_hd__tap_1 TAP_997 (  );
sky130_fd_sc_hd__tap_1 TAP_9970 (  );
sky130_fd_sc_hd__tap_1 TAP_9971 (  );
sky130_fd_sc_hd__tap_1 TAP_9972 (  );
sky130_fd_sc_hd__tap_1 TAP_9973 (  );
sky130_fd_sc_hd__tap_1 TAP_9974 (  );
sky130_fd_sc_hd__tap_1 TAP_9975 (  );
sky130_fd_sc_hd__tap_1 TAP_9976 (  );
sky130_fd_sc_hd__tap_1 TAP_9977 (  );
sky130_fd_sc_hd__tap_1 TAP_9978 (  );
sky130_fd_sc_hd__tap_1 TAP_9979 (  );
sky130_fd_sc_hd__tap_1 TAP_998 (  );
sky130_fd_sc_hd__tap_1 TAP_9980 (  );
sky130_fd_sc_hd__tap_1 TAP_9981 (  );
sky130_fd_sc_hd__tap_1 TAP_9982 (  );
sky130_fd_sc_hd__tap_1 TAP_9983 (  );
sky130_fd_sc_hd__tap_1 TAP_9984 (  );
sky130_fd_sc_hd__tap_1 TAP_9985 (  );
sky130_fd_sc_hd__tap_1 TAP_9986 (  );
sky130_fd_sc_hd__tap_1 TAP_9987 (  );
sky130_fd_sc_hd__tap_1 TAP_9988 (  );
sky130_fd_sc_hd__tap_1 TAP_9989 (  );
sky130_fd_sc_hd__tap_1 TAP_999 (  );
sky130_fd_sc_hd__tap_1 TAP_9990 (  );
sky130_fd_sc_hd__tap_1 TAP_9991 (  );
sky130_fd_sc_hd__tap_1 TAP_9992 (  );
sky130_fd_sc_hd__tap_1 TAP_9993 (  );
sky130_fd_sc_hd__tap_1 TAP_9994 (  );
sky130_fd_sc_hd__tap_1 TAP_9995 (  );
sky130_fd_sc_hd__tap_1 TAP_9996 (  );
sky130_fd_sc_hd__tap_1 TAP_9997 (  );
sky130_fd_sc_hd__tap_1 TAP_9998 (  );
sky130_fd_sc_hd__tap_1 TAP_9999 (  );
sky130_fd_sc_hd__clkbuf_1 _1940_ ( .A(ld ), .X(_1278_ ) );
sky130_fd_sc_hd__buf_2 _1941_ ( .A(_1278_ ), .X(_1279_ ) );
sky130_fd_sc_hd__inv_1 _1942_ ( .A(\dcnt\[0\] ), .Y(_1280_ ) );
sky130_fd_sc_hd__nor2_1 _1943_ ( .A(\dcnt\[1\] ), .B(\dcnt\[2\] ), .Y(_1281_ ) );
sky130_fd_sc_hd__clkbuf_1 _1944_ ( .A(ld ), .X(_1282_ ) );
sky130_fd_sc_hd__inv_1 _1945_ ( .A(_1282_ ), .Y(_1283_ ) );
sky130_fd_sc_hd__nand3b_1 _1946_ ( .A_N(\dcnt\[3\] ), .B(_1281_ ), .C(_1283_ ), .Y(_1284_ ) );
sky130_fd_sc_hd__o211a_1 _1947_ ( .A1(_1279_ ), .A2(_1280_ ), .B1(rst ), .C1(_1284_ ), .X(_0261_ ) );
sky130_fd_sc_hd__or2b_1 _1948_ ( .A(\dcnt\[3\] ), .B_N(_1281_ ), .X(_1285_ ) );
sky130_fd_sc_hd__nor2_1 _1949_ ( .A(\dcnt\[0\] ), .B(\dcnt\[1\] ), .Y(_1286_ ) );
sky130_fd_sc_hd__nand2_1 _1950_ ( .A(_1285_ ), .B(_1286_ ), .Y(_1287_ ) );
sky130_fd_sc_hd__nand2_1 _1951_ ( .A(\dcnt\[0\] ), .B(\dcnt\[1\] ), .Y(_1288_ ) );
sky130_fd_sc_hd__inv_1 _1952_ ( .A(rst ), .Y(_1289_ ) );
sky130_fd_sc_hd__a31oi_1 _1953_ ( .A1(_1287_ ), .A2(_1283_ ), .A3(_1288_ ), .B1(_1289_ ), .Y(_0262_ ) );
sky130_fd_sc_hd__or2b_1 _1954_ ( .A(_1285_ ), .B_N(_1280_ ), .X(_1290_ ) );
sky130_fd_sc_hd__xor2_1 _1955_ ( .A(\dcnt\[2\] ), .B(_1286_ ), .X(_1291_ ) );
sky130_fd_sc_hd__and4_1 _1956_ ( .A(_1290_ ), .B(_1283_ ), .C(rst ), .D(_1291_ ), .X(_0263_ ) );
sky130_fd_sc_hd__o31ai_1 _1957_ ( .A1(\dcnt\[0\] ), .A2(\dcnt\[1\] ), .A3(\dcnt\[2\] ), .B1(\dcnt\[3\] ), .Y(_1292_ ) );
sky130_fd_sc_hd__a21oi_1 _1958_ ( .A1(_1292_ ), .A2(_1283_ ), .B1(_1289_ ), .Y(_0264_ ) );
sky130_fd_sc_hd__mux2_1 _1959_ ( .A0(\text_in_r\[0\] ), .A1(\text_in[0] ), .S(_1279_ ), .X(_0266_ ) );
sky130_fd_sc_hd__mux2_1 _1960_ ( .A0(\text_in_r\[1\] ), .A1(\text_in[1] ), .S(_1279_ ), .X(_0305_ ) );
sky130_fd_sc_hd__mux2_1 _1961_ ( .A0(\text_in_r\[2\] ), .A1(\text_in[2] ), .S(_1279_ ), .X(_0316_ ) );
sky130_fd_sc_hd__mux2_1 _1962_ ( .A0(\text_in_r\[3\] ), .A1(\text_in[3] ), .S(_1279_ ), .X(_0327_ ) );
sky130_fd_sc_hd__mux2_1 _1963_ ( .A0(\text_in_r\[4\] ), .A1(\text_in[4] ), .S(_1279_ ), .X(_0338_ ) );
sky130_fd_sc_hd__mux2_1 _1964_ ( .A0(\text_in_r\[5\] ), .A1(\text_in[5] ), .S(_1279_ ), .X(_0349_ ) );
sky130_fd_sc_hd__mux2_1 _1965_ ( .A0(\text_in_r\[6\] ), .A1(\text_in[6] ), .S(_1279_ ), .X(_0360_ ) );
sky130_fd_sc_hd__mux2_1 _1966_ ( .A0(\text_in_r\[7\] ), .A1(\text_in[7] ), .S(_1279_ ), .X(_0371_ ) );
sky130_fd_sc_hd__mux2_1 _1967_ ( .A0(\text_in_r\[8\] ), .A1(\text_in[8] ), .S(_1279_ ), .X(_0382_ ) );
sky130_fd_sc_hd__buf_2 _1968_ ( .A(_1278_ ), .X(_1293_ ) );
sky130_fd_sc_hd__mux2_1 _1969_ ( .A0(\text_in_r\[9\] ), .A1(\text_in[9] ), .S(_1293_ ), .X(_0393_ ) );
sky130_fd_sc_hd__mux2_1 _1970_ ( .A0(\text_in_r\[10\] ), .A1(\text_in[10] ), .S(_1293_ ), .X(_0277_ ) );
sky130_fd_sc_hd__mux2_1 _1971_ ( .A0(\text_in_r\[11\] ), .A1(\text_in[11] ), .S(_1293_ ), .X(_0288_ ) );
sky130_fd_sc_hd__mux2_1 _1972_ ( .A0(\text_in_r\[12\] ), .A1(\text_in[12] ), .S(_1293_ ), .X(_0297_ ) );
sky130_fd_sc_hd__mux2_1 _1973_ ( .A0(\text_in_r\[13\] ), .A1(\text_in[13] ), .S(_1293_ ), .X(_0298_ ) );
sky130_fd_sc_hd__mux2_1 _1974_ ( .A0(\text_in_r\[14\] ), .A1(\text_in[14] ), .S(_1293_ ), .X(_0299_ ) );
sky130_fd_sc_hd__mux2_1 _1975_ ( .A0(\text_in_r\[15\] ), .A1(\text_in[15] ), .S(_1293_ ), .X(_0300_ ) );
sky130_fd_sc_hd__mux2_1 _1976_ ( .A0(\text_in_r\[16\] ), .A1(\text_in[16] ), .S(_1293_ ), .X(_0301_ ) );
sky130_fd_sc_hd__mux2_1 _1977_ ( .A0(\text_in_r\[17\] ), .A1(\text_in[17] ), .S(_1293_ ), .X(_0302_ ) );
sky130_fd_sc_hd__mux2_1 _1978_ ( .A0(\text_in_r\[18\] ), .A1(\text_in[18] ), .S(_1293_ ), .X(_0303_ ) );
sky130_fd_sc_hd__buf_2 _1979_ ( .A(_1278_ ), .X(_1294_ ) );
sky130_fd_sc_hd__mux2_1 _1980_ ( .A0(\text_in_r\[19\] ), .A1(\text_in[19] ), .S(_1294_ ), .X(_0304_ ) );
sky130_fd_sc_hd__mux2_1 _1981_ ( .A0(\text_in_r\[20\] ), .A1(\text_in[20] ), .S(_1294_ ), .X(_0306_ ) );
sky130_fd_sc_hd__mux2_1 _1982_ ( .A0(\text_in_r\[21\] ), .A1(\text_in[21] ), .S(_1294_ ), .X(_0307_ ) );
sky130_fd_sc_hd__mux2_1 _1983_ ( .A0(\text_in_r\[22\] ), .A1(\text_in[22] ), .S(_1294_ ), .X(_0308_ ) );
sky130_fd_sc_hd__mux2_1 _1984_ ( .A0(\text_in_r\[23\] ), .A1(\text_in[23] ), .S(_1294_ ), .X(_0309_ ) );
sky130_fd_sc_hd__mux2_1 _1985_ ( .A0(\text_in_r\[24\] ), .A1(\text_in[24] ), .S(_1294_ ), .X(_0310_ ) );
sky130_fd_sc_hd__mux2_1 _1986_ ( .A0(\text_in_r\[25\] ), .A1(\text_in[25] ), .S(_1294_ ), .X(_0311_ ) );
sky130_fd_sc_hd__mux2_1 _1987_ ( .A0(\text_in_r\[26\] ), .A1(\text_in[26] ), .S(_1294_ ), .X(_0312_ ) );
sky130_fd_sc_hd__mux2_1 _1988_ ( .A0(\text_in_r\[27\] ), .A1(\text_in[27] ), .S(_1294_ ), .X(_0313_ ) );
sky130_fd_sc_hd__mux2_1 _1989_ ( .A0(\text_in_r\[28\] ), .A1(\text_in[28] ), .S(_1294_ ), .X(_0314_ ) );
sky130_fd_sc_hd__buf_2 _1990_ ( .A(_1278_ ), .X(_1295_ ) );
sky130_fd_sc_hd__mux2_1 _1991_ ( .A0(\text_in_r\[29\] ), .A1(\text_in[29] ), .S(_1295_ ), .X(_0315_ ) );
sky130_fd_sc_hd__mux2_1 _1992_ ( .A0(\text_in_r\[30\] ), .A1(\text_in[30] ), .S(_1295_ ), .X(_0317_ ) );
sky130_fd_sc_hd__mux2_1 _1993_ ( .A0(\text_in_r\[31\] ), .A1(\text_in[31] ), .S(_1295_ ), .X(_0318_ ) );
sky130_fd_sc_hd__mux2_1 _1994_ ( .A0(\text_in_r\[32\] ), .A1(\text_in[32] ), .S(_1295_ ), .X(_0319_ ) );
sky130_fd_sc_hd__mux2_1 _1995_ ( .A0(\text_in_r\[33\] ), .A1(\text_in[33] ), .S(_1295_ ), .X(_0320_ ) );
sky130_fd_sc_hd__mux2_1 _1996_ ( .A0(\text_in_r\[34\] ), .A1(\text_in[34] ), .S(_1295_ ), .X(_0321_ ) );
sky130_fd_sc_hd__mux2_1 _1997_ ( .A0(\text_in_r\[35\] ), .A1(\text_in[35] ), .S(_1295_ ), .X(_0322_ ) );
sky130_fd_sc_hd__mux2_1 _1998_ ( .A0(\text_in_r\[36\] ), .A1(\text_in[36] ), .S(_1295_ ), .X(_0323_ ) );
sky130_fd_sc_hd__mux2_1 _1999_ ( .A0(\text_in_r\[37\] ), .A1(\text_in[37] ), .S(_1295_ ), .X(_0324_ ) );
sky130_fd_sc_hd__mux2_1 _2000_ ( .A0(\text_in_r\[38\] ), .A1(\text_in[38] ), .S(_1295_ ), .X(_0325_ ) );
sky130_fd_sc_hd__buf_2 _2001_ ( .A(_1278_ ), .X(_1296_ ) );
sky130_fd_sc_hd__mux2_1 _2002_ ( .A0(\text_in_r\[39\] ), .A1(\text_in[39] ), .S(_1296_ ), .X(_0326_ ) );
sky130_fd_sc_hd__mux2_1 _2003_ ( .A0(\text_in_r\[40\] ), .A1(\text_in[40] ), .S(_1296_ ), .X(_0328_ ) );
sky130_fd_sc_hd__mux2_1 _2004_ ( .A0(\text_in_r\[41\] ), .A1(\text_in[41] ), .S(_1296_ ), .X(_0329_ ) );
sky130_fd_sc_hd__mux2_1 _2005_ ( .A0(\text_in_r\[42\] ), .A1(\text_in[42] ), .S(_1296_ ), .X(_0330_ ) );
sky130_fd_sc_hd__mux2_1 _2006_ ( .A0(\text_in_r\[43\] ), .A1(\text_in[43] ), .S(_1296_ ), .X(_0331_ ) );
sky130_fd_sc_hd__mux2_1 _2007_ ( .A0(\text_in_r\[44\] ), .A1(\text_in[44] ), .S(_1296_ ), .X(_0332_ ) );
sky130_fd_sc_hd__mux2_1 _2008_ ( .A0(\text_in_r\[45\] ), .A1(\text_in[45] ), .S(_1296_ ), .X(_0333_ ) );
sky130_fd_sc_hd__mux2_1 _2009_ ( .A0(\text_in_r\[46\] ), .A1(\text_in[46] ), .S(_1296_ ), .X(_0334_ ) );
sky130_fd_sc_hd__mux2_1 _2010_ ( .A0(\text_in_r\[47\] ), .A1(\text_in[47] ), .S(_1296_ ), .X(_0335_ ) );
sky130_fd_sc_hd__mux2_1 _2011_ ( .A0(\text_in_r\[48\] ), .A1(\text_in[48] ), .S(_1296_ ), .X(_0336_ ) );
sky130_fd_sc_hd__buf_2 _2012_ ( .A(_1278_ ), .X(_1297_ ) );
sky130_fd_sc_hd__mux2_1 _2013_ ( .A0(\text_in_r\[49\] ), .A1(\text_in[49] ), .S(_1297_ ), .X(_0337_ ) );
sky130_fd_sc_hd__mux2_1 _2014_ ( .A0(\text_in_r\[50\] ), .A1(\text_in[50] ), .S(_1297_ ), .X(_0339_ ) );
sky130_fd_sc_hd__mux2_1 _2015_ ( .A0(\text_in_r\[51\] ), .A1(\text_in[51] ), .S(_1297_ ), .X(_0340_ ) );
sky130_fd_sc_hd__mux2_1 _2016_ ( .A0(\text_in_r\[52\] ), .A1(\text_in[52] ), .S(_1297_ ), .X(_0341_ ) );
sky130_fd_sc_hd__mux2_1 _2017_ ( .A0(\text_in_r\[53\] ), .A1(\text_in[53] ), .S(_1297_ ), .X(_0342_ ) );
sky130_fd_sc_hd__mux2_1 _2018_ ( .A0(\text_in_r\[54\] ), .A1(\text_in[54] ), .S(_1297_ ), .X(_0343_ ) );
sky130_fd_sc_hd__mux2_1 _2019_ ( .A0(\text_in_r\[55\] ), .A1(\text_in[55] ), .S(_1297_ ), .X(_0344_ ) );
sky130_fd_sc_hd__mux2_1 _2020_ ( .A0(\text_in_r\[56\] ), .A1(\text_in[56] ), .S(_1297_ ), .X(_0345_ ) );
sky130_fd_sc_hd__mux2_1 _2021_ ( .A0(\text_in_r\[57\] ), .A1(\text_in[57] ), .S(_1297_ ), .X(_0346_ ) );
sky130_fd_sc_hd__mux2_1 _2022_ ( .A0(\text_in_r\[58\] ), .A1(\text_in[58] ), .S(_1297_ ), .X(_0347_ ) );
sky130_fd_sc_hd__buf_2 _2023_ ( .A(_1278_ ), .X(_1298_ ) );
sky130_fd_sc_hd__mux2_1 _2024_ ( .A0(\text_in_r\[59\] ), .A1(\text_in[59] ), .S(_1298_ ), .X(_0348_ ) );
sky130_fd_sc_hd__mux2_1 _2025_ ( .A0(\text_in_r\[60\] ), .A1(\text_in[60] ), .S(_1298_ ), .X(_0350_ ) );
sky130_fd_sc_hd__mux2_1 _2026_ ( .A0(\text_in_r\[61\] ), .A1(\text_in[61] ), .S(_1298_ ), .X(_0351_ ) );
sky130_fd_sc_hd__mux2_1 _2027_ ( .A0(\text_in_r\[62\] ), .A1(\text_in[62] ), .S(_1298_ ), .X(_0352_ ) );
sky130_fd_sc_hd__mux2_1 _2028_ ( .A0(\text_in_r\[63\] ), .A1(\text_in[63] ), .S(_1298_ ), .X(_0353_ ) );
sky130_fd_sc_hd__mux2_1 _2029_ ( .A0(\text_in_r\[64\] ), .A1(\text_in[64] ), .S(_1298_ ), .X(_0354_ ) );
sky130_fd_sc_hd__mux2_1 _2030_ ( .A0(\text_in_r\[65\] ), .A1(\text_in[65] ), .S(_1298_ ), .X(_0355_ ) );
sky130_fd_sc_hd__mux2_1 _2031_ ( .A0(\text_in_r\[66\] ), .A1(\text_in[66] ), .S(_1298_ ), .X(_0356_ ) );
sky130_fd_sc_hd__mux2_1 _2032_ ( .A0(\text_in_r\[67\] ), .A1(\text_in[67] ), .S(_1298_ ), .X(_0357_ ) );
sky130_fd_sc_hd__mux2_1 _2033_ ( .A0(\text_in_r\[68\] ), .A1(\text_in[68] ), .S(_1298_ ), .X(_0358_ ) );
sky130_fd_sc_hd__mux2_1 _2035_ ( .A0(\text_in_r\[69\] ), .A1(\text_in[69] ), .S(_1295_ ), .X(_0359_ ) );
sky130_fd_sc_hd__mux2_1 _2036_ ( .A0(\text_in_r\[70\] ), .A1(\text_in[70] ), .S(_1295_ ), .X(_0361_ ) );
sky130_fd_sc_hd__mux2_1 _2037_ ( .A0(\text_in_r\[71\] ), .A1(\text_in[71] ), .S(_1295_ ), .X(_0362_ ) );
sky130_fd_sc_hd__mux2_1 _2038_ ( .A0(\text_in_r\[72\] ), .A1(\text_in[72] ), .S(_1295_ ), .X(_0363_ ) );
sky130_fd_sc_hd__mux2_1 _2039_ ( .A0(\text_in_r\[73\] ), .A1(\text_in[73] ), .S(_1295_ ), .X(_0364_ ) );
sky130_fd_sc_hd__mux2_1 _2040_ ( .A0(\text_in_r\[74\] ), .A1(\text_in[74] ), .S(_1295_ ), .X(_0365_ ) );
sky130_fd_sc_hd__mux2_1 _2041_ ( .A0(\text_in_r\[75\] ), .A1(\text_in[75] ), .S(_1295_ ), .X(_0366_ ) );
sky130_fd_sc_hd__mux2_1 _2042_ ( .A0(\text_in_r\[76\] ), .A1(\text_in[76] ), .S(_1295_ ), .X(_0367_ ) );
sky130_fd_sc_hd__mux2_1 _2043_ ( .A0(\text_in_r\[77\] ), .A1(\text_in[77] ), .S(_1295_ ), .X(_0368_ ) );
sky130_fd_sc_hd__mux2_1 _2044_ ( .A0(\text_in_r\[78\] ), .A1(\text_in[78] ), .S(_1295_ ), .X(_0369_ ) );
sky130_fd_sc_hd__buf_2 _2045_ ( .A(_1278_ ), .X(_0529_ ) );
sky130_fd_sc_hd__mux2_1 _2046_ ( .A0(\text_in_r\[79\] ), .A1(\text_in[79] ), .S(_0529_ ), .X(_0370_ ) );
sky130_fd_sc_hd__mux2_1 _2047_ ( .A0(\text_in_r\[80\] ), .A1(\text_in[80] ), .S(_0529_ ), .X(_0372_ ) );
sky130_fd_sc_hd__mux2_1 _2048_ ( .A0(\text_in_r\[81\] ), .A1(\text_in[81] ), .S(_0529_ ), .X(_0373_ ) );
sky130_fd_sc_hd__mux2_1 _2049_ ( .A0(\text_in_r\[82\] ), .A1(\text_in[82] ), .S(_0529_ ), .X(_0374_ ) );
sky130_fd_sc_hd__mux2_1 _2050_ ( .A0(\text_in_r\[83\] ), .A1(\text_in[83] ), .S(_0529_ ), .X(_0375_ ) );
sky130_fd_sc_hd__mux2_1 _2051_ ( .A0(\text_in_r\[84\] ), .A1(\text_in[84] ), .S(_0529_ ), .X(_0376_ ) );
sky130_fd_sc_hd__mux2_1 _2052_ ( .A0(\text_in_r\[85\] ), .A1(\text_in[85] ), .S(_0529_ ), .X(_0377_ ) );
sky130_fd_sc_hd__mux2_1 _2053_ ( .A0(\text_in_r\[86\] ), .A1(\text_in[86] ), .S(_0529_ ), .X(_0378_ ) );
sky130_fd_sc_hd__mux2_1 _2054_ ( .A0(\text_in_r\[87\] ), .A1(\text_in[87] ), .S(_0529_ ), .X(_0379_ ) );
sky130_fd_sc_hd__mux2_1 _2055_ ( .A0(\text_in_r\[88\] ), .A1(\text_in[88] ), .S(_0529_ ), .X(_0380_ ) );
sky130_fd_sc_hd__buf_2 _2056_ ( .A(_1278_ ), .X(_0530_ ) );
sky130_fd_sc_hd__mux2_1 _2057_ ( .A0(\text_in_r\[89\] ), .A1(\text_in[89] ), .S(_0530_ ), .X(_0381_ ) );
sky130_fd_sc_hd__mux2_1 _2058_ ( .A0(\text_in_r\[90\] ), .A1(\text_in[90] ), .S(_0530_ ), .X(_0383_ ) );
sky130_fd_sc_hd__mux2_1 _2059_ ( .A0(\text_in_r\[91\] ), .A1(\text_in[91] ), .S(_0530_ ), .X(_0384_ ) );
sky130_fd_sc_hd__mux2_1 _2060_ ( .A0(\text_in_r\[92\] ), .A1(\text_in[92] ), .S(_0530_ ), .X(_0385_ ) );
sky130_fd_sc_hd__mux2_1 _2061_ ( .A0(\text_in_r\[93\] ), .A1(\text_in[93] ), .S(_0530_ ), .X(_0386_ ) );
sky130_fd_sc_hd__mux2_1 _2062_ ( .A0(\text_in_r\[94\] ), .A1(\text_in[94] ), .S(_0530_ ), .X(_0387_ ) );
sky130_fd_sc_hd__mux2_1 _2063_ ( .A0(\text_in_r\[95\] ), .A1(\text_in[95] ), .S(_0530_ ), .X(_0388_ ) );
sky130_fd_sc_hd__mux2_1 _2064_ ( .A0(\text_in_r\[96\] ), .A1(\text_in[96] ), .S(_0530_ ), .X(_0389_ ) );
sky130_fd_sc_hd__mux2_1 _2065_ ( .A0(\text_in_r\[97\] ), .A1(\text_in[97] ), .S(_0530_ ), .X(_0390_ ) );
sky130_fd_sc_hd__mux2_1 _2066_ ( .A0(\text_in_r\[98\] ), .A1(\text_in[98] ), .S(_0530_ ), .X(_0391_ ) );
sky130_fd_sc_hd__buf_2 _2067_ ( .A(ld ), .X(_0531_ ) );
sky130_fd_sc_hd__mux2_1 _2068_ ( .A0(\text_in_r\[99\] ), .A1(\text_in[99] ), .S(_0531_ ), .X(_0392_ ) );
sky130_fd_sc_hd__mux2_1 _2069_ ( .A0(\text_in_r\[100\] ), .A1(\text_in[100] ), .S(_0531_ ), .X(_0267_ ) );
sky130_fd_sc_hd__mux2_1 _2070_ ( .A0(\text_in_r\[101\] ), .A1(\text_in[101] ), .S(_0531_ ), .X(_0268_ ) );
sky130_fd_sc_hd__mux2_1 _2071_ ( .A0(\text_in_r\[102\] ), .A1(\text_in[102] ), .S(_0531_ ), .X(_0269_ ) );
sky130_fd_sc_hd__mux2_1 _2072_ ( .A0(\text_in_r\[103\] ), .A1(\text_in[103] ), .S(_0531_ ), .X(_0270_ ) );
sky130_fd_sc_hd__mux2_1 _2073_ ( .A0(\text_in_r\[104\] ), .A1(\text_in[104] ), .S(_0531_ ), .X(_0271_ ) );
sky130_fd_sc_hd__mux2_1 _2074_ ( .A0(\text_in_r\[105\] ), .A1(\text_in[105] ), .S(_0531_ ), .X(_0272_ ) );
sky130_fd_sc_hd__mux2_1 _2075_ ( .A0(\text_in_r\[106\] ), .A1(\text_in[106] ), .S(_0531_ ), .X(_0273_ ) );
sky130_fd_sc_hd__mux2_1 _2076_ ( .A0(\text_in_r\[107\] ), .A1(\text_in[107] ), .S(_0531_ ), .X(_0274_ ) );
sky130_fd_sc_hd__mux2_1 _2077_ ( .A0(\text_in_r\[108\] ), .A1(\text_in[108] ), .S(_0531_ ), .X(_0275_ ) );
sky130_fd_sc_hd__buf_2 _2078_ ( .A(ld ), .X(_0532_ ) );
sky130_fd_sc_hd__mux2_1 _2079_ ( .A0(\text_in_r\[109\] ), .A1(\text_in[109] ), .S(_0532_ ), .X(_0276_ ) );
sky130_fd_sc_hd__mux2_1 _2080_ ( .A0(\text_in_r\[110\] ), .A1(\text_in[110] ), .S(_0532_ ), .X(_0278_ ) );
sky130_fd_sc_hd__mux2_1 _2081_ ( .A0(\text_in_r\[111\] ), .A1(\text_in[111] ), .S(_0532_ ), .X(_0279_ ) );
sky130_fd_sc_hd__mux2_1 _2082_ ( .A0(\text_in_r\[112\] ), .A1(\text_in[112] ), .S(_0532_ ), .X(_0280_ ) );
sky130_fd_sc_hd__mux2_1 _2083_ ( .A0(\text_in_r\[113\] ), .A1(\text_in[113] ), .S(_0532_ ), .X(_0281_ ) );
sky130_fd_sc_hd__mux2_1 _2084_ ( .A0(\text_in_r\[114\] ), .A1(\text_in[114] ), .S(_0532_ ), .X(_0282_ ) );
sky130_fd_sc_hd__mux2_1 _2085_ ( .A0(\text_in_r\[115\] ), .A1(\text_in[115] ), .S(_0532_ ), .X(_0283_ ) );
sky130_fd_sc_hd__mux2_1 _2086_ ( .A0(\text_in_r\[116\] ), .A1(\text_in[116] ), .S(_0532_ ), .X(_0284_ ) );
sky130_fd_sc_hd__mux2_1 _2087_ ( .A0(\text_in_r\[117\] ), .A1(\text_in[117] ), .S(_0532_ ), .X(_0285_ ) );
sky130_fd_sc_hd__mux2_1 _2088_ ( .A0(\text_in_r\[118\] ), .A1(\text_in[118] ), .S(_0532_ ), .X(_0286_ ) );
sky130_fd_sc_hd__mux2_1 _2089_ ( .A0(\text_in_r\[119\] ), .A1(\text_in[119] ), .S(_1282_ ), .X(_0287_ ) );
sky130_fd_sc_hd__mux2_1 _2090_ ( .A0(\text_in_r\[120\] ), .A1(\text_in[120] ), .S(_1282_ ), .X(_0289_ ) );
sky130_fd_sc_hd__mux2_1 _2091_ ( .A0(\text_in_r\[121\] ), .A1(\text_in[121] ), .S(_1282_ ), .X(_0290_ ) );
sky130_fd_sc_hd__mux2_1 _2092_ ( .A0(\text_in_r\[122\] ), .A1(\text_in[122] ), .S(_1282_ ), .X(_0291_ ) );
sky130_fd_sc_hd__mux2_1 _2093_ ( .A0(\text_in_r\[123\] ), .A1(\text_in[123] ), .S(_1282_ ), .X(_0292_ ) );
sky130_fd_sc_hd__mux2_1 _2094_ ( .A0(\text_in_r\[124\] ), .A1(\text_in[124] ), .S(_1282_ ), .X(_0293_ ) );
sky130_fd_sc_hd__mux2_1 _2095_ ( .A0(\text_in_r\[125\] ), .A1(\text_in[125] ), .S(_1282_ ), .X(_0294_ ) );
sky130_fd_sc_hd__mux2_1 _2096_ ( .A0(\text_in_r\[126\] ), .A1(\text_in[126] ), .S(_1282_ ), .X(_0295_ ) );
sky130_fd_sc_hd__mux2_1 _2097_ ( .A0(\text_in_r\[127\] ), .A1(\text_in[127] ), .S(_1282_ ), .X(_0296_ ) );
sky130_fd_sc_hd__nor2_1 _2098_ ( .A(_1280_ ), .B(_1284_ ), .Y(_0265_ ) );
sky130_fd_sc_hd__xnor2_1 _2099_ ( .A(\us11\/_0008_ ), .B(\us22\/_0008_ ), .Y(_0533_ ) );
sky130_fd_sc_hd__xor2_1 _2100_ ( .A(_1379_ ), .B(\us33\/_0008_ ), .X(_0534_ ) );
sky130_fd_sc_hd__xor3_1 _2101_ ( .A(\us00\/_0015_ ), .B(_0533_ ), .C(_0534_ ), .X(_0535_ ) );
sky130_fd_sc_hd__clkbuf_1 _2102_ ( .A(ld_r ), .X(_0536_ ) );
sky130_fd_sc_hd__inv_2 _2103_ ( .A(_0536_ ), .Y(_0537_ ) );
sky130_fd_sc_hd__clkbuf_1 _2104_ ( .A(_0537_ ), .X(_0538_ ) );
sky130_fd_sc_hd__nand2_1 _2105_ ( .A(_0535_ ), .B(_0538_ ), .Y(_0539_ ) );
sky130_fd_sc_hd__or2b_1 _2107_ ( .A(\text_in_r\[120\] ), .B_N(_0549_ ), .X(_0541_ ) );
sky130_fd_sc_hd__nand2_1 _2108_ ( .A(_0539_ ), .B(_0541_ ), .Y(_0542_ ) );
sky130_fd_sc_hd__xnor2_1 _2109_ ( .A(\w0\[24\] ), .B(_0542_ ), .Y(_1300_ ) );
sky130_fd_sc_hd__xor2_1 _2110_ ( .A(\us00\/_0015_ ), .B(\us00\/_0008_ ), .X(_0543_ ) );
sky130_fd_sc_hd__xor2_1 _2111_ ( .A(\us22\/_0009_ ), .B(\us33\/_0009_ ), .X(_0544_ ) );
sky130_fd_sc_hd__xnor3_1 _2112_ ( .A(_1379_ ), .B(\us11\/_0008_ ), .C(_1373_ ), .X(_0545_ ) );
sky130_fd_sc_hd__xnor3_1 _2113_ ( .A(_0543_ ), .B(_0544_ ), .C(_0545_ ), .X(_0546_ ) );
sky130_fd_sc_hd__clkbuf_1 _2114_ ( .A(_0537_ ), .X(_0547_ ) );
sky130_fd_sc_hd__nand2_1 _2115_ ( .A(_0546_ ), .B(_0547_ ), .Y(_0548_ ) );
sky130_fd_sc_hd__buf_2 _2116_ ( .A(_0536_ ), .X(_0549_ ) );
sky130_fd_sc_hd__buf_2 _2117_ ( .A(_0549_ ), .X(_0550_ ) );
sky130_fd_sc_hd__nand2_1 _2118_ ( .A(\text_in_r\[121\] ), .B(_0550_ ), .Y(_0551_ ) );
sky130_fd_sc_hd__nand2_1 _2119_ ( .A(_0548_ ), .B(_0551_ ), .Y(_0552_ ) );
sky130_fd_sc_hd__xor2_1 _2120_ ( .A(\w0\[25\] ), .B(_0552_ ), .X(_1301_ ) );
sky130_fd_sc_hd__and2_0 _2122_ ( .A(\text_in_r\[122\] ), .B(ld_r ), .X(_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 _2123_ ( .A(_0549_ ), .X(_0555_ ) );
sky130_fd_sc_hd__inv_1 _2124_ ( .A(\us22\/_0010_ ), .Y(_0556_ ) );
sky130_fd_sc_hd__xnor2_1 _2125_ ( .A(_1373_ ), .B(\us00\/_0009_ ), .Y(_0557_ ) );
sky130_fd_sc_hd__xor2_1 _2126_ ( .A(\us11\/_0010_ ), .B(\us33\/_0010_ ), .X(_0558_ ) );
sky130_fd_sc_hd__xnor3_1 _2127_ ( .A(_0556_ ), .B(_0557_ ), .C(_0558_ ), .X(_0559_ ) );
sky130_fd_sc_hd__nor2_1 _2128_ ( .A(_0555_ ), .B(_0559_ ), .Y(_0560_ ) );
sky130_fd_sc_hd__nor2_1 _2129_ ( .A(_0554_ ), .B(_0560_ ), .Y(_0561_ ) );
sky130_fd_sc_hd__xnor2_1 _2130_ ( .A(\w0\[26\] ), .B(_0561_ ), .Y(_1302_ ) );
sky130_fd_sc_hd__clkbuf_1 _2131_ ( .A(ld_r ), .X(_0562_ ) );
sky130_fd_sc_hd__and2b_1 _2132_ ( .A_N(\text_in_r\[123\] ), .B(_0562_ ), .X(_0563_ ) );
sky130_fd_sc_hd__clkbuf_1 _2133_ ( .A(_0549_ ), .X(_0564_ ) );
sky130_fd_sc_hd__xor2_1 _2134_ ( .A(\us00\/_0015_ ), .B(\us00\/_0010_ ), .X(_0565_ ) );
sky130_fd_sc_hd__xor2_1 _2135_ ( .A(\us22\/_0011_ ), .B(\us33\/_0011_ ), .X(_0566_ ) );
sky130_fd_sc_hd__xnor3_1 _2136_ ( .A(_1379_ ), .B(\us11\/_0010_ ), .C(\us11\/_0011_ ), .X(_0567_ ) );
sky130_fd_sc_hd__xnor3_1 _2137_ ( .A(_0565_ ), .B(_0566_ ), .C(_0567_ ), .X(_0568_ ) );
sky130_fd_sc_hd__nor2_1 _2138_ ( .A(_0564_ ), .B(_0568_ ), .Y(_0569_ ) );
sky130_fd_sc_hd__nor2_1 _2139_ ( .A(_0563_ ), .B(_0569_ ), .Y(_0570_ ) );
sky130_fd_sc_hd__xor2_1 _2140_ ( .A(\w0\[27\] ), .B(_0570_ ), .X(_1303_ ) );
sky130_fd_sc_hd__and2b_1 _2141_ ( .A_N(\text_in_r\[124\] ), .B(_0562_ ), .X(_0571_ ) );
sky130_fd_sc_hd__xnor2_1 _2142_ ( .A(\us00\/_0015_ ), .B(\us00\/_0011_ ), .Y(_0572_ ) );
sky130_fd_sc_hd__xnor2_1 _2143_ ( .A(\us22\/_0012_ ), .B(\us33\/_0012_ ), .Y(_0573_ ) );
sky130_fd_sc_hd__xnor3_1 _2144_ ( .A(_1379_ ), .B(\us11\/_0011_ ), .C(\us11\/_0012_ ), .X(_0574_ ) );
sky130_fd_sc_hd__xnor3_1 _2145_ ( .A(_0572_ ), .B(_0573_ ), .C(_0574_ ), .X(_0575_ ) );
sky130_fd_sc_hd__nor2_1 _2146_ ( .A(_0564_ ), .B(_0575_ ), .Y(_0576_ ) );
sky130_fd_sc_hd__nor2_1 _2147_ ( .A(_0571_ ), .B(_0576_ ), .Y(_0577_ ) );
sky130_fd_sc_hd__xor2_1 _2148_ ( .A(\w0\[28\] ), .B(_0577_ ), .X(_1304_ ) );
sky130_fd_sc_hd__xnor2_1 _2149_ ( .A(_1377_ ), .B(\us22\/_0013_ ), .Y(_0578_ ) );
sky130_fd_sc_hd__xnor2_1 _2150_ ( .A(\us11\/_0012_ ), .B(\us00\/_0012_ ), .Y(_0579_ ) );
sky130_fd_sc_hd__xnor3_1 _2151_ ( .A(\us33\/_0013_ ), .B(_0578_ ), .C(_0579_ ), .X(_0580_ ) );
sky130_fd_sc_hd__nand2_1 _2152_ ( .A(_0580_ ), .B(_0538_ ), .Y(_0581_ ) );
sky130_fd_sc_hd__or2b_1 _2153_ ( .A(\text_in_r\[125\] ), .B_N(_0549_ ), .X(_0582_ ) );
sky130_fd_sc_hd__nand2_1 _2154_ ( .A(_0581_ ), .B(_0582_ ), .Y(_0583_ ) );
sky130_fd_sc_hd__xnor2_1 _2155_ ( .A(\w0\[29\] ), .B(_0583_ ), .Y(_1305_ ) );
sky130_fd_sc_hd__and2_0 _2156_ ( .A(\text_in_r\[126\] ), .B(ld_r ), .X(_0584_ ) );
sky130_fd_sc_hd__xor2_1 _2157_ ( .A(_1377_ ), .B(\us00\/_0013_ ), .X(_0585_ ) );
sky130_fd_sc_hd__xor2_1 _2158_ ( .A(\us11\/_0014_ ), .B(\us33\/_0014_ ), .X(_0586_ ) );
sky130_fd_sc_hd__xnor3_1 _2159_ ( .A(\us22\/_0014_ ), .B(_0585_ ), .C(_0586_ ), .X(_0587_ ) );
sky130_fd_sc_hd__nor2_1 _2160_ ( .A(_0555_ ), .B(_0587_ ), .Y(_0588_ ) );
sky130_fd_sc_hd__nor2_1 _2161_ ( .A(_0584_ ), .B(_0588_ ), .Y(_0589_ ) );
sky130_fd_sc_hd__xnor2_1 _2162_ ( .A(\w0\[30\] ), .B(_0589_ ), .Y(_1306_ ) );
sky130_fd_sc_hd__xnor2_1 _2164_ ( .A(\us11\/_0014_ ), .B(\us33\/_0015_ ), .Y(_0591_ ) );
sky130_fd_sc_hd__xnor2_1 _2165_ ( .A(\us00\/_0014_ ), .B(\us22\/_0015_ ), .Y(_0592_ ) );
sky130_fd_sc_hd__xnor3_1 _2166_ ( .A(_1379_ ), .B(_0591_ ), .C(_0592_ ), .X(_0593_ ) );
sky130_fd_sc_hd__nand2_1 _2167_ ( .A(_0593_ ), .B(_0538_ ), .Y(_0594_ ) );
sky130_fd_sc_hd__or2b_1 _2168_ ( .A(\text_in_r\[127\] ), .B_N(_0549_ ), .X(_0595_ ) );
sky130_fd_sc_hd__nand2_1 _2169_ ( .A(_0594_ ), .B(_0595_ ), .Y(_0596_ ) );
sky130_fd_sc_hd__xnor2_1 _2170_ ( .A(\w0\[31\] ), .B(_0596_ ), .Y(_1307_ ) );
sky130_fd_sc_hd__and2_0 _2171_ ( .A(\text_in_r\[88\] ), .B(ld_r ), .X(_0597_ ) );
sky130_fd_sc_hd__inv_1 _2172_ ( .A(\us01\/_0015_ ), .Y(_0598_ ) );
sky130_fd_sc_hd__xnor2_1 _2173_ ( .A(\us12\/_0008_ ), .B(\us23\/_0008_ ), .Y(_0599_ ) );
sky130_fd_sc_hd__xor2_1 _2174_ ( .A(\us12\/_0015_ ), .B(\us30\/_0008_ ), .X(_0600_ ) );
sky130_fd_sc_hd__xnor3_1 _2175_ ( .A(_0598_ ), .B(_0599_ ), .C(_0600_ ), .X(_0601_ ) );
sky130_fd_sc_hd__nor2_1 _2176_ ( .A(_0555_ ), .B(_0601_ ), .Y(_0602_ ) );
sky130_fd_sc_hd__nor2_1 _2177_ ( .A(_0597_ ), .B(_0602_ ), .Y(_0603_ ) );
sky130_fd_sc_hd__xnor2_1 _2178_ ( .A(\w1\[24\] ), .B(_0603_ ), .Y(_1316_ ) );
sky130_fd_sc_hd__xor2_1 _2179_ ( .A(\us01\/_0015_ ), .B(\us01\/_0008_ ), .X(_0604_ ) );
sky130_fd_sc_hd__xor2_1 _2180_ ( .A(\us23\/_0009_ ), .B(\us30\/_0009_ ), .X(_0605_ ) );
sky130_fd_sc_hd__xnor3_1 _2181_ ( .A(\us12\/_0015_ ), .B(\us12\/_0008_ ), .C(\us12\/_0009_ ), .X(_0606_ ) );
sky130_fd_sc_hd__xnor3_1 _2182_ ( .A(_0604_ ), .B(_0605_ ), .C(_0606_ ), .X(_0607_ ) );
sky130_fd_sc_hd__nand2_1 _2183_ ( .A(_0607_ ), .B(_0547_ ), .Y(_0608_ ) );
sky130_fd_sc_hd__nand2_1 _2184_ ( .A(\text_in_r\[89\] ), .B(_0550_ ), .Y(_0609_ ) );
sky130_fd_sc_hd__nand2_1 _2185_ ( .A(_0608_ ), .B(_0609_ ), .Y(_0610_ ) );
sky130_fd_sc_hd__xor2_1 _2186_ ( .A(\w1\[25\] ), .B(_0610_ ), .X(_1317_ ) );
sky130_fd_sc_hd__and2_0 _2187_ ( .A(\text_in_r\[90\] ), .B(ld_r ), .X(_0611_ ) );
sky130_fd_sc_hd__inv_1 _2188_ ( .A(\us23\/_0010_ ), .Y(_0612_ ) );
sky130_fd_sc_hd__xnor2_1 _2189_ ( .A(\us12\/_0009_ ), .B(\us01\/_0009_ ), .Y(_0613_ ) );
sky130_fd_sc_hd__xor2_1 _2190_ ( .A(\us12\/_0010_ ), .B(\us30\/_0010_ ), .X(_0614_ ) );
sky130_fd_sc_hd__xnor3_1 _2191_ ( .A(_0612_ ), .B(_0613_ ), .C(_0614_ ), .X(_0615_ ) );
sky130_fd_sc_hd__nor2_1 _2192_ ( .A(_0555_ ), .B(_0615_ ), .Y(_0616_ ) );
sky130_fd_sc_hd__nor2_1 _2193_ ( .A(_0611_ ), .B(_0616_ ), .Y(_0617_ ) );
sky130_fd_sc_hd__xnor2_1 _2194_ ( .A(\w1\[26\] ), .B(_0617_ ), .Y(_1318_ ) );
sky130_fd_sc_hd__and2b_1 _2195_ ( .A_N(\text_in_r\[91\] ), .B(_0562_ ), .X(_0618_ ) );
sky130_fd_sc_hd__xor2_1 _2196_ ( .A(\us01\/_0015_ ), .B(\us01\/_0010_ ), .X(_0619_ ) );
sky130_fd_sc_hd__xor2_1 _2197_ ( .A(\us23\/_0011_ ), .B(\us30\/_0011_ ), .X(_0620_ ) );
sky130_fd_sc_hd__xnor3_1 _2198_ ( .A(\us12\/_0015_ ), .B(\us12\/_0010_ ), .C(\us12\/_0011_ ), .X(_0621_ ) );
sky130_fd_sc_hd__xnor3_1 _2199_ ( .A(_0619_ ), .B(_0620_ ), .C(_0621_ ), .X(_0622_ ) );
sky130_fd_sc_hd__nor2_1 _2200_ ( .A(_0564_ ), .B(_0622_ ), .Y(_0623_ ) );
sky130_fd_sc_hd__nor2_1 _2201_ ( .A(_0618_ ), .B(_0623_ ), .Y(_0624_ ) );
sky130_fd_sc_hd__xor2_1 _2202_ ( .A(\w1\[27\] ), .B(_0624_ ), .X(_1319_ ) );
sky130_fd_sc_hd__xnor2_1 _2203_ ( .A(\us01\/_0015_ ), .B(\us01\/_0011_ ), .Y(_0625_ ) );
sky130_fd_sc_hd__xnor2_1 _2204_ ( .A(\us23\/_0012_ ), .B(\us30\/_0012_ ), .Y(_0626_ ) );
sky130_fd_sc_hd__xnor3_1 _2205_ ( .A(\us12\/_0015_ ), .B(\us12\/_0011_ ), .C(\us12\/_0012_ ), .X(_0627_ ) );
sky130_fd_sc_hd__xnor3_1 _2206_ ( .A(_0625_ ), .B(_0626_ ), .C(_0627_ ), .X(_0628_ ) );
sky130_fd_sc_hd__nand2_1 _2207_ ( .A(_0628_ ), .B(_0547_ ), .Y(_0629_ ) );
sky130_fd_sc_hd__nand2_1 _2208_ ( .A(\text_in_r\[92\] ), .B(_0550_ ), .Y(_0630_ ) );
sky130_fd_sc_hd__nand2_1 _2209_ ( .A(_0629_ ), .B(_0630_ ), .Y(_0631_ ) );
sky130_fd_sc_hd__xor2_1 _2210_ ( .A(\w1\[28\] ), .B(_0631_ ), .X(_1320_ ) );
sky130_fd_sc_hd__xnor2_1 _2211_ ( .A(\us12\/_0013_ ), .B(\us23\/_0013_ ), .Y(_0632_ ) );
sky130_fd_sc_hd__xnor2_1 _2212_ ( .A(\us12\/_0012_ ), .B(\us01\/_0012_ ), .Y(_0633_ ) );
sky130_fd_sc_hd__xnor3_1 _2213_ ( .A(\us30\/_0013_ ), .B(_0632_ ), .C(_0633_ ), .X(_0634_ ) );
sky130_fd_sc_hd__nand2_1 _2214_ ( .A(_0634_ ), .B(_0538_ ), .Y(_0635_ ) );
sky130_fd_sc_hd__or2b_1 _2215_ ( .A(\text_in_r\[93\] ), .B_N(_0549_ ), .X(_0636_ ) );
sky130_fd_sc_hd__nand2_1 _2216_ ( .A(_0635_ ), .B(_0636_ ), .Y(_0637_ ) );
sky130_fd_sc_hd__xnor2_1 _2217_ ( .A(\w1\[29\] ), .B(_0637_ ), .Y(_1321_ ) );
sky130_fd_sc_hd__xor2_1 _2218_ ( .A(\us12\/_0013_ ), .B(\us01\/_0013_ ), .X(_0638_ ) );
sky130_fd_sc_hd__xor2_1 _2219_ ( .A(\us12\/_0014_ ), .B(\us30\/_0014_ ), .X(_0639_ ) );
sky130_fd_sc_hd__xnor3_1 _2220_ ( .A(\us23\/_0014_ ), .B(_0638_ ), .C(_0639_ ), .X(_0640_ ) );
sky130_fd_sc_hd__nand2_1 _2221_ ( .A(_0640_ ), .B(_0538_ ), .Y(_0641_ ) );
sky130_fd_sc_hd__or2b_1 _2223_ ( .A(\text_in_r\[94\] ), .B_N(_0911_ ), .X(_0643_ ) );
sky130_fd_sc_hd__nand2_1 _2224_ ( .A(_0641_ ), .B(_0643_ ), .Y(_0644_ ) );
sky130_fd_sc_hd__xnor2_1 _2225_ ( .A(\w1\[30\] ), .B(_0644_ ), .Y(_1322_ ) );
sky130_fd_sc_hd__and2_0 _2226_ ( .A(\text_in_r\[95\] ), .B(ld_r ), .X(_0645_ ) );
sky130_fd_sc_hd__clkbuf_1 _2227_ ( .A(\us30\/_0015_ ), .X(_0646_ ) );
sky130_fd_sc_hd__xnor2_1 _2228_ ( .A(\us12\/_0014_ ), .B(_0646_ ), .Y(_0647_ ) );
sky130_fd_sc_hd__xnor2_1 _2229_ ( .A(\us01\/_0014_ ), .B(\us23\/_0015_ ), .Y(_0648_ ) );
sky130_fd_sc_hd__xnor3_1 _2230_ ( .A(\us12\/_0015_ ), .B(_0647_ ), .C(_0648_ ), .X(_0649_ ) );
sky130_fd_sc_hd__nor2_1 _2231_ ( .A(_0555_ ), .B(_0649_ ), .Y(_0650_ ) );
sky130_fd_sc_hd__nor2_1 _2232_ ( .A(_0645_ ), .B(_0650_ ), .Y(_0651_ ) );
sky130_fd_sc_hd__xnor2_1 _2233_ ( .A(\w1\[31\] ), .B(_0651_ ), .Y(_1323_ ) );
sky130_fd_sc_hd__and2_0 _2234_ ( .A(\text_in_r\[56\] ), .B(ld_r ), .X(_0652_ ) );
sky130_fd_sc_hd__clkbuf_1 _2235_ ( .A(_0549_ ), .X(_0653_ ) );
sky130_fd_sc_hd__inv_1 _2236_ ( .A(\us02\/_0015_ ), .Y(_0654_ ) );
sky130_fd_sc_hd__xnor2_1 _2237_ ( .A(\us13\/_0008_ ), .B(\us20\/_0008_ ), .Y(_0655_ ) );
sky130_fd_sc_hd__xor2_1 _2238_ ( .A(_1419_ ), .B(\us31\/_0008_ ), .X(_0656_ ) );
sky130_fd_sc_hd__xnor3_1 _2239_ ( .A(_0654_ ), .B(_0655_ ), .C(_0656_ ), .X(_0657_ ) );
sky130_fd_sc_hd__nor2_1 _2240_ ( .A(_0653_ ), .B(_0657_ ), .Y(_0658_ ) );
sky130_fd_sc_hd__nor2_1 _2241_ ( .A(_0652_ ), .B(_0658_ ), .Y(_0659_ ) );
sky130_fd_sc_hd__xnor2_1 _2242_ ( .A(\w2\[24\] ), .B(_0659_ ), .Y(_1332_ ) );
sky130_fd_sc_hd__xor2_1 _2243_ ( .A(\us02\/_0015_ ), .B(\us02\/_0008_ ), .X(_0660_ ) );
sky130_fd_sc_hd__xor2_1 _2244_ ( .A(\us20\/_0009_ ), .B(\us31\/_0009_ ), .X(_0661_ ) );
sky130_fd_sc_hd__xnor3_1 _2245_ ( .A(_1419_ ), .B(\us13\/_0008_ ), .C(\us13\/_0009_ ), .X(_0662_ ) );
sky130_fd_sc_hd__xnor3_1 _2246_ ( .A(_0660_ ), .B(_0661_ ), .C(_0662_ ), .X(_0663_ ) );
sky130_fd_sc_hd__clkbuf_1 _2247_ ( .A(_0537_ ), .X(_0664_ ) );
sky130_fd_sc_hd__nand2_1 _2248_ ( .A(_0663_ ), .B(_0664_ ), .Y(_0665_ ) );
sky130_fd_sc_hd__nand2_1 _2249_ ( .A(\text_in_r\[57\] ), .B(_0550_ ), .Y(_0666_ ) );
sky130_fd_sc_hd__nand2_1 _2250_ ( .A(_0665_ ), .B(_0666_ ), .Y(_0667_ ) );
sky130_fd_sc_hd__xor2_1 _2251_ ( .A(\w2\[25\] ), .B(_0667_ ), .X(_1333_ ) );
sky130_fd_sc_hd__inv_1 _2252_ ( .A(\us20\/_0010_ ), .Y(_0668_ ) );
sky130_fd_sc_hd__xnor2_1 _2253_ ( .A(\us13\/_0009_ ), .B(\us02\/_0009_ ), .Y(_0669_ ) );
sky130_fd_sc_hd__xor2_1 _2254_ ( .A(\us13\/_0010_ ), .B(\us31\/_0010_ ), .X(_0670_ ) );
sky130_fd_sc_hd__xnor3_1 _2255_ ( .A(_0668_ ), .B(_0669_ ), .C(_0670_ ), .X(_0671_ ) );
sky130_fd_sc_hd__nand2_1 _2256_ ( .A(_0671_ ), .B(_0538_ ), .Y(_0672_ ) );
sky130_fd_sc_hd__or2b_1 _2257_ ( .A(\text_in_r\[58\] ), .B_N(_0911_ ), .X(_0673_ ) );
sky130_fd_sc_hd__nand2_1 _2258_ ( .A(_0672_ ), .B(_0673_ ), .Y(_0674_ ) );
sky130_fd_sc_hd__xnor2_1 _2259_ ( .A(\w2\[26\] ), .B(_0674_ ), .Y(_1334_ ) );
sky130_fd_sc_hd__xor2_1 _2260_ ( .A(\us02\/_0015_ ), .B(\us02\/_0010_ ), .X(_0675_ ) );
sky130_fd_sc_hd__xor2_1 _2261_ ( .A(\us20\/_0011_ ), .B(\us31\/_0011_ ), .X(_0676_ ) );
sky130_fd_sc_hd__xnor3_1 _2262_ ( .A(_1419_ ), .B(\us13\/_0010_ ), .C(\us13\/_0011_ ), .X(_0677_ ) );
sky130_fd_sc_hd__xnor3_1 _2263_ ( .A(_0675_ ), .B(_0676_ ), .C(_0677_ ), .X(_0678_ ) );
sky130_fd_sc_hd__nand2_1 _2264_ ( .A(_0678_ ), .B(_0664_ ), .Y(_0679_ ) );
sky130_fd_sc_hd__nand2_1 _2265_ ( .A(\text_in_r\[59\] ), .B(_0550_ ), .Y(_0680_ ) );
sky130_fd_sc_hd__nand2_1 _2266_ ( .A(_0679_ ), .B(_0680_ ), .Y(_0681_ ) );
sky130_fd_sc_hd__xor2_1 _2267_ ( .A(\w2\[27\] ), .B(_0681_ ), .X(_1335_ ) );
sky130_fd_sc_hd__and2b_1 _2268_ ( .A_N(\text_in_r\[60\] ), .B(_0562_ ), .X(_0682_ ) );
sky130_fd_sc_hd__clkbuf_1 _2269_ ( .A(_0549_ ), .X(_0683_ ) );
sky130_fd_sc_hd__xnor2_1 _2270_ ( .A(\us02\/_0015_ ), .B(\us02\/_0011_ ), .Y(_0684_ ) );
sky130_fd_sc_hd__xnor2_1 _2271_ ( .A(\us20\/_0012_ ), .B(\us31\/_0012_ ), .Y(_0685_ ) );
sky130_fd_sc_hd__xnor3_1 _2272_ ( .A(_1419_ ), .B(\us13\/_0011_ ), .C(\us13\/_0012_ ), .X(_0686_ ) );
sky130_fd_sc_hd__xnor3_1 _2273_ ( .A(_0684_ ), .B(_0685_ ), .C(_0686_ ), .X(_0687_ ) );
sky130_fd_sc_hd__nor2_1 _2274_ ( .A(_0683_ ), .B(_0687_ ), .Y(_0688_ ) );
sky130_fd_sc_hd__nor2_1 _2275_ ( .A(_0682_ ), .B(_0688_ ), .Y(_0689_ ) );
sky130_fd_sc_hd__xor2_1 _2276_ ( .A(\w2\[28\] ), .B(_0689_ ), .X(_1336_ ) );
sky130_fd_sc_hd__and2_0 _2277_ ( .A(\text_in_r\[61\] ), .B(ld_r ), .X(_0690_ ) );
sky130_fd_sc_hd__xnor2_1 _2278_ ( .A(\us13\/_0013_ ), .B(\us20\/_0013_ ), .Y(_0691_ ) );
sky130_fd_sc_hd__xnor2_1 _2279_ ( .A(\us13\/_0012_ ), .B(\us02\/_0012_ ), .Y(_0692_ ) );
sky130_fd_sc_hd__xnor3_1 _2280_ ( .A(\us31\/_0013_ ), .B(_0691_ ), .C(_0692_ ), .X(_0693_ ) );
sky130_fd_sc_hd__nor2_1 _2281_ ( .A(_0653_ ), .B(_0693_ ), .Y(_0694_ ) );
sky130_fd_sc_hd__nor2_1 _2282_ ( .A(_0690_ ), .B(_0694_ ), .Y(_0695_ ) );
sky130_fd_sc_hd__xnor2_1 _2283_ ( .A(\w2\[29\] ), .B(_0695_ ), .Y(_1337_ ) );
sky130_fd_sc_hd__and2_0 _2284_ ( .A(\text_in_r\[62\] ), .B(ld_r ), .X(_0696_ ) );
sky130_fd_sc_hd__xor2_1 _2285_ ( .A(\us13\/_0013_ ), .B(\us02\/_0013_ ), .X(_0697_ ) );
sky130_fd_sc_hd__xor2_1 _2286_ ( .A(\us13\/_0014_ ), .B(\us31\/_0014_ ), .X(_0698_ ) );
sky130_fd_sc_hd__xnor3_1 _2287_ ( .A(\us20\/_0014_ ), .B(_0697_ ), .C(_0698_ ), .X(_0699_ ) );
sky130_fd_sc_hd__nor2_1 _2288_ ( .A(_0653_ ), .B(_0699_ ), .Y(_0700_ ) );
sky130_fd_sc_hd__nor2_1 _2289_ ( .A(_0696_ ), .B(_0700_ ), .Y(_0701_ ) );
sky130_fd_sc_hd__xnor2_1 _2290_ ( .A(\w2\[30\] ), .B(_0701_ ), .Y(_1338_ ) );
sky130_fd_sc_hd__and2_0 _2291_ ( .A(\text_in_r\[63\] ), .B(ld_r ), .X(_0702_ ) );
sky130_fd_sc_hd__xnor2_1 _2293_ ( .A(\us13\/_0014_ ), .B(\us31\/_0015_ ), .Y(_0704_ ) );
sky130_fd_sc_hd__xnor2_1 _2294_ ( .A(\us02\/_0014_ ), .B(_1451_ ), .Y(_0705_ ) );
sky130_fd_sc_hd__xnor3_1 _2295_ ( .A(_1419_ ), .B(_0704_ ), .C(_0705_ ), .X(_0706_ ) );
sky130_fd_sc_hd__nor2_1 _2296_ ( .A(_0653_ ), .B(_0706_ ), .Y(_0707_ ) );
sky130_fd_sc_hd__nor2_1 _2297_ ( .A(_0702_ ), .B(_0707_ ), .Y(_0708_ ) );
sky130_fd_sc_hd__xnor2_1 _2298_ ( .A(\w2\[31\] ), .B(_0708_ ), .Y(_1339_ ) );
sky130_fd_sc_hd__clkbuf_1 _2299_ ( .A(_0536_ ), .X(_0709_ ) );
sky130_fd_sc_hd__and2_0 _2300_ ( .A(\text_in_r\[24\] ), .B(_0709_ ), .X(_0710_ ) );
sky130_fd_sc_hd__inv_1 _2301_ ( .A(\us03\/_0015_ ), .Y(_0711_ ) );
sky130_fd_sc_hd__xnor2_1 _2302_ ( .A(\us10\/_0008_ ), .B(\us21\/_0008_ ), .Y(_0712_ ) );
sky130_fd_sc_hd__xor2_1 _2303_ ( .A(_1387_ ), .B(\us32\/_0008_ ), .X(_0713_ ) );
sky130_fd_sc_hd__xnor3_1 _2304_ ( .A(_0711_ ), .B(_0712_ ), .C(_0713_ ), .X(_0714_ ) );
sky130_fd_sc_hd__nor2_1 _2305_ ( .A(_0653_ ), .B(_0714_ ), .Y(_0715_ ) );
sky130_fd_sc_hd__nor2_1 _2306_ ( .A(_0710_ ), .B(_0715_ ), .Y(_0716_ ) );
sky130_fd_sc_hd__xnor2_1 _2307_ ( .A(\w3\[24\] ), .B(_0716_ ), .Y(_1348_ ) );
sky130_fd_sc_hd__and2b_1 _2308_ ( .A_N(\text_in_r\[25\] ), .B(_0562_ ), .X(_0717_ ) );
sky130_fd_sc_hd__xor2_1 _2309_ ( .A(\us03\/_0015_ ), .B(\us03\/_0008_ ), .X(_0718_ ) );
sky130_fd_sc_hd__xor2_1 _2310_ ( .A(\us21\/_0009_ ), .B(\us32\/_0009_ ), .X(_0719_ ) );
sky130_fd_sc_hd__xnor3_1 _2311_ ( .A(_1387_ ), .B(\us10\/_0008_ ), .C(\us10\/_0009_ ), .X(_0720_ ) );
sky130_fd_sc_hd__xnor3_1 _2312_ ( .A(_0718_ ), .B(_0719_ ), .C(_0720_ ), .X(_0721_ ) );
sky130_fd_sc_hd__nor2_1 _2313_ ( .A(_0683_ ), .B(_0721_ ), .Y(_0722_ ) );
sky130_fd_sc_hd__nor2_1 _2314_ ( .A(_0717_ ), .B(_0722_ ), .Y(_0723_ ) );
sky130_fd_sc_hd__xor2_1 _2315_ ( .A(\w3\[25\] ), .B(_0723_ ), .X(_1349_ ) );
sky130_fd_sc_hd__inv_1 _2316_ ( .A(\us21\/_0010_ ), .Y(_0724_ ) );
sky130_fd_sc_hd__xnor2_1 _2317_ ( .A(\us10\/_0009_ ), .B(\us03\/_0009_ ), .Y(_0725_ ) );
sky130_fd_sc_hd__xor2_1 _2318_ ( .A(\us10\/_0010_ ), .B(\us32\/_0010_ ), .X(_0726_ ) );
sky130_fd_sc_hd__xnor3_1 _2319_ ( .A(_0724_ ), .B(_0725_ ), .C(_0726_ ), .X(_0727_ ) );
sky130_fd_sc_hd__nand2_1 _2320_ ( .A(_0727_ ), .B(_0538_ ), .Y(_0728_ ) );
sky130_fd_sc_hd__or2b_1 _2321_ ( .A(\text_in_r\[26\] ), .B_N(_0911_ ), .X(_0729_ ) );
sky130_fd_sc_hd__nand2_1 _2322_ ( .A(_0728_ ), .B(_0729_ ), .Y(_0730_ ) );
sky130_fd_sc_hd__xnor2_1 _2323_ ( .A(\w3\[26\] ), .B(_0730_ ), .Y(_1350_ ) );
sky130_fd_sc_hd__and2b_1 _2324_ ( .A_N(\text_in_r\[27\] ), .B(_0562_ ), .X(_0731_ ) );
sky130_fd_sc_hd__xor2_1 _2325_ ( .A(\us03\/_0015_ ), .B(\us03\/_0010_ ), .X(_0732_ ) );
sky130_fd_sc_hd__xor2_1 _2326_ ( .A(\us21\/_0011_ ), .B(\us32\/_0011_ ), .X(_0733_ ) );
sky130_fd_sc_hd__xnor3_1 _2327_ ( .A(_1387_ ), .B(\us10\/_0010_ ), .C(\us10\/_0011_ ), .X(_0734_ ) );
sky130_fd_sc_hd__xnor3_1 _2328_ ( .A(_0732_ ), .B(_0733_ ), .C(_0734_ ), .X(_0735_ ) );
sky130_fd_sc_hd__nor2_1 _2329_ ( .A(_0683_ ), .B(_0735_ ), .Y(_0736_ ) );
sky130_fd_sc_hd__nor2_1 _2330_ ( .A(_0731_ ), .B(_0736_ ), .Y(_0737_ ) );
sky130_fd_sc_hd__xor2_1 _2331_ ( .A(\w3\[27\] ), .B(_0737_ ), .X(_1351_ ) );
sky130_fd_sc_hd__xnor2_1 _2332_ ( .A(\us03\/_0015_ ), .B(\us03\/_0011_ ), .Y(_0738_ ) );
sky130_fd_sc_hd__xnor2_1 _2333_ ( .A(\us21\/_0012_ ), .B(\us32\/_0012_ ), .Y(_0739_ ) );
sky130_fd_sc_hd__xnor3_1 _2334_ ( .A(_1387_ ), .B(\us10\/_0011_ ), .C(\us10\/_0012_ ), .X(_0740_ ) );
sky130_fd_sc_hd__xnor3_1 _2335_ ( .A(_0738_ ), .B(_0739_ ), .C(_0740_ ), .X(_0741_ ) );
sky130_fd_sc_hd__nand2_1 _2336_ ( .A(_0741_ ), .B(_0664_ ), .Y(_0742_ ) );
sky130_fd_sc_hd__nand2_1 _2337_ ( .A(\text_in_r\[28\] ), .B(_0550_ ), .Y(_0743_ ) );
sky130_fd_sc_hd__nand2_1 _2338_ ( .A(_0742_ ), .B(_0743_ ), .Y(_0744_ ) );
sky130_fd_sc_hd__xor2_1 _2339_ ( .A(\w3\[28\] ), .B(_0744_ ), .X(_1352_ ) );
sky130_fd_sc_hd__and2_0 _2340_ ( .A(\text_in_r\[29\] ), .B(_0709_ ), .X(_0745_ ) );
sky130_fd_sc_hd__xnor2_1 _2341_ ( .A(\us10\/_0013_ ), .B(\us21\/_0013_ ), .Y(_0746_ ) );
sky130_fd_sc_hd__xnor2_1 _2342_ ( .A(\us10\/_0012_ ), .B(\us03\/_0012_ ), .Y(_0747_ ) );
sky130_fd_sc_hd__xnor3_1 _2343_ ( .A(\us32\/_0013_ ), .B(_0746_ ), .C(_0747_ ), .X(_0748_ ) );
sky130_fd_sc_hd__nor2_1 _2344_ ( .A(_0653_ ), .B(_0748_ ), .Y(_0749_ ) );
sky130_fd_sc_hd__nor2_1 _2345_ ( .A(_0745_ ), .B(_0749_ ), .Y(_0750_ ) );
sky130_fd_sc_hd__xnor2_1 _2346_ ( .A(\w3\[29\] ), .B(_0750_ ), .Y(_1353_ ) );
sky130_fd_sc_hd__xor2_1 _2347_ ( .A(\us10\/_0013_ ), .B(\us03\/_0013_ ), .X(_0751_ ) );
sky130_fd_sc_hd__xor2_1 _2348_ ( .A(\us10\/_0014_ ), .B(\us32\/_0014_ ), .X(_0752_ ) );
sky130_fd_sc_hd__xnor3_1 _2349_ ( .A(\us21\/_0014_ ), .B(_0751_ ), .C(_0752_ ), .X(_0753_ ) );
sky130_fd_sc_hd__nand2_1 _2350_ ( .A(_0753_ ), .B(_0538_ ), .Y(_0754_ ) );
sky130_fd_sc_hd__or2b_1 _2351_ ( .A(\text_in_r\[30\] ), .B_N(_0911_ ), .X(_0755_ ) );
sky130_fd_sc_hd__nand2_1 _2352_ ( .A(_0754_ ), .B(_0755_ ), .Y(_0756_ ) );
sky130_fd_sc_hd__xnor2_1 _2353_ ( .A(\w3\[30\] ), .B(_0756_ ), .Y(_1354_ ) );
sky130_fd_sc_hd__xnor2_1 _2355_ ( .A(\us10\/_0014_ ), .B(\us32\/_0015_ ), .Y(_0758_ ) );
sky130_fd_sc_hd__xnor2_1 _2356_ ( .A(\us03\/_0014_ ), .B(\us21\/_0015_ ), .Y(_0759_ ) );
sky130_fd_sc_hd__xnor3_1 _2357_ ( .A(_1387_ ), .B(_0758_ ), .C(_0759_ ), .X(_0760_ ) );
sky130_fd_sc_hd__nand2_1 _2358_ ( .A(_0760_ ), .B(_0538_ ), .Y(_0761_ ) );
sky130_fd_sc_hd__or2b_1 _2359_ ( .A(\text_in_r\[31\] ), .B_N(_0911_ ), .X(_0762_ ) );
sky130_fd_sc_hd__nand2_1 _2360_ ( .A(_0761_ ), .B(_0762_ ), .Y(_0763_ ) );
sky130_fd_sc_hd__xnor2_1 _2361_ ( .A(\u0\/_0842_ ), .B(_0763_ ), .Y(_1355_ ) );
sky130_fd_sc_hd__and2_0 _2362_ ( .A(\text_in_r\[112\] ), .B(_0709_ ), .X(_0764_ ) );
sky130_fd_sc_hd__xnor2_1 _2363_ ( .A(\us22\/_0008_ ), .B(\us22\/_0015_ ), .Y(_0765_ ) );
sky130_fd_sc_hd__xor3_1 _2364_ ( .A(\us00\/_0008_ ), .B(_0765_ ), .C(_0534_ ), .X(_0766_ ) );
sky130_fd_sc_hd__nor2_1 _2365_ ( .A(_0653_ ), .B(_0766_ ), .Y(_0767_ ) );
sky130_fd_sc_hd__nor2_1 _2366_ ( .A(_0764_ ), .B(_0767_ ), .Y(_0768_ ) );
sky130_fd_sc_hd__xnor2_1 _2367_ ( .A(\w0\[16\] ), .B(_0768_ ), .Y(_1364_ ) );
sky130_fd_sc_hd__and2b_1 _2368_ ( .A_N(\text_in_r\[113\] ), .B(_0562_ ), .X(_0769_ ) );
sky130_fd_sc_hd__xnor2_1 _2369_ ( .A(_1379_ ), .B(\us11\/_0008_ ), .Y(_0770_ ) );
sky130_fd_sc_hd__xor2_1 _2370_ ( .A(\us00\/_0009_ ), .B(_0770_ ), .X(_0771_ ) );
sky130_fd_sc_hd__xor3_1 _2371_ ( .A(_0544_ ), .B(_0765_ ), .C(_0771_ ), .X(_0772_ ) );
sky130_fd_sc_hd__nor2_1 _2372_ ( .A(_0683_ ), .B(_0772_ ), .Y(_0773_ ) );
sky130_fd_sc_hd__nor2_1 _2373_ ( .A(_0769_ ), .B(_0773_ ), .Y(_0774_ ) );
sky130_fd_sc_hd__xor2_1 _2374_ ( .A(\w0\[17\] ), .B(_0774_ ), .X(_1365_ ) );
sky130_fd_sc_hd__xnor3_1 _2375_ ( .A(\us33\/_0010_ ), .B(\us00\/_0010_ ), .C(_0556_ ), .X(_0775_ ) );
sky130_fd_sc_hd__xor3_1 _2376_ ( .A(_1373_ ), .B(\us22\/_0009_ ), .C(_0775_ ), .X(_0776_ ) );
sky130_fd_sc_hd__nand2_1 _2377_ ( .A(_0776_ ), .B(_0664_ ), .Y(_0777_ ) );
sky130_fd_sc_hd__nand2_1 _2378_ ( .A(\text_in_r\[114\] ), .B(_0550_ ), .Y(_0778_ ) );
sky130_fd_sc_hd__nand2_1 _2379_ ( .A(_0777_ ), .B(_0778_ ), .Y(_0779_ ) );
sky130_fd_sc_hd__xor2_1 _2380_ ( .A(\w0\[18\] ), .B(_0779_ ), .X(_1366_ ) );
sky130_fd_sc_hd__clkbuf_1 _2381_ ( .A(ld_r ), .X(_0780_ ) );
sky130_fd_sc_hd__and2b_1 _2382_ ( .A_N(\text_in_r\[115\] ), .B(_0780_ ), .X(_0781_ ) );
sky130_fd_sc_hd__xor2_1 _2383_ ( .A(\us22\/_0010_ ), .B(\us22\/_0015_ ), .X(_0782_ ) );
sky130_fd_sc_hd__xnor2_1 _2384_ ( .A(_1379_ ), .B(\us11\/_0010_ ), .Y(_0783_ ) );
sky130_fd_sc_hd__xor2_1 _2385_ ( .A(\us00\/_0011_ ), .B(_0783_ ), .X(_0784_ ) );
sky130_fd_sc_hd__xnor3_1 _2386_ ( .A(_0566_ ), .B(_0782_ ), .C(_0784_ ), .X(_0785_ ) );
sky130_fd_sc_hd__nor2_1 _2387_ ( .A(_0683_ ), .B(_0785_ ), .Y(_0786_ ) );
sky130_fd_sc_hd__nor2_1 _2388_ ( .A(_0781_ ), .B(_0786_ ), .Y(_0787_ ) );
sky130_fd_sc_hd__xor2_1 _2389_ ( .A(\w0\[19\] ), .B(_0787_ ), .X(_1367_ ) );
sky130_fd_sc_hd__xnor2_1 _2390_ ( .A(\us22\/_0011_ ), .B(\us22\/_0015_ ), .Y(_0788_ ) );
sky130_fd_sc_hd__xnor2_1 _2391_ ( .A(_1379_ ), .B(\us11\/_0011_ ), .Y(_0789_ ) );
sky130_fd_sc_hd__xor2_1 _2392_ ( .A(\us00\/_0012_ ), .B(_0789_ ), .X(_0790_ ) );
sky130_fd_sc_hd__xnor3_1 _2393_ ( .A(_0573_ ), .B(_0788_ ), .C(_0790_ ), .X(_0791_ ) );
sky130_fd_sc_hd__nand2_1 _2394_ ( .A(_0791_ ), .B(_0664_ ), .Y(_0792_ ) );
sky130_fd_sc_hd__nand2_1 _2395_ ( .A(\text_in_r\[116\] ), .B(_0550_ ), .Y(_0793_ ) );
sky130_fd_sc_hd__nand2_1 _2396_ ( .A(_0792_ ), .B(_0793_ ), .Y(_0794_ ) );
sky130_fd_sc_hd__xor2_1 _2397_ ( .A(\w0\[20\] ), .B(_0794_ ), .X(_1368_ ) );
sky130_fd_sc_hd__inv_1 _2398_ ( .A(\us33\/_0013_ ), .Y(_0795_ ) );
sky130_fd_sc_hd__inv_1 _2399_ ( .A(\us22\/_0012_ ), .Y(_0796_ ) );
sky130_fd_sc_hd__xnor3_1 _2400_ ( .A(\us11\/_0012_ ), .B(\us00\/_0013_ ), .C(_0796_ ), .X(_0797_ ) );
sky130_fd_sc_hd__xor3_1 _2401_ ( .A(\us22\/_0013_ ), .B(_0795_ ), .C(_0797_ ), .X(_0798_ ) );
sky130_fd_sc_hd__nand2_1 _2402_ ( .A(_0798_ ), .B(_0538_ ), .Y(_0799_ ) );
sky130_fd_sc_hd__or2b_1 _2403_ ( .A(\text_in_r\[117\] ), .B_N(_0911_ ), .X(_0800_ ) );
sky130_fd_sc_hd__nand2_1 _2404_ ( .A(_0799_ ), .B(_0800_ ), .Y(_0801_ ) );
sky130_fd_sc_hd__xnor2_1 _2405_ ( .A(\w0\[21\] ), .B(_0801_ ), .Y(_1369_ ) );
sky130_fd_sc_hd__xnor2_1 _2406_ ( .A(\us22\/_0014_ ), .B(\us33\/_0014_ ), .Y(_0802_ ) );
sky130_fd_sc_hd__xnor3_1 _2407_ ( .A(\us00\/_0014_ ), .B(_0578_ ), .C(_0802_ ), .X(_0803_ ) );
sky130_fd_sc_hd__nand2_1 _2409_ ( .A(_0803_ ), .B(_1024_ ), .Y(_0805_ ) );
sky130_fd_sc_hd__or2b_1 _2410_ ( .A(\text_in_r\[118\] ), .B_N(_0911_ ), .X(_0806_ ) );
sky130_fd_sc_hd__nand2_1 _2411_ ( .A(_0805_ ), .B(_0806_ ), .Y(_0807_ ) );
sky130_fd_sc_hd__xnor2_1 _2412_ ( .A(\w0\[22\] ), .B(_0807_ ), .Y(_1370_ ) );
sky130_fd_sc_hd__and2_0 _2413_ ( .A(\text_in_r\[119\] ), .B(_0709_ ), .X(_0808_ ) );
sky130_fd_sc_hd__xnor3_1 _2414_ ( .A(\us22\/_0014_ ), .B(\us22\/_0015_ ), .C(\us33\/_0015_ ), .X(_0809_ ) );
sky130_fd_sc_hd__xor3_1 _2415_ ( .A(\us00\/_0015_ ), .B(\us11\/_0014_ ), .C(_0809_ ), .X(_0810_ ) );
sky130_fd_sc_hd__nor2_1 _2416_ ( .A(_0653_ ), .B(_0810_ ), .Y(_0811_ ) );
sky130_fd_sc_hd__nor2_1 _2417_ ( .A(_0808_ ), .B(_0811_ ), .Y(_0812_ ) );
sky130_fd_sc_hd__xnor2_1 _2418_ ( .A(\w0\[23\] ), .B(_0812_ ), .Y(_1371_ ) );
sky130_fd_sc_hd__xnor2_1 _2419_ ( .A(\us23\/_0008_ ), .B(\us23\/_0015_ ), .Y(_0813_ ) );
sky130_fd_sc_hd__xor3_1 _2420_ ( .A(\us01\/_0008_ ), .B(_0813_ ), .C(_0600_ ), .X(_0814_ ) );
sky130_fd_sc_hd__nand2_1 _2421_ ( .A(_0814_ ), .B(_1024_ ), .Y(_0815_ ) );
sky130_fd_sc_hd__or2b_1 _2422_ ( .A(\text_in_r\[80\] ), .B_N(_0911_ ), .X(_0816_ ) );
sky130_fd_sc_hd__nand2_1 _2423_ ( .A(_0815_ ), .B(_0816_ ), .Y(_0817_ ) );
sky130_fd_sc_hd__xnor2_1 _2424_ ( .A(\w1\[16\] ), .B(_0817_ ), .Y(_1388_ ) );
sky130_fd_sc_hd__and2b_1 _2425_ ( .A_N(\text_in_r\[81\] ), .B(_0780_ ), .X(_0818_ ) );
sky130_fd_sc_hd__xnor2_1 _2426_ ( .A(\us12\/_0015_ ), .B(\us12\/_0008_ ), .Y(_0819_ ) );
sky130_fd_sc_hd__xor2_1 _2427_ ( .A(\us01\/_0009_ ), .B(_0819_ ), .X(_0820_ ) );
sky130_fd_sc_hd__xor3_1 _2428_ ( .A(_0605_ ), .B(_0813_ ), .C(_0820_ ), .X(_0821_ ) );
sky130_fd_sc_hd__nor2_1 _2429_ ( .A(_0683_ ), .B(_0821_ ), .Y(_0822_ ) );
sky130_fd_sc_hd__nor2_1 _2430_ ( .A(_0818_ ), .B(_0822_ ), .Y(_0823_ ) );
sky130_fd_sc_hd__xor2_1 _2431_ ( .A(\w1\[17\] ), .B(_0823_ ), .X(_1389_ ) );
sky130_fd_sc_hd__xnor3_1 _2432_ ( .A(\us30\/_0010_ ), .B(\us01\/_0010_ ), .C(_0612_ ), .X(_0824_ ) );
sky130_fd_sc_hd__xor3_1 _2433_ ( .A(\us12\/_0009_ ), .B(\us23\/_0009_ ), .C(_0824_ ), .X(_0825_ ) );
sky130_fd_sc_hd__nand2_1 _2434_ ( .A(_0825_ ), .B(_0664_ ), .Y(_0826_ ) );
sky130_fd_sc_hd__nand2_1 _2435_ ( .A(\text_in_r\[82\] ), .B(_0550_ ), .Y(_0827_ ) );
sky130_fd_sc_hd__nand2_1 _2436_ ( .A(_0826_ ), .B(_0827_ ), .Y(_0828_ ) );
sky130_fd_sc_hd__xor2_1 _2437_ ( .A(\w1\[18\] ), .B(_0828_ ), .X(_1390_ ) );
sky130_fd_sc_hd__xor2_1 _2438_ ( .A(\us23\/_0010_ ), .B(\us23\/_0015_ ), .X(_0829_ ) );
sky130_fd_sc_hd__xnor2_1 _2439_ ( .A(\us12\/_0015_ ), .B(\us12\/_0010_ ), .Y(_0830_ ) );
sky130_fd_sc_hd__xor2_1 _2440_ ( .A(\us01\/_0011_ ), .B(_0830_ ), .X(_0831_ ) );
sky130_fd_sc_hd__xnor3_1 _2441_ ( .A(_0620_ ), .B(_0829_ ), .C(_0831_ ), .X(_0832_ ) );
sky130_fd_sc_hd__nand2_1 _2442_ ( .A(_0832_ ), .B(_0664_ ), .Y(_0833_ ) );
sky130_fd_sc_hd__nand2_1 _2443_ ( .A(\text_in_r\[83\] ), .B(_0550_ ), .Y(_0834_ ) );
sky130_fd_sc_hd__nand2_1 _2444_ ( .A(_0833_ ), .B(_0834_ ), .Y(_0835_ ) );
sky130_fd_sc_hd__xor2_1 _2445_ ( .A(\w1\[19\] ), .B(_0835_ ), .X(_1391_ ) );
sky130_fd_sc_hd__xnor2_1 _2446_ ( .A(\us23\/_0011_ ), .B(\us23\/_0015_ ), .Y(_0836_ ) );
sky130_fd_sc_hd__xnor2_1 _2447_ ( .A(\us12\/_0015_ ), .B(\us12\/_0011_ ), .Y(_0837_ ) );
sky130_fd_sc_hd__xor2_1 _2448_ ( .A(\us01\/_0012_ ), .B(_0837_ ), .X(_0838_ ) );
sky130_fd_sc_hd__xnor3_1 _2449_ ( .A(_0626_ ), .B(_0836_ ), .C(_0838_ ), .X(_0839_ ) );
sky130_fd_sc_hd__nand2_1 _2450_ ( .A(_0839_ ), .B(_0664_ ), .Y(_0840_ ) );
sky130_fd_sc_hd__buf_2 _2451_ ( .A(_0549_ ), .X(_0841_ ) );
sky130_fd_sc_hd__nand2_1 _2452_ ( .A(\text_in_r\[84\] ), .B(_0841_ ), .Y(_0842_ ) );
sky130_fd_sc_hd__nand2_1 _2453_ ( .A(_0840_ ), .B(_0842_ ), .Y(_0843_ ) );
sky130_fd_sc_hd__xor2_1 _2454_ ( .A(\w1\[20\] ), .B(_0843_ ), .X(_1392_ ) );
sky130_fd_sc_hd__and2_0 _2455_ ( .A(\text_in_r\[85\] ), .B(_0709_ ), .X(_0844_ ) );
sky130_fd_sc_hd__xor2_1 _2456_ ( .A(\us23\/_0013_ ), .B(\us30\/_0013_ ), .X(_0845_ ) );
sky130_fd_sc_hd__xor2_1 _2457_ ( .A(\us12\/_0012_ ), .B(\us23\/_0012_ ), .X(_0846_ ) );
sky130_fd_sc_hd__xnor3_1 _2458_ ( .A(\us01\/_0013_ ), .B(_0845_ ), .C(_0846_ ), .X(_0847_ ) );
sky130_fd_sc_hd__nor2_1 _2459_ ( .A(_0653_ ), .B(_0847_ ), .Y(_0848_ ) );
sky130_fd_sc_hd__nor2_1 _2460_ ( .A(_0844_ ), .B(_0848_ ), .Y(_0849_ ) );
sky130_fd_sc_hd__xnor2_1 _2461_ ( .A(\w1\[21\] ), .B(_0849_ ), .Y(_1393_ ) );
sky130_fd_sc_hd__xnor2_1 _2462_ ( .A(\us23\/_0014_ ), .B(\us30\/_0014_ ), .Y(_0850_ ) );
sky130_fd_sc_hd__xnor3_1 _2463_ ( .A(\us01\/_0014_ ), .B(_0632_ ), .C(_0850_ ), .X(_0851_ ) );
sky130_fd_sc_hd__nand2_1 _2464_ ( .A(_0851_ ), .B(_1024_ ), .Y(_0852_ ) );
sky130_fd_sc_hd__or2b_1 _2465_ ( .A(\text_in_r\[86\] ), .B_N(_0911_ ), .X(_0853_ ) );
sky130_fd_sc_hd__nand2_1 _2466_ ( .A(_0852_ ), .B(_0853_ ), .Y(_0854_ ) );
sky130_fd_sc_hd__xnor2_1 _2467_ ( .A(\w1\[22\] ), .B(_0854_ ), .Y(_1394_ ) );
sky130_fd_sc_hd__xnor3_1 _2468_ ( .A(\us23\/_0014_ ), .B(\us23\/_0015_ ), .C(_0646_ ), .X(_0855_ ) );
sky130_fd_sc_hd__xor3_1 _2469_ ( .A(_0598_ ), .B(\us12\/_0014_ ), .C(_0855_ ), .X(_0856_ ) );
sky130_fd_sc_hd__nand2_1 _2470_ ( .A(_0856_ ), .B(_0664_ ), .Y(_0857_ ) );
sky130_fd_sc_hd__nand2_1 _2471_ ( .A(\text_in_r\[87\] ), .B(_0841_ ), .Y(_0858_ ) );
sky130_fd_sc_hd__nand2_1 _2472_ ( .A(_0857_ ), .B(_0858_ ), .Y(_0859_ ) );
sky130_fd_sc_hd__xor2_1 _2473_ ( .A(\w1\[23\] ), .B(_0859_ ), .X(_1395_ ) );
sky130_fd_sc_hd__and2_0 _2474_ ( .A(\text_in_r\[48\] ), .B(_0709_ ), .X(_0860_ ) );
sky130_fd_sc_hd__xnor2_1 _2475_ ( .A(\us20\/_0008_ ), .B(_1451_ ), .Y(_0861_ ) );
sky130_fd_sc_hd__xor3_1 _2476_ ( .A(\us02\/_0008_ ), .B(_0861_ ), .C(_0656_ ), .X(_0862_ ) );
sky130_fd_sc_hd__nor2_1 _2477_ ( .A(_0653_ ), .B(_0862_ ), .Y(_0863_ ) );
sky130_fd_sc_hd__nor2_1 _2478_ ( .A(_0860_ ), .B(_0863_ ), .Y(_0864_ ) );
sky130_fd_sc_hd__xnor2_1 _2479_ ( .A(\w2\[16\] ), .B(_0864_ ), .Y(_1404_ ) );
sky130_fd_sc_hd__and2b_1 _2480_ ( .A_N(\text_in_r\[49\] ), .B(_0780_ ), .X(_0865_ ) );
sky130_fd_sc_hd__xnor2_1 _2481_ ( .A(_1419_ ), .B(\us13\/_0008_ ), .Y(_0866_ ) );
sky130_fd_sc_hd__xor2_1 _2482_ ( .A(\us02\/_0009_ ), .B(_0866_ ), .X(_0867_ ) );
sky130_fd_sc_hd__xor3_1 _2483_ ( .A(_0661_ ), .B(_0861_ ), .C(_0867_ ), .X(_0868_ ) );
sky130_fd_sc_hd__nor2_1 _2484_ ( .A(_0683_ ), .B(_0868_ ), .Y(_0869_ ) );
sky130_fd_sc_hd__nor2_1 _2485_ ( .A(_0865_ ), .B(_0869_ ), .Y(_0870_ ) );
sky130_fd_sc_hd__xor2_1 _2486_ ( .A(\w2\[17\] ), .B(_0870_ ), .X(_1405_ ) );
sky130_fd_sc_hd__xnor3_1 _2487_ ( .A(\us31\/_0010_ ), .B(\us02\/_0010_ ), .C(_0668_ ), .X(_0871_ ) );
sky130_fd_sc_hd__xor3_1 _2488_ ( .A(\us13\/_0009_ ), .B(\us20\/_0009_ ), .C(_0871_ ), .X(_0872_ ) );
sky130_fd_sc_hd__nand2_1 _2489_ ( .A(_0872_ ), .B(_0664_ ), .Y(_0873_ ) );
sky130_fd_sc_hd__nand2_1 _2490_ ( .A(\text_in_r\[50\] ), .B(_0841_ ), .Y(_0874_ ) );
sky130_fd_sc_hd__nand2_1 _2491_ ( .A(_0873_ ), .B(_0874_ ), .Y(_0875_ ) );
sky130_fd_sc_hd__xor2_1 _2492_ ( .A(\w2\[18\] ), .B(_0875_ ), .X(_1406_ ) );
sky130_fd_sc_hd__xor2_1 _2493_ ( .A(\us20\/_0010_ ), .B(_1451_ ), .X(_0876_ ) );
sky130_fd_sc_hd__xnor2_1 _2494_ ( .A(_1419_ ), .B(\us13\/_0010_ ), .Y(_0877_ ) );
sky130_fd_sc_hd__xor2_1 _2495_ ( .A(\us02\/_0011_ ), .B(_0877_ ), .X(_0878_ ) );
sky130_fd_sc_hd__xnor3_1 _2496_ ( .A(_0676_ ), .B(_0876_ ), .C(_0878_ ), .X(_0879_ ) );
sky130_fd_sc_hd__clkbuf_1 _2497_ ( .A(_0537_ ), .X(_0880_ ) );
sky130_fd_sc_hd__nand2_1 _2498_ ( .A(_0879_ ), .B(_0880_ ), .Y(_0881_ ) );
sky130_fd_sc_hd__nand2_1 _2499_ ( .A(\text_in_r\[51\] ), .B(_0841_ ), .Y(_0882_ ) );
sky130_fd_sc_hd__nand2_1 _2500_ ( .A(_0881_ ), .B(_0882_ ), .Y(_0883_ ) );
sky130_fd_sc_hd__xor2_1 _2501_ ( .A(\w2\[19\] ), .B(_0883_ ), .X(_1407_ ) );
sky130_fd_sc_hd__and2b_1 _2502_ ( .A_N(\text_in_r\[52\] ), .B(_0780_ ), .X(_0884_ ) );
sky130_fd_sc_hd__xnor2_1 _2503_ ( .A(\us20\/_0011_ ), .B(_1451_ ), .Y(_0885_ ) );
sky130_fd_sc_hd__xnor2_1 _2504_ ( .A(_1419_ ), .B(\us13\/_0011_ ), .Y(_0886_ ) );
sky130_fd_sc_hd__xor2_1 _2505_ ( .A(\us02\/_0012_ ), .B(_0886_ ), .X(_0887_ ) );
sky130_fd_sc_hd__xnor3_1 _2506_ ( .A(_0685_ ), .B(_0885_ ), .C(_0887_ ), .X(_0888_ ) );
sky130_fd_sc_hd__nor2_1 _2507_ ( .A(_0683_ ), .B(_0888_ ), .Y(_0889_ ) );
sky130_fd_sc_hd__nor2_1 _2508_ ( .A(_0884_ ), .B(_0889_ ), .Y(_0890_ ) );
sky130_fd_sc_hd__xor2_1 _2509_ ( .A(\w2\[20\] ), .B(_0890_ ), .X(_1408_ ) );
sky130_fd_sc_hd__xor2_1 _2510_ ( .A(\us20\/_0013_ ), .B(\us31\/_0013_ ), .X(_0891_ ) );
sky130_fd_sc_hd__xor2_1 _2511_ ( .A(\us13\/_0012_ ), .B(\us20\/_0012_ ), .X(_0892_ ) );
sky130_fd_sc_hd__xnor3_1 _2512_ ( .A(\us02\/_0013_ ), .B(_0891_ ), .C(_0892_ ), .X(_0893_ ) );
sky130_fd_sc_hd__nand2_1 _2513_ ( .A(_0893_ ), .B(_1024_ ), .Y(_0894_ ) );
sky130_fd_sc_hd__or2b_1 _2514_ ( .A(\text_in_r\[53\] ), .B_N(_0911_ ), .X(_0895_ ) );
sky130_fd_sc_hd__nand2_1 _2515_ ( .A(_0894_ ), .B(_0895_ ), .Y(_0896_ ) );
sky130_fd_sc_hd__xnor2_1 _2516_ ( .A(\w2\[21\] ), .B(_0896_ ), .Y(_1409_ ) );
sky130_fd_sc_hd__and2_0 _2517_ ( .A(\text_in_r\[54\] ), .B(_0709_ ), .X(_0897_ ) );
sky130_fd_sc_hd__clkbuf_1 _2518_ ( .A(_0549_ ), .X(_0898_ ) );
sky130_fd_sc_hd__xnor2_1 _2519_ ( .A(\us20\/_0014_ ), .B(\us31\/_0014_ ), .Y(_0899_ ) );
sky130_fd_sc_hd__xnor3_1 _2520_ ( .A(\us02\/_0014_ ), .B(_0691_ ), .C(_0899_ ), .X(_0900_ ) );
sky130_fd_sc_hd__nor2_1 _2521_ ( .A(_0898_ ), .B(_0900_ ), .Y(_0901_ ) );
sky130_fd_sc_hd__nor2_1 _2522_ ( .A(_0897_ ), .B(_0901_ ), .Y(_0902_ ) );
sky130_fd_sc_hd__xnor2_1 _2523_ ( .A(\w2\[22\] ), .B(_0902_ ), .Y(_1410_ ) );
sky130_fd_sc_hd__and2b_1 _2524_ ( .A_N(\text_in_r\[55\] ), .B(_0780_ ), .X(_0903_ ) );
sky130_fd_sc_hd__xnor3_1 _2525_ ( .A(\us20\/_0014_ ), .B(_1451_ ), .C(\us31\/_0015_ ), .X(_0904_ ) );
sky130_fd_sc_hd__xor3_1 _2526_ ( .A(_0654_ ), .B(\us13\/_0014_ ), .C(_0904_ ), .X(_0905_ ) );
sky130_fd_sc_hd__nor2_1 _2527_ ( .A(_0683_ ), .B(_0905_ ), .Y(_0906_ ) );
sky130_fd_sc_hd__nor2_1 _2528_ ( .A(_0903_ ), .B(_0906_ ), .Y(_0907_ ) );
sky130_fd_sc_hd__xor2_1 _2529_ ( .A(\w2\[23\] ), .B(_0907_ ), .X(_1411_ ) );
sky130_fd_sc_hd__xnor2_1 _2530_ ( .A(\us21\/_0008_ ), .B(\us21\/_0015_ ), .Y(_0908_ ) );
sky130_fd_sc_hd__xor3_1 _2531_ ( .A(\us03\/_0008_ ), .B(_0908_ ), .C(_0713_ ), .X(_0909_ ) );
sky130_fd_sc_hd__nand2_1 _2532_ ( .A(_0909_ ), .B(_1024_ ), .Y(_0910_ ) );
sky130_fd_sc_hd__buf_2 _2533_ ( .A(_0536_ ), .X(_0911_ ) );
sky130_fd_sc_hd__or2b_1 _2534_ ( .A(\text_in_r\[16\] ), .B_N(_0911_ ), .X(_0912_ ) );
sky130_fd_sc_hd__nand2_1 _2535_ ( .A(_0910_ ), .B(_0912_ ), .Y(_0913_ ) );
sky130_fd_sc_hd__xnor2_1 _2536_ ( .A(\w3\[16\] ), .B(_0913_ ), .Y(_1420_ ) );
sky130_fd_sc_hd__and2b_1 _2537_ ( .A_N(\text_in_r\[17\] ), .B(_0780_ ), .X(_0914_ ) );
sky130_fd_sc_hd__xnor2_1 _2538_ ( .A(_1387_ ), .B(\us10\/_0008_ ), .Y(_0915_ ) );
sky130_fd_sc_hd__xor2_1 _2539_ ( .A(\us03\/_0009_ ), .B(_0915_ ), .X(_0916_ ) );
sky130_fd_sc_hd__xor3_1 _2540_ ( .A(_0719_ ), .B(_0908_ ), .C(_0916_ ), .X(_0917_ ) );
sky130_fd_sc_hd__nor2_1 _2541_ ( .A(_0683_ ), .B(_0917_ ), .Y(_0918_ ) );
sky130_fd_sc_hd__nor2_1 _2542_ ( .A(_0914_ ), .B(_0918_ ), .Y(_0919_ ) );
sky130_fd_sc_hd__xor2_1 _2543_ ( .A(\w3\[17\] ), .B(_0919_ ), .X(_1421_ ) );
sky130_fd_sc_hd__and2b_1 _2544_ ( .A_N(\text_in_r\[18\] ), .B(_0780_ ), .X(_0920_ ) );
sky130_fd_sc_hd__clkbuf_1 _2545_ ( .A(_0549_ ), .X(_0921_ ) );
sky130_fd_sc_hd__xnor3_1 _2546_ ( .A(\us32\/_0010_ ), .B(\us03\/_0010_ ), .C(_0724_ ), .X(_0922_ ) );
sky130_fd_sc_hd__xor3_1 _2547_ ( .A(\us10\/_0009_ ), .B(\us21\/_0009_ ), .C(_0922_ ), .X(_0923_ ) );
sky130_fd_sc_hd__nor2_1 _2548_ ( .A(_0921_ ), .B(_0923_ ), .Y(_0924_ ) );
sky130_fd_sc_hd__nor2_1 _2549_ ( .A(_0920_ ), .B(_0924_ ), .Y(_0925_ ) );
sky130_fd_sc_hd__xor2_1 _2550_ ( .A(\w3\[18\] ), .B(_0925_ ), .X(_1422_ ) );
sky130_fd_sc_hd__xor2_1 _2551_ ( .A(\us21\/_0010_ ), .B(\us21\/_0015_ ), .X(_0926_ ) );
sky130_fd_sc_hd__xnor2_1 _2552_ ( .A(_1387_ ), .B(\us10\/_0010_ ), .Y(_0927_ ) );
sky130_fd_sc_hd__xor2_1 _2553_ ( .A(\us03\/_0011_ ), .B(_0927_ ), .X(_0928_ ) );
sky130_fd_sc_hd__xnor3_1 _2554_ ( .A(_0733_ ), .B(_0926_ ), .C(_0928_ ), .X(_0929_ ) );
sky130_fd_sc_hd__nand2_1 _2555_ ( .A(_0929_ ), .B(_0880_ ), .Y(_0930_ ) );
sky130_fd_sc_hd__nand2_1 _2556_ ( .A(\text_in_r\[19\] ), .B(_0841_ ), .Y(_0931_ ) );
sky130_fd_sc_hd__nand2_1 _2557_ ( .A(_0930_ ), .B(_0931_ ), .Y(_0932_ ) );
sky130_fd_sc_hd__xor2_1 _2558_ ( .A(\w3\[19\] ), .B(_0932_ ), .X(_1423_ ) );
sky130_fd_sc_hd__xnor2_1 _2559_ ( .A(\us21\/_0011_ ), .B(\us21\/_0015_ ), .Y(_0933_ ) );
sky130_fd_sc_hd__xnor2_1 _2560_ ( .A(_1387_ ), .B(\us10\/_0011_ ), .Y(_0934_ ) );
sky130_fd_sc_hd__xor2_1 _2561_ ( .A(\us03\/_0012_ ), .B(_0934_ ), .X(_0935_ ) );
sky130_fd_sc_hd__xnor3_1 _2562_ ( .A(_0739_ ), .B(_0933_ ), .C(_0935_ ), .X(_0936_ ) );
sky130_fd_sc_hd__nand2_1 _2563_ ( .A(_0936_ ), .B(_0880_ ), .Y(_0937_ ) );
sky130_fd_sc_hd__nand2_1 _2564_ ( .A(\text_in_r\[20\] ), .B(_0841_ ), .Y(_0938_ ) );
sky130_fd_sc_hd__nand2_1 _2565_ ( .A(_0937_ ), .B(_0938_ ), .Y(_0939_ ) );
sky130_fd_sc_hd__xor2_1 _2566_ ( .A(\w3\[20\] ), .B(_0939_ ), .X(_1424_ ) );
sky130_fd_sc_hd__xor2_1 _2567_ ( .A(\us21\/_0013_ ), .B(\us32\/_0013_ ), .X(_0940_ ) );
sky130_fd_sc_hd__xor2_1 _2568_ ( .A(\us10\/_0012_ ), .B(\us21\/_0012_ ), .X(_0941_ ) );
sky130_fd_sc_hd__xnor3_1 _2569_ ( .A(\us03\/_0013_ ), .B(_0940_ ), .C(_0941_ ), .X(_0942_ ) );
sky130_fd_sc_hd__nand2_1 _2570_ ( .A(_0942_ ), .B(_1024_ ), .Y(_0943_ ) );
sky130_fd_sc_hd__or2b_1 _2571_ ( .A(\text_in_r\[21\] ), .B_N(_0911_ ), .X(_0944_ ) );
sky130_fd_sc_hd__nand2_1 _2572_ ( .A(_0943_ ), .B(_0944_ ), .Y(_0945_ ) );
sky130_fd_sc_hd__xnor2_1 _2573_ ( .A(\w3\[21\] ), .B(_0945_ ), .Y(_1425_ ) );
sky130_fd_sc_hd__and2_0 _2574_ ( .A(\text_in_r\[22\] ), .B(_0709_ ), .X(_0946_ ) );
sky130_fd_sc_hd__xnor2_1 _2575_ ( .A(\us21\/_0014_ ), .B(\us32\/_0014_ ), .Y(_0947_ ) );
sky130_fd_sc_hd__xnor3_1 _2576_ ( .A(\us03\/_0014_ ), .B(_0746_ ), .C(_0947_ ), .X(_0948_ ) );
sky130_fd_sc_hd__nor2_1 _2577_ ( .A(_0898_ ), .B(_0948_ ), .Y(_0949_ ) );
sky130_fd_sc_hd__nor2_1 _2578_ ( .A(_0946_ ), .B(_0949_ ), .Y(_0950_ ) );
sky130_fd_sc_hd__xnor2_1 _2579_ ( .A(\w3\[22\] ), .B(_0950_ ), .Y(_1426_ ) );
sky130_fd_sc_hd__and2b_1 _2580_ ( .A_N(\text_in_r\[23\] ), .B(_0780_ ), .X(_0951_ ) );
sky130_fd_sc_hd__xnor3_1 _2581_ ( .A(\us21\/_0014_ ), .B(\us21\/_0015_ ), .C(\us32\/_0015_ ), .X(_0952_ ) );
sky130_fd_sc_hd__xor3_1 _2582_ ( .A(_0711_ ), .B(\us10\/_0014_ ), .C(_0952_ ), .X(_0953_ ) );
sky130_fd_sc_hd__nor2_1 _2583_ ( .A(_0921_ ), .B(_0953_ ), .Y(_0954_ ) );
sky130_fd_sc_hd__nor2_1 _2584_ ( .A(_0951_ ), .B(_0954_ ), .Y(_0955_ ) );
sky130_fd_sc_hd__xor2_1 _2585_ ( .A(\w3\[23\] ), .B(_0955_ ), .X(_1427_ ) );
sky130_fd_sc_hd__xor2_1 _2586_ ( .A(\us11\/_0008_ ), .B(\us00\/_0008_ ), .X(_0956_ ) );
sky130_fd_sc_hd__xor2_1 _2587_ ( .A(\us33\/_0008_ ), .B(\us33\/_0015_ ), .X(_0957_ ) );
sky130_fd_sc_hd__xnor3_1 _2588_ ( .A(\us22\/_0015_ ), .B(_0956_ ), .C(_0957_ ), .X(_0958_ ) );
sky130_fd_sc_hd__nand2_1 _2589_ ( .A(_0958_ ), .B(_1024_ ), .Y(_0959_ ) );
sky130_fd_sc_hd__or2b_1 _2590_ ( .A(\text_in_r\[104\] ), .B_N(_0911_ ), .X(_0960_ ) );
sky130_fd_sc_hd__nand2_1 _2591_ ( .A(_0959_ ), .B(_0960_ ), .Y(_0961_ ) );
sky130_fd_sc_hd__xnor2_1 _2592_ ( .A(\w0\[8\] ), .B(_0961_ ), .Y(_1428_ ) );
sky130_fd_sc_hd__xnor3_1 _2593_ ( .A(\us33\/_0008_ ), .B(\us33\/_0009_ ), .C(\us33\/_0015_ ), .X(_0962_ ) );
sky130_fd_sc_hd__xnor3_1 _2594_ ( .A(_0557_ ), .B(_0765_ ), .C(_0962_ ), .X(_0963_ ) );
sky130_fd_sc_hd__nand2_1 _2595_ ( .A(_0963_ ), .B(_0880_ ), .Y(_0964_ ) );
sky130_fd_sc_hd__nand2_1 _2596_ ( .A(\text_in_r\[105\] ), .B(_0841_ ), .Y(_0965_ ) );
sky130_fd_sc_hd__nand2_1 _2597_ ( .A(_0964_ ), .B(_0965_ ), .Y(_0966_ ) );
sky130_fd_sc_hd__xor2_1 _2598_ ( .A(\w0\[9\] ), .B(_0966_ ), .X(_1429_ ) );
sky130_fd_sc_hd__and2b_1 _2599_ ( .A_N(\text_in_r\[106\] ), .B(_0780_ ), .X(_0967_ ) );
sky130_fd_sc_hd__xor3_1 _2600_ ( .A(\us00\/_0010_ ), .B(_0544_ ), .C(_0558_ ), .X(_0968_ ) );
sky130_fd_sc_hd__nor2_1 _2601_ ( .A(_0921_ ), .B(_0968_ ), .Y(_0969_ ) );
sky130_fd_sc_hd__nor2_1 _2602_ ( .A(_0967_ ), .B(_0969_ ), .Y(_0970_ ) );
sky130_fd_sc_hd__xor2_1 _2603_ ( .A(\w0\[10\] ), .B(_0970_ ), .X(_1430_ ) );
sky130_fd_sc_hd__xor2_1 _2604_ ( .A(\us11\/_0011_ ), .B(\us00\/_0011_ ), .X(_0971_ ) );
sky130_fd_sc_hd__xnor3_1 _2605_ ( .A(\us33\/_0010_ ), .B(\us33\/_0011_ ), .C(\us33\/_0015_ ), .X(_0972_ ) );
sky130_fd_sc_hd__xnor3_1 _2606_ ( .A(_0782_ ), .B(_0971_ ), .C(_0972_ ), .X(_0973_ ) );
sky130_fd_sc_hd__nand2_1 _2607_ ( .A(_0973_ ), .B(_0880_ ), .Y(_0974_ ) );
sky130_fd_sc_hd__nand2_1 _2608_ ( .A(\text_in_r\[107\] ), .B(_0841_ ), .Y(_0975_ ) );
sky130_fd_sc_hd__nand2_1 _2609_ ( .A(_0974_ ), .B(_0975_ ), .Y(_0976_ ) );
sky130_fd_sc_hd__xor2_1 _2610_ ( .A(\w0\[11\] ), .B(_0976_ ), .X(_1431_ ) );
sky130_fd_sc_hd__xnor3_1 _2611_ ( .A(\us33\/_0011_ ), .B(\us33\/_0012_ ), .C(\us33\/_0015_ ), .X(_0977_ ) );
sky130_fd_sc_hd__xnor3_1 _2612_ ( .A(_0579_ ), .B(_0788_ ), .C(_0977_ ), .X(_0978_ ) );
sky130_fd_sc_hd__nand2_1 _2613_ ( .A(_0978_ ), .B(_0880_ ), .Y(_0979_ ) );
sky130_fd_sc_hd__nand2_1 _2614_ ( .A(\text_in_r\[108\] ), .B(_0841_ ), .Y(_0980_ ) );
sky130_fd_sc_hd__nand2_1 _2615_ ( .A(_0979_ ), .B(_0980_ ), .Y(_0981_ ) );
sky130_fd_sc_hd__xor2_1 _2616_ ( .A(\w0\[12\] ), .B(_0981_ ), .X(_1432_ ) );
sky130_fd_sc_hd__xnor3_1 _2617_ ( .A(_0795_ ), .B(_0573_ ), .C(_0585_ ), .X(_0982_ ) );
sky130_fd_sc_hd__nand2_1 _2618_ ( .A(_0982_ ), .B(_1024_ ), .Y(_0983_ ) );
sky130_fd_sc_hd__or2b_1 _2619_ ( .A(\text_in_r\[109\] ), .B_N(_0911_ ), .X(_0984_ ) );
sky130_fd_sc_hd__nand2_1 _2620_ ( .A(_0983_ ), .B(_0984_ ), .Y(_0985_ ) );
sky130_fd_sc_hd__xnor2_1 _2621_ ( .A(\w0\[13\] ), .B(_0985_ ), .Y(_1433_ ) );
sky130_fd_sc_hd__and2_0 _2622_ ( .A(\text_in_r\[110\] ), .B(_0709_ ), .X(_0986_ ) );
sky130_fd_sc_hd__xor2_1 _2623_ ( .A(\us22\/_0013_ ), .B(\us33\/_0013_ ), .X(_0987_ ) );
sky130_fd_sc_hd__xnor3_1 _2624_ ( .A(\us00\/_0014_ ), .B(_0586_ ), .C(_0987_ ), .X(_0988_ ) );
sky130_fd_sc_hd__nor2_1 _2625_ ( .A(_0898_ ), .B(_0988_ ), .Y(_0989_ ) );
sky130_fd_sc_hd__nor2_1 _2626_ ( .A(_0986_ ), .B(_0989_ ), .Y(_0990_ ) );
sky130_fd_sc_hd__xnor2_1 _2627_ ( .A(\w0\[14\] ), .B(_0990_ ), .Y(_1434_ ) );
sky130_fd_sc_hd__xor2_1 _2628_ ( .A(_1379_ ), .B(\us00\/_0015_ ), .X(_0991_ ) );
sky130_fd_sc_hd__xor3_1 _2629_ ( .A(\us33\/_0015_ ), .B(_0802_ ), .C(_0991_ ), .X(_0992_ ) );
sky130_fd_sc_hd__nand2_1 _2630_ ( .A(_0992_ ), .B(_1024_ ), .Y(_0993_ ) );
sky130_fd_sc_hd__or2b_1 _2631_ ( .A(\text_in_r\[111\] ), .B_N(_0911_ ), .X(_0994_ ) );
sky130_fd_sc_hd__nand2_1 _2632_ ( .A(_0993_ ), .B(_0994_ ), .Y(_0995_ ) );
sky130_fd_sc_hd__xnor2_1 _2633_ ( .A(\w0\[15\] ), .B(_0995_ ), .Y(_1435_ ) );
sky130_fd_sc_hd__xor2_1 _2634_ ( .A(\us12\/_0008_ ), .B(\us01\/_0008_ ), .X(_0996_ ) );
sky130_fd_sc_hd__xor2_1 _2635_ ( .A(\us30\/_0008_ ), .B(_0646_ ), .X(_0997_ ) );
sky130_fd_sc_hd__xnor3_1 _2636_ ( .A(\us23\/_0015_ ), .B(_0996_ ), .C(_0997_ ), .X(_0998_ ) );
sky130_fd_sc_hd__nand2_1 _2637_ ( .A(_0998_ ), .B(_1024_ ), .Y(_0999_ ) );
sky130_fd_sc_hd__or2b_1 _2638_ ( .A(\text_in_r\[72\] ), .B_N(_0911_ ), .X(_1000_ ) );
sky130_fd_sc_hd__nand2_1 _2639_ ( .A(_0999_ ), .B(_1000_ ), .Y(_1001_ ) );
sky130_fd_sc_hd__xnor2_1 _2640_ ( .A(\w1\[8\] ), .B(_1001_ ), .Y(_1452_ ) );
sky130_fd_sc_hd__xnor3_1 _2641_ ( .A(\us30\/_0008_ ), .B(\us30\/_0009_ ), .C(_0646_ ), .X(_1002_ ) );
sky130_fd_sc_hd__xnor3_1 _2642_ ( .A(_0613_ ), .B(_0813_ ), .C(_1002_ ), .X(_1003_ ) );
sky130_fd_sc_hd__nand2_1 _2643_ ( .A(_1003_ ), .B(_0880_ ), .Y(_1004_ ) );
sky130_fd_sc_hd__nand2_1 _2644_ ( .A(\text_in_r\[73\] ), .B(_0841_ ), .Y(_1005_ ) );
sky130_fd_sc_hd__nand2_1 _2645_ ( .A(_1004_ ), .B(_1005_ ), .Y(_1006_ ) );
sky130_fd_sc_hd__xor2_1 _2646_ ( .A(\w1\[9\] ), .B(_1006_ ), .X(_1453_ ) );
sky130_fd_sc_hd__xor3_1 _2647_ ( .A(\us01\/_0010_ ), .B(_0605_ ), .C(_0614_ ), .X(_1007_ ) );
sky130_fd_sc_hd__nand2_1 _2648_ ( .A(_1007_ ), .B(_0880_ ), .Y(_1008_ ) );
sky130_fd_sc_hd__buf_2 _2649_ ( .A(_0549_ ), .X(_1009_ ) );
sky130_fd_sc_hd__nand2_1 _2650_ ( .A(\text_in_r\[74\] ), .B(_1009_ ), .Y(_1010_ ) );
sky130_fd_sc_hd__nand2_1 _2651_ ( .A(_1008_ ), .B(_1010_ ), .Y(_1011_ ) );
sky130_fd_sc_hd__xor2_1 _2652_ ( .A(\w1\[10\] ), .B(_1011_ ), .X(_1454_ ) );
sky130_fd_sc_hd__xor2_1 _2653_ ( .A(\us12\/_0011_ ), .B(\us01\/_0011_ ), .X(_1012_ ) );
sky130_fd_sc_hd__xnor3_1 _2654_ ( .A(\us30\/_0010_ ), .B(\us30\/_0011_ ), .C(_0646_ ), .X(_1013_ ) );
sky130_fd_sc_hd__xnor3_1 _2655_ ( .A(_0829_ ), .B(_1012_ ), .C(_1013_ ), .X(_1014_ ) );
sky130_fd_sc_hd__nand2_1 _2656_ ( .A(_1014_ ), .B(_0880_ ), .Y(_1015_ ) );
sky130_fd_sc_hd__nand2_1 _2657_ ( .A(\text_in_r\[75\] ), .B(_1009_ ), .Y(_1016_ ) );
sky130_fd_sc_hd__nand2_1 _2658_ ( .A(_1015_ ), .B(_1016_ ), .Y(_1017_ ) );
sky130_fd_sc_hd__xor2_1 _2659_ ( .A(\w1\[11\] ), .B(_1017_ ), .X(_1455_ ) );
sky130_fd_sc_hd__and2b_1 _2660_ ( .A_N(\text_in_r\[76\] ), .B(_0780_ ), .X(_1018_ ) );
sky130_fd_sc_hd__xnor3_1 _2661_ ( .A(\us30\/_0011_ ), .B(\us30\/_0012_ ), .C(\us30\/_0015_ ), .X(_1019_ ) );
sky130_fd_sc_hd__xnor3_1 _2662_ ( .A(_0633_ ), .B(_0836_ ), .C(_1019_ ), .X(_1020_ ) );
sky130_fd_sc_hd__nor2_1 _2663_ ( .A(_0921_ ), .B(_1020_ ), .Y(_1021_ ) );
sky130_fd_sc_hd__nor2_1 _2664_ ( .A(_1018_ ), .B(_1021_ ), .Y(_1022_ ) );
sky130_fd_sc_hd__xor2_1 _2665_ ( .A(\w1\[12\] ), .B(_1022_ ), .X(_1456_ ) );
sky130_fd_sc_hd__xor3_1 _2666_ ( .A(\us30\/_0013_ ), .B(_0626_ ), .C(_0638_ ), .X(_1023_ ) );
sky130_fd_sc_hd__buf_2 _2667_ ( .A(_0537_ ), .X(_1024_ ) );
sky130_fd_sc_hd__nand2_1 _2668_ ( .A(_1023_ ), .B(_1024_ ), .Y(_1025_ ) );
sky130_fd_sc_hd__or2b_1 _2669_ ( .A(\text_in_r\[77\] ), .B_N(_0911_ ), .X(_1026_ ) );
sky130_fd_sc_hd__nand2_1 _2670_ ( .A(_1025_ ), .B(_1026_ ), .Y(_1027_ ) );
sky130_fd_sc_hd__xnor2_1 _2671_ ( .A(\w1\[13\] ), .B(_1027_ ), .Y(_1457_ ) );
sky130_fd_sc_hd__xnor3_1 _2672_ ( .A(\us01\/_0014_ ), .B(_0639_ ), .C(_0845_ ), .X(_1028_ ) );
sky130_fd_sc_hd__nand2_1 _2673_ ( .A(_1028_ ), .B(_1024_ ), .Y(_1029_ ) );
sky130_fd_sc_hd__or2b_1 _2674_ ( .A(\text_in_r\[78\] ), .B_N(_0911_ ), .X(_1030_ ) );
sky130_fd_sc_hd__nand2_1 _2675_ ( .A(_1029_ ), .B(_1030_ ), .Y(_1031_ ) );
sky130_fd_sc_hd__xnor2_1 _2676_ ( .A(\w1\[14\] ), .B(_1031_ ), .Y(_1458_ ) );
sky130_fd_sc_hd__xor2_1 _2677_ ( .A(\us12\/_0015_ ), .B(\us01\/_0015_ ), .X(_1032_ ) );
sky130_fd_sc_hd__xor3_1 _2678_ ( .A(_0646_ ), .B(_0850_ ), .C(_1032_ ), .X(_1033_ ) );
sky130_fd_sc_hd__nand2_1 _2679_ ( .A(_1033_ ), .B(_1024_ ), .Y(_1034_ ) );
sky130_fd_sc_hd__or2b_1 _2680_ ( .A(\text_in_r\[79\] ), .B_N(_0911_ ), .X(_1035_ ) );
sky130_fd_sc_hd__nand2_1 _2681_ ( .A(_1034_ ), .B(_1035_ ), .Y(_1036_ ) );
sky130_fd_sc_hd__xnor2_1 _2682_ ( .A(\w1\[15\] ), .B(_1036_ ), .Y(_1459_ ) );
sky130_fd_sc_hd__and2_0 _2683_ ( .A(\text_in_r\[40\] ), .B(_0709_ ), .X(_1037_ ) );
sky130_fd_sc_hd__xor2_1 _2684_ ( .A(\us13\/_0008_ ), .B(\us02\/_0008_ ), .X(_1038_ ) );
sky130_fd_sc_hd__xor2_1 _2685_ ( .A(\us31\/_0008_ ), .B(\us31\/_0015_ ), .X(_1039_ ) );
sky130_fd_sc_hd__xnor3_1 _2686_ ( .A(_1451_ ), .B(_1038_ ), .C(_1039_ ), .X(_1040_ ) );
sky130_fd_sc_hd__nor2_1 _2687_ ( .A(_0898_ ), .B(_1040_ ), .Y(_1041_ ) );
sky130_fd_sc_hd__nor2_1 _2688_ ( .A(_1037_ ), .B(_1041_ ), .Y(_1042_ ) );
sky130_fd_sc_hd__xnor2_1 _2689_ ( .A(\w2\[8\] ), .B(_1042_ ), .Y(_1476_ ) );
sky130_fd_sc_hd__and2b_1 _2690_ ( .A_N(\text_in_r\[41\] ), .B(_0549_ ), .X(_1043_ ) );
sky130_fd_sc_hd__xnor3_1 _2691_ ( .A(\us31\/_0008_ ), .B(\us31\/_0009_ ), .C(\us31\/_0015_ ), .X(_1044_ ) );
sky130_fd_sc_hd__xnor3_1 _2692_ ( .A(_0669_ ), .B(_0861_ ), .C(_1044_ ), .X(_1045_ ) );
sky130_fd_sc_hd__nor2_1 _2693_ ( .A(_0921_ ), .B(_1045_ ), .Y(_1046_ ) );
sky130_fd_sc_hd__nor2_1 _2694_ ( .A(_1043_ ), .B(_1046_ ), .Y(_1047_ ) );
sky130_fd_sc_hd__xor2_1 _2695_ ( .A(\w2\[9\] ), .B(_1047_ ), .X(_1477_ ) );
sky130_fd_sc_hd__xor3_1 _2696_ ( .A(\us02\/_0010_ ), .B(_0661_ ), .C(_0670_ ), .X(_1048_ ) );
sky130_fd_sc_hd__nand2_1 _2697_ ( .A(_1048_ ), .B(_0880_ ), .Y(_1049_ ) );
sky130_fd_sc_hd__nand2_1 _2698_ ( .A(\text_in_r\[42\] ), .B(_1009_ ), .Y(_1050_ ) );
sky130_fd_sc_hd__nand2_1 _2699_ ( .A(_1049_ ), .B(_1050_ ), .Y(_1051_ ) );
sky130_fd_sc_hd__xor2_1 _2700_ ( .A(\w2\[10\] ), .B(_1051_ ), .X(_1478_ ) );
sky130_fd_sc_hd__and2b_1 _2701_ ( .A_N(\text_in_r\[43\] ), .B(_0549_ ), .X(_1052_ ) );
sky130_fd_sc_hd__xor2_1 _2702_ ( .A(\us13\/_0011_ ), .B(\us02\/_0011_ ), .X(_1053_ ) );
sky130_fd_sc_hd__xnor3_1 _2703_ ( .A(\us31\/_0010_ ), .B(\us31\/_0011_ ), .C(\us31\/_0015_ ), .X(_1054_ ) );
sky130_fd_sc_hd__xnor3_1 _2704_ ( .A(_0876_ ), .B(_1053_ ), .C(_1054_ ), .X(_1055_ ) );
sky130_fd_sc_hd__nor2_1 _2705_ ( .A(_0921_ ), .B(_1055_ ), .Y(_1056_ ) );
sky130_fd_sc_hd__nor2_1 _2706_ ( .A(_1052_ ), .B(_1056_ ), .Y(_1057_ ) );
sky130_fd_sc_hd__xor2_1 _2707_ ( .A(\w2\[11\] ), .B(_1057_ ), .X(_1479_ ) );
sky130_fd_sc_hd__and2b_1 _2708_ ( .A_N(\text_in_r\[44\] ), .B(_0549_ ), .X(_1058_ ) );
sky130_fd_sc_hd__xnor3_1 _2709_ ( .A(\us31\/_0011_ ), .B(\us31\/_0012_ ), .C(\us31\/_0015_ ), .X(_1059_ ) );
sky130_fd_sc_hd__xnor3_1 _2710_ ( .A(_0692_ ), .B(_0885_ ), .C(_1059_ ), .X(_1060_ ) );
sky130_fd_sc_hd__nor2_1 _2711_ ( .A(_0921_ ), .B(_1060_ ), .Y(_1061_ ) );
sky130_fd_sc_hd__nor2_1 _2712_ ( .A(_1058_ ), .B(_1061_ ), .Y(_1062_ ) );
sky130_fd_sc_hd__xor2_1 _2713_ ( .A(\w2\[12\] ), .B(_1062_ ), .X(_1480_ ) );
sky130_fd_sc_hd__xor3_1 _2714_ ( .A(\us31\/_0013_ ), .B(_0685_ ), .C(_0697_ ), .X(_1063_ ) );
sky130_fd_sc_hd__nand2_1 _2715_ ( .A(_1063_ ), .B(_1024_ ), .Y(_1064_ ) );
sky130_fd_sc_hd__or2b_1 _2716_ ( .A(\text_in_r\[45\] ), .B_N(_0911_ ), .X(_1065_ ) );
sky130_fd_sc_hd__nand2_1 _2717_ ( .A(_1064_ ), .B(_1065_ ), .Y(_1066_ ) );
sky130_fd_sc_hd__xnor2_1 _2718_ ( .A(\w2\[13\] ), .B(_1066_ ), .Y(_1481_ ) );
sky130_fd_sc_hd__xnor3_1 _2719_ ( .A(\us02\/_0014_ ), .B(_0698_ ), .C(_0891_ ), .X(_1067_ ) );
sky130_fd_sc_hd__nand2_1 _2720_ ( .A(_1067_ ), .B(_1024_ ), .Y(_1068_ ) );
sky130_fd_sc_hd__clkbuf_1 _2721_ ( .A(ld_r ), .X(_1069_ ) );
sky130_fd_sc_hd__or2b_1 _2722_ ( .A(\text_in_r\[46\] ), .B_N(_1069_ ), .X(_1070_ ) );
sky130_fd_sc_hd__nand2_1 _2723_ ( .A(_1068_ ), .B(_1070_ ), .Y(_1071_ ) );
sky130_fd_sc_hd__xnor2_1 _2724_ ( .A(\w2\[14\] ), .B(_1071_ ), .Y(_1482_ ) );
sky130_fd_sc_hd__xor2_1 _2725_ ( .A(_1419_ ), .B(\us02\/_0015_ ), .X(_1072_ ) );
sky130_fd_sc_hd__xor3_1 _2726_ ( .A(\us31\/_0015_ ), .B(_0899_ ), .C(_1072_ ), .X(_1073_ ) );
sky130_fd_sc_hd__nand2_1 _2727_ ( .A(_1073_ ), .B(_1024_ ), .Y(_1074_ ) );
sky130_fd_sc_hd__or2b_1 _2728_ ( .A(\text_in_r\[47\] ), .B_N(_1069_ ), .X(_1075_ ) );
sky130_fd_sc_hd__nand2_1 _2729_ ( .A(_1074_ ), .B(_1075_ ), .Y(_1076_ ) );
sky130_fd_sc_hd__xnor2_1 _2730_ ( .A(\w2\[15\] ), .B(_1076_ ), .Y(_1483_ ) );
sky130_fd_sc_hd__clkbuf_1 _2731_ ( .A(_0536_ ), .X(_1077_ ) );
sky130_fd_sc_hd__and2_0 _2732_ ( .A(\text_in_r\[8\] ), .B(_1077_ ), .X(_1078_ ) );
sky130_fd_sc_hd__xor2_1 _2733_ ( .A(\us10\/_0008_ ), .B(\us03\/_0008_ ), .X(_1079_ ) );
sky130_fd_sc_hd__xor2_1 _2734_ ( .A(\us32\/_0008_ ), .B(\us32\/_0015_ ), .X(_1080_ ) );
sky130_fd_sc_hd__xnor3_1 _2735_ ( .A(\us21\/_0015_ ), .B(_1079_ ), .C(_1080_ ), .X(_1081_ ) );
sky130_fd_sc_hd__nor2_1 _2736_ ( .A(_0898_ ), .B(_1081_ ), .Y(_1082_ ) );
sky130_fd_sc_hd__nor2_1 _2737_ ( .A(_1078_ ), .B(_1082_ ), .Y(_1083_ ) );
sky130_fd_sc_hd__xnor2_1 _2738_ ( .A(\w3\[8\] ), .B(_1083_ ), .Y(_1484_ ) );
sky130_fd_sc_hd__xnor3_1 _2739_ ( .A(\us32\/_0008_ ), .B(\us32\/_0009_ ), .C(\us32\/_0015_ ), .X(_1084_ ) );
sky130_fd_sc_hd__xnor3_1 _2740_ ( .A(_0725_ ), .B(_0908_ ), .C(_1084_ ), .X(_1085_ ) );
sky130_fd_sc_hd__clkbuf_1 _2741_ ( .A(_0537_ ), .X(_1086_ ) );
sky130_fd_sc_hd__nand2_1 _2742_ ( .A(_1085_ ), .B(_1086_ ), .Y(_1087_ ) );
sky130_fd_sc_hd__nand2_1 _2743_ ( .A(\text_in_r\[9\] ), .B(_1009_ ), .Y(_1088_ ) );
sky130_fd_sc_hd__nand2_1 _2744_ ( .A(_1087_ ), .B(_1088_ ), .Y(_1089_ ) );
sky130_fd_sc_hd__xor2_1 _2745_ ( .A(\w3\[9\] ), .B(_1089_ ), .X(_1485_ ) );
sky130_fd_sc_hd__xor3_1 _2746_ ( .A(\us03\/_0010_ ), .B(_0719_ ), .C(_0726_ ), .X(_1090_ ) );
sky130_fd_sc_hd__nand2_1 _2747_ ( .A(_1090_ ), .B(_1086_ ), .Y(_1091_ ) );
sky130_fd_sc_hd__nand2_1 _2748_ ( .A(\text_in_r\[10\] ), .B(_1009_ ), .Y(_1092_ ) );
sky130_fd_sc_hd__nand2_1 _2749_ ( .A(_1091_ ), .B(_1092_ ), .Y(_1093_ ) );
sky130_fd_sc_hd__xor2_1 _2750_ ( .A(\w3\[10\] ), .B(_1093_ ), .X(_1486_ ) );
sky130_fd_sc_hd__xor2_1 _2751_ ( .A(\us10\/_0011_ ), .B(\us03\/_0011_ ), .X(_1094_ ) );
sky130_fd_sc_hd__xnor3_1 _2752_ ( .A(\us32\/_0010_ ), .B(\us32\/_0011_ ), .C(\us32\/_0015_ ), .X(_1095_ ) );
sky130_fd_sc_hd__xnor3_1 _2753_ ( .A(_0926_ ), .B(_1094_ ), .C(_1095_ ), .X(_1096_ ) );
sky130_fd_sc_hd__nand2_1 _2754_ ( .A(_1096_ ), .B(_1086_ ), .Y(_1097_ ) );
sky130_fd_sc_hd__nand2_1 _2755_ ( .A(\text_in_r\[11\] ), .B(_1009_ ), .Y(_1098_ ) );
sky130_fd_sc_hd__nand2_1 _2756_ ( .A(_1097_ ), .B(_1098_ ), .Y(_1099_ ) );
sky130_fd_sc_hd__xor2_1 _2757_ ( .A(\w3\[11\] ), .B(_1099_ ), .X(_1487_ ) );
sky130_fd_sc_hd__xnor3_1 _2758_ ( .A(\us32\/_0011_ ), .B(\us32\/_0012_ ), .C(\us32\/_0015_ ), .X(_1100_ ) );
sky130_fd_sc_hd__xnor3_1 _2759_ ( .A(_0747_ ), .B(_0933_ ), .C(_1100_ ), .X(_1101_ ) );
sky130_fd_sc_hd__nand2_1 _2760_ ( .A(_1101_ ), .B(_1086_ ), .Y(_1102_ ) );
sky130_fd_sc_hd__nand2_1 _2761_ ( .A(\text_in_r\[12\] ), .B(_1009_ ), .Y(_1103_ ) );
sky130_fd_sc_hd__nand2_1 _2762_ ( .A(_1102_ ), .B(_1103_ ), .Y(_1104_ ) );
sky130_fd_sc_hd__xor2_1 _2763_ ( .A(\w3\[12\] ), .B(_1104_ ), .X(_1488_ ) );
sky130_fd_sc_hd__xor3_1 _2764_ ( .A(\us32\/_0013_ ), .B(_0739_ ), .C(_0751_ ), .X(_1105_ ) );
sky130_fd_sc_hd__nand2_1 _2765_ ( .A(_1105_ ), .B(_1024_ ), .Y(_1106_ ) );
sky130_fd_sc_hd__or2b_1 _2766_ ( .A(\text_in_r\[13\] ), .B_N(_1069_ ), .X(_1107_ ) );
sky130_fd_sc_hd__nand2_1 _2767_ ( .A(_1106_ ), .B(_1107_ ), .Y(_1108_ ) );
sky130_fd_sc_hd__xnor2_1 _2768_ ( .A(\w3\[13\] ), .B(_1108_ ), .Y(_1489_ ) );
sky130_fd_sc_hd__xnor3_1 _2769_ ( .A(\us03\/_0014_ ), .B(_0752_ ), .C(_0940_ ), .X(_1109_ ) );
sky130_fd_sc_hd__nand2_1 _2770_ ( .A(_1109_ ), .B(_1024_ ), .Y(_1110_ ) );
sky130_fd_sc_hd__or2b_1 _2771_ ( .A(\text_in_r\[14\] ), .B_N(_1069_ ), .X(_1111_ ) );
sky130_fd_sc_hd__nand2_1 _2772_ ( .A(_1110_ ), .B(_1111_ ), .Y(_1112_ ) );
sky130_fd_sc_hd__xnor2_1 _2773_ ( .A(\w3\[14\] ), .B(_1112_ ), .Y(_1490_ ) );
sky130_fd_sc_hd__and2_0 _2774_ ( .A(\text_in_r\[15\] ), .B(_1077_ ), .X(_1113_ ) );
sky130_fd_sc_hd__xor2_1 _2775_ ( .A(_1387_ ), .B(\us03\/_0015_ ), .X(_1114_ ) );
sky130_fd_sc_hd__xor3_1 _2776_ ( .A(\us32\/_0015_ ), .B(_0947_ ), .C(_1114_ ), .X(_1115_ ) );
sky130_fd_sc_hd__nor2_1 _2777_ ( .A(_0898_ ), .B(_1115_ ), .Y(_1116_ ) );
sky130_fd_sc_hd__nor2_1 _2778_ ( .A(_1113_ ), .B(_1116_ ), .Y(_1117_ ) );
sky130_fd_sc_hd__xnor2_1 _2779_ ( .A(\w3\[15\] ), .B(_1117_ ), .Y(_1491_ ) );
sky130_fd_sc_hd__and2_0 _2780_ ( .A(\text_in_r\[96\] ), .B(_1077_ ), .X(_1118_ ) );
sky130_fd_sc_hd__xor3_1 _2781_ ( .A(\us33\/_0015_ ), .B(_0533_ ), .C(_0543_ ), .X(_1119_ ) );
sky130_fd_sc_hd__nor2_1 _2782_ ( .A(_0898_ ), .B(_1119_ ), .Y(_1120_ ) );
sky130_fd_sc_hd__nor2_1 _2783_ ( .A(_1118_ ), .B(_1120_ ), .Y(_1121_ ) );
sky130_fd_sc_hd__xnor2_1 _2784_ ( .A(\w0\[0\] ), .B(_1121_ ), .Y(_1492_ ) );
sky130_fd_sc_hd__and2_0 _2785_ ( .A(\text_in_r\[97\] ), .B(_1077_ ), .X(_1122_ ) );
sky130_fd_sc_hd__xnor3_1 _2786_ ( .A(\us00\/_0015_ ), .B(\us00\/_0008_ ), .C(\us22\/_0009_ ), .X(_1123_ ) );
sky130_fd_sc_hd__xnor3_1 _2787_ ( .A(_0557_ ), .B(_0957_ ), .C(_1123_ ), .X(_1124_ ) );
sky130_fd_sc_hd__nor2_1 _2788_ ( .A(_0898_ ), .B(_1124_ ), .Y(_1125_ ) );
sky130_fd_sc_hd__nor2_1 _2789_ ( .A(_1122_ ), .B(_1125_ ), .Y(_1126_ ) );
sky130_fd_sc_hd__xnor2_1 _2790_ ( .A(\w0\[1\] ), .B(_1126_ ), .Y(_1493_ ) );
sky130_fd_sc_hd__xnor3_1 _2791_ ( .A(\us33\/_0009_ ), .B(\us00\/_0010_ ), .C(_0556_ ), .X(_1127_ ) );
sky130_fd_sc_hd__xor3_1 _2792_ ( .A(\us00\/_0009_ ), .B(\us11\/_0010_ ), .C(_1127_ ), .X(_1128_ ) );
sky130_fd_sc_hd__nand2_1 _2793_ ( .A(_1128_ ), .B(_1086_ ), .Y(_1129_ ) );
sky130_fd_sc_hd__nand2_1 _2794_ ( .A(\text_in_r\[98\] ), .B(_1009_ ), .Y(_1130_ ) );
sky130_fd_sc_hd__nand2_1 _2795_ ( .A(_1129_ ), .B(_1130_ ), .Y(_1131_ ) );
sky130_fd_sc_hd__xor2_1 _2796_ ( .A(\w0\[2\] ), .B(_1131_ ), .X(_1494_ ) );
sky130_fd_sc_hd__xnor2_1 _2797_ ( .A(\us33\/_0010_ ), .B(\us33\/_0015_ ), .Y(_1132_ ) );
sky130_fd_sc_hd__xor2_1 _2798_ ( .A(\us22\/_0011_ ), .B(_0565_ ), .X(_1133_ ) );
sky130_fd_sc_hd__xor3_1 _2799_ ( .A(_0971_ ), .B(_1132_ ), .C(_1133_ ), .X(_1134_ ) );
sky130_fd_sc_hd__nand2_1 _2800_ ( .A(_1134_ ), .B(_1024_ ), .Y(_1135_ ) );
sky130_fd_sc_hd__or2b_1 _2801_ ( .A(\text_in_r\[99\] ), .B_N(_1069_ ), .X(_1136_ ) );
sky130_fd_sc_hd__nand2_1 _2802_ ( .A(_1135_ ), .B(_1136_ ), .Y(_1137_ ) );
sky130_fd_sc_hd__xnor2_1 _2803_ ( .A(\w0\[3\] ), .B(_1137_ ), .Y(_1495_ ) );
sky130_fd_sc_hd__xor2_1 _2804_ ( .A(\us33\/_0011_ ), .B(\us33\/_0015_ ), .X(_1138_ ) );
sky130_fd_sc_hd__xor2_1 _2805_ ( .A(_0796_ ), .B(_0572_ ), .X(_1139_ ) );
sky130_fd_sc_hd__xor3_1 _2806_ ( .A(_0579_ ), .B(_1138_ ), .C(_1139_ ), .X(_1140_ ) );
sky130_fd_sc_hd__nand2_1 _2807_ ( .A(_1140_ ), .B(_1024_ ), .Y(_1141_ ) );
sky130_fd_sc_hd__or2b_1 _2808_ ( .A(\text_in_r\[100\] ), .B_N(_1069_ ), .X(_1142_ ) );
sky130_fd_sc_hd__nand2_1 _2809_ ( .A(_1141_ ), .B(_1142_ ), .Y(_1143_ ) );
sky130_fd_sc_hd__xnor2_1 _2810_ ( .A(\w0\[4\] ), .B(_1143_ ), .Y(_1496_ ) );
sky130_fd_sc_hd__and2b_1 _2811_ ( .A_N(\text_in_r\[101\] ), .B(_0549_ ), .X(_1144_ ) );
sky130_fd_sc_hd__xnor3_1 _2812_ ( .A(\us33\/_0012_ ), .B(\us22\/_0013_ ), .C(\us00\/_0013_ ), .X(_1145_ ) );
sky130_fd_sc_hd__xnor3_1 _2813_ ( .A(\us00\/_0012_ ), .B(_1377_ ), .C(_1145_ ), .X(_1146_ ) );
sky130_fd_sc_hd__nor2_1 _2814_ ( .A(_0921_ ), .B(_1146_ ), .Y(_1147_ ) );
sky130_fd_sc_hd__nor2_1 _2815_ ( .A(_1144_ ), .B(_1147_ ), .Y(_1148_ ) );
sky130_fd_sc_hd__xor2_1 _2816_ ( .A(\w0\[5\] ), .B(_1148_ ), .X(_1497_ ) );
sky130_fd_sc_hd__and2b_1 _2817_ ( .A_N(\text_in_r\[102\] ), .B(_0549_ ), .X(_1149_ ) );
sky130_fd_sc_hd__xnor3_1 _2818_ ( .A(\us22\/_0014_ ), .B(\us00\/_0014_ ), .C(_0795_ ), .X(_1150_ ) );
sky130_fd_sc_hd__xor3_1 _2819_ ( .A(\us00\/_0013_ ), .B(\us11\/_0014_ ), .C(_1150_ ), .X(_1151_ ) );
sky130_fd_sc_hd__nor2_1 _2820_ ( .A(_0921_ ), .B(_1151_ ), .Y(_1152_ ) );
sky130_fd_sc_hd__nor2_1 _2821_ ( .A(_1149_ ), .B(_1152_ ), .Y(_1153_ ) );
sky130_fd_sc_hd__xor2_1 _2822_ ( .A(\w0\[6\] ), .B(_1153_ ), .X(_1498_ ) );
sky130_fd_sc_hd__xor3_1 _2823_ ( .A(\us33\/_0014_ ), .B(_0592_ ), .C(_0991_ ), .X(_1154_ ) );
sky130_fd_sc_hd__nand2_1 _2824_ ( .A(_1154_ ), .B(_0547_ ), .Y(_1155_ ) );
sky130_fd_sc_hd__or2b_1 _2825_ ( .A(\text_in_r\[103\] ), .B_N(_1069_ ), .X(_1156_ ) );
sky130_fd_sc_hd__nand2_1 _2826_ ( .A(_1155_ ), .B(_1156_ ), .Y(_1157_ ) );
sky130_fd_sc_hd__xnor2_1 _2827_ ( .A(\w0\[7\] ), .B(_1157_ ), .Y(_1499_ ) );
sky130_fd_sc_hd__xor3_1 _2828_ ( .A(_0646_ ), .B(_0599_ ), .C(_0604_ ), .X(_1158_ ) );
sky130_fd_sc_hd__nand2_1 _2829_ ( .A(_1158_ ), .B(_0547_ ), .Y(_1159_ ) );
sky130_fd_sc_hd__or2b_1 _2830_ ( .A(\text_in_r\[64\] ), .B_N(_1069_ ), .X(_1160_ ) );
sky130_fd_sc_hd__nand2_1 _2831_ ( .A(_1159_ ), .B(_1160_ ), .Y(_1161_ ) );
sky130_fd_sc_hd__xnor2_1 _2832_ ( .A(\w1\[0\] ), .B(_1161_ ), .Y(_1516_ ) );
sky130_fd_sc_hd__xnor3_1 _2833_ ( .A(\us01\/_0015_ ), .B(\us01\/_0008_ ), .C(\us23\/_0009_ ), .X(_1162_ ) );
sky130_fd_sc_hd__xnor3_1 _2834_ ( .A(_0613_ ), .B(_0997_ ), .C(_1162_ ), .X(_1163_ ) );
sky130_fd_sc_hd__nand2_1 _2835_ ( .A(_1163_ ), .B(_0547_ ), .Y(_1164_ ) );
sky130_fd_sc_hd__or2b_1 _2836_ ( .A(\text_in_r\[65\] ), .B_N(_1069_ ), .X(_1165_ ) );
sky130_fd_sc_hd__nand2_1 _2837_ ( .A(_1164_ ), .B(_1165_ ), .Y(_1166_ ) );
sky130_fd_sc_hd__xnor2_1 _2838_ ( .A(\w1\[1\] ), .B(_1166_ ), .Y(_1517_ ) );
sky130_fd_sc_hd__xnor3_1 _2839_ ( .A(\us30\/_0009_ ), .B(\us01\/_0010_ ), .C(_0612_ ), .X(_1167_ ) );
sky130_fd_sc_hd__xor3_1 _2840_ ( .A(\us01\/_0009_ ), .B(\us12\/_0010_ ), .C(_1167_ ), .X(_1168_ ) );
sky130_fd_sc_hd__nand2_1 _2841_ ( .A(_1168_ ), .B(_1086_ ), .Y(_1169_ ) );
sky130_fd_sc_hd__nand2_1 _2842_ ( .A(\text_in_r\[66\] ), .B(_1009_ ), .Y(_1170_ ) );
sky130_fd_sc_hd__nand2_1 _2843_ ( .A(_1169_ ), .B(_1170_ ), .Y(_1171_ ) );
sky130_fd_sc_hd__xor2_1 _2844_ ( .A(\w1\[2\] ), .B(_1171_ ), .X(_1518_ ) );
sky130_fd_sc_hd__and2_0 _2845_ ( .A(\text_in_r\[67\] ), .B(_1077_ ), .X(_1172_ ) );
sky130_fd_sc_hd__xnor2_1 _2846_ ( .A(\us30\/_0010_ ), .B(_0646_ ), .Y(_1173_ ) );
sky130_fd_sc_hd__xor2_1 _2847_ ( .A(\us23\/_0011_ ), .B(_0619_ ), .X(_1174_ ) );
sky130_fd_sc_hd__xor3_1 _2848_ ( .A(_1012_ ), .B(_1173_ ), .C(_1174_ ), .X(_1175_ ) );
sky130_fd_sc_hd__nor2_1 _2849_ ( .A(_0898_ ), .B(_1175_ ), .Y(_1176_ ) );
sky130_fd_sc_hd__nor2_1 _2850_ ( .A(_1172_ ), .B(_1176_ ), .Y(_1177_ ) );
sky130_fd_sc_hd__xnor2_1 _2851_ ( .A(\w1\[3\] ), .B(_1177_ ), .Y(_1519_ ) );
sky130_fd_sc_hd__and2_0 _2852_ ( .A(\text_in_r\[68\] ), .B(_1077_ ), .X(_1178_ ) );
sky130_fd_sc_hd__xor2_1 _2853_ ( .A(\us30\/_0011_ ), .B(_0646_ ), .X(_1179_ ) );
sky130_fd_sc_hd__xor2_1 _2854_ ( .A(\us23\/_0012_ ), .B(_0625_ ), .X(_1180_ ) );
sky130_fd_sc_hd__xnor3_1 _2855_ ( .A(_0633_ ), .B(_1179_ ), .C(_1180_ ), .X(_1181_ ) );
sky130_fd_sc_hd__nor2_1 _2856_ ( .A(_0898_ ), .B(_1181_ ), .Y(_1182_ ) );
sky130_fd_sc_hd__nor2_1 _2857_ ( .A(_1178_ ), .B(_1182_ ), .Y(_1183_ ) );
sky130_fd_sc_hd__xnor2_1 _2858_ ( .A(\w1\[4\] ), .B(_1183_ ), .Y(_1520_ ) );
sky130_fd_sc_hd__xnor3_1 _2859_ ( .A(\us30\/_0012_ ), .B(\us23\/_0013_ ), .C(\us01\/_0013_ ), .X(_1184_ ) );
sky130_fd_sc_hd__xnor3_1 _2860_ ( .A(\us01\/_0012_ ), .B(\us12\/_0013_ ), .C(_1184_ ), .X(_1185_ ) );
sky130_fd_sc_hd__nand2_1 _2861_ ( .A(_1185_ ), .B(_1086_ ), .Y(_1186_ ) );
sky130_fd_sc_hd__nand2_1 _2862_ ( .A(\text_in_r\[69\] ), .B(_1009_ ), .Y(_1187_ ) );
sky130_fd_sc_hd__nand2_1 _2863_ ( .A(_1186_ ), .B(_1187_ ), .Y(_1188_ ) );
sky130_fd_sc_hd__xor2_1 _2864_ ( .A(\w1\[5\] ), .B(_1188_ ), .X(_1521_ ) );
sky130_fd_sc_hd__and2b_1 _2865_ ( .A_N(\text_in_r\[70\] ), .B(_0549_ ), .X(_1189_ ) );
sky130_fd_sc_hd__xnor3_1 _2866_ ( .A(\us30\/_0013_ ), .B(\us23\/_0014_ ), .C(\us01\/_0014_ ), .X(_1190_ ) );
sky130_fd_sc_hd__xnor3_1 _2867_ ( .A(\us01\/_0013_ ), .B(\us12\/_0014_ ), .C(_1190_ ), .X(_1191_ ) );
sky130_fd_sc_hd__nor2_1 _2868_ ( .A(_0921_ ), .B(_1191_ ), .Y(_1192_ ) );
sky130_fd_sc_hd__nor2_1 _2869_ ( .A(_1189_ ), .B(_1192_ ), .Y(_1193_ ) );
sky130_fd_sc_hd__xor2_1 _2870_ ( .A(\w1\[6\] ), .B(_1193_ ), .X(_1522_ ) );
sky130_fd_sc_hd__xor3_1 _2871_ ( .A(\us30\/_0014_ ), .B(_0648_ ), .C(_1032_ ), .X(_1194_ ) );
sky130_fd_sc_hd__nand2_1 _2872_ ( .A(_1194_ ), .B(_0547_ ), .Y(_1195_ ) );
sky130_fd_sc_hd__or2b_1 _2873_ ( .A(\text_in_r\[71\] ), .B_N(_1069_ ), .X(_1196_ ) );
sky130_fd_sc_hd__nand2_1 _2874_ ( .A(_1195_ ), .B(_1196_ ), .Y(_1197_ ) );
sky130_fd_sc_hd__xnor2_1 _2875_ ( .A(\w1\[7\] ), .B(_1197_ ), .Y(_1523_ ) );
sky130_fd_sc_hd__xor3_1 _2876_ ( .A(\us31\/_0015_ ), .B(_0655_ ), .C(_0660_ ), .X(_1198_ ) );
sky130_fd_sc_hd__nand2_1 _2877_ ( .A(_1198_ ), .B(_0547_ ), .Y(_1199_ ) );
sky130_fd_sc_hd__or2b_1 _2878_ ( .A(\text_in_r\[32\] ), .B_N(_0536_ ), .X(_1200_ ) );
sky130_fd_sc_hd__nand2_1 _2879_ ( .A(_1199_ ), .B(_1200_ ), .Y(_1201_ ) );
sky130_fd_sc_hd__xnor2_1 _2880_ ( .A(\w2\[0\] ), .B(_1201_ ), .Y(_1532_ ) );
sky130_fd_sc_hd__and2_0 _2881_ ( .A(\text_in_r\[33\] ), .B(_1077_ ), .X(_1202_ ) );
sky130_fd_sc_hd__xnor3_1 _2882_ ( .A(\us02\/_0015_ ), .B(\us02\/_0008_ ), .C(\us20\/_0009_ ), .X(_1203_ ) );
sky130_fd_sc_hd__xnor3_1 _2883_ ( .A(_0669_ ), .B(_1039_ ), .C(_1203_ ), .X(_1204_ ) );
sky130_fd_sc_hd__nor2_1 _2884_ ( .A(_0564_ ), .B(_1204_ ), .Y(_1205_ ) );
sky130_fd_sc_hd__nor2_1 _2885_ ( .A(_1202_ ), .B(_1205_ ), .Y(_1206_ ) );
sky130_fd_sc_hd__xnor2_1 _2886_ ( .A(\w2\[1\] ), .B(_1206_ ), .Y(_1533_ ) );
sky130_fd_sc_hd__xnor3_1 _2887_ ( .A(\us31\/_0009_ ), .B(\us02\/_0010_ ), .C(_0668_ ), .X(_1207_ ) );
sky130_fd_sc_hd__xor3_1 _2888_ ( .A(\us02\/_0009_ ), .B(\us13\/_0010_ ), .C(_1207_ ), .X(_1208_ ) );
sky130_fd_sc_hd__nand2_1 _2889_ ( .A(_1208_ ), .B(_1086_ ), .Y(_1209_ ) );
sky130_fd_sc_hd__nand2_1 _2890_ ( .A(\text_in_r\[34\] ), .B(_0555_ ), .Y(_1210_ ) );
sky130_fd_sc_hd__nand2_1 _2891_ ( .A(_1209_ ), .B(_1210_ ), .Y(_1211_ ) );
sky130_fd_sc_hd__xor2_1 _2892_ ( .A(\w2\[2\] ), .B(_1211_ ), .X(_1534_ ) );
sky130_fd_sc_hd__and2_0 _2893_ ( .A(\text_in_r\[35\] ), .B(_1077_ ), .X(_1212_ ) );
sky130_fd_sc_hd__xnor2_1 _2894_ ( .A(\us31\/_0010_ ), .B(\us31\/_0015_ ), .Y(_1213_ ) );
sky130_fd_sc_hd__xor2_1 _2895_ ( .A(\us20\/_0011_ ), .B(_0675_ ), .X(_1214_ ) );
sky130_fd_sc_hd__xor3_1 _2896_ ( .A(_1053_ ), .B(_1213_ ), .C(_1214_ ), .X(_1215_ ) );
sky130_fd_sc_hd__nor2_1 _2897_ ( .A(_0564_ ), .B(_1215_ ), .Y(_1216_ ) );
sky130_fd_sc_hd__nor2_1 _2898_ ( .A(_1212_ ), .B(_1216_ ), .Y(_1217_ ) );
sky130_fd_sc_hd__xnor2_1 _2899_ ( .A(\w2\[3\] ), .B(_1217_ ), .Y(_1535_ ) );
sky130_fd_sc_hd__and2_0 _2900_ ( .A(\text_in_r\[36\] ), .B(_1077_ ), .X(_1218_ ) );
sky130_fd_sc_hd__xor2_1 _2901_ ( .A(\us31\/_0011_ ), .B(\us31\/_0015_ ), .X(_1219_ ) );
sky130_fd_sc_hd__xor2_1 _2902_ ( .A(\us20\/_0012_ ), .B(_0684_ ), .X(_1220_ ) );
sky130_fd_sc_hd__xnor3_1 _2903_ ( .A(_0692_ ), .B(_1219_ ), .C(_1220_ ), .X(_1221_ ) );
sky130_fd_sc_hd__nor2_1 _2904_ ( .A(_0564_ ), .B(_1221_ ), .Y(_1222_ ) );
sky130_fd_sc_hd__nor2_1 _2905_ ( .A(_1218_ ), .B(_1222_ ), .Y(_1223_ ) );
sky130_fd_sc_hd__xnor2_1 _2906_ ( .A(\w2\[4\] ), .B(_1223_ ), .Y(_1536_ ) );
sky130_fd_sc_hd__xnor3_1 _2907_ ( .A(\us31\/_0012_ ), .B(\us20\/_0013_ ), .C(\us02\/_0013_ ), .X(_1224_ ) );
sky130_fd_sc_hd__xnor3_1 _2908_ ( .A(\us02\/_0012_ ), .B(\us13\/_0013_ ), .C(_1224_ ), .X(_1225_ ) );
sky130_fd_sc_hd__nand2_1 _2909_ ( .A(_1225_ ), .B(_1086_ ), .Y(_1226_ ) );
sky130_fd_sc_hd__nand2_1 _2910_ ( .A(\text_in_r\[37\] ), .B(_0555_ ), .Y(_1227_ ) );
sky130_fd_sc_hd__nand2_1 _2911_ ( .A(_1226_ ), .B(_1227_ ), .Y(_1228_ ) );
sky130_fd_sc_hd__xor2_1 _2912_ ( .A(\w2\[5\] ), .B(_1228_ ), .X(_1537_ ) );
sky130_fd_sc_hd__xnor3_1 _2913_ ( .A(\us31\/_0013_ ), .B(\us20\/_0014_ ), .C(\us02\/_0014_ ), .X(_1229_ ) );
sky130_fd_sc_hd__xnor3_1 _2914_ ( .A(\us02\/_0013_ ), .B(\us13\/_0014_ ), .C(_1229_ ), .X(_1230_ ) );
sky130_fd_sc_hd__nand2_1 _2915_ ( .A(_1230_ ), .B(_1086_ ), .Y(_1231_ ) );
sky130_fd_sc_hd__nand2_1 _2916_ ( .A(\text_in_r\[38\] ), .B(_0555_ ), .Y(_1232_ ) );
sky130_fd_sc_hd__nand2_1 _2917_ ( .A(_1231_ ), .B(_1232_ ), .Y(_1233_ ) );
sky130_fd_sc_hd__xor2_1 _2918_ ( .A(\w2\[6\] ), .B(_1233_ ), .X(_1538_ ) );
sky130_fd_sc_hd__and2_0 _2919_ ( .A(\text_in_r\[39\] ), .B(_1077_ ), .X(_1234_ ) );
sky130_fd_sc_hd__xor3_1 _2920_ ( .A(\us31\/_0014_ ), .B(_0705_ ), .C(_1072_ ), .X(_1235_ ) );
sky130_fd_sc_hd__nor2_1 _2921_ ( .A(_0564_ ), .B(_1235_ ), .Y(_1236_ ) );
sky130_fd_sc_hd__nor2_1 _2922_ ( .A(_1234_ ), .B(_1236_ ), .Y(_1237_ ) );
sky130_fd_sc_hd__xnor2_1 _2923_ ( .A(\w2\[7\] ), .B(_1237_ ), .Y(_1539_ ) );
sky130_fd_sc_hd__and2_0 _2924_ ( .A(\text_in_r\[0\] ), .B(_0562_ ), .X(_1238_ ) );
sky130_fd_sc_hd__xor3_1 _2925_ ( .A(\us32\/_0015_ ), .B(_0712_ ), .C(_0718_ ), .X(_1239_ ) );
sky130_fd_sc_hd__nor2_1 _2926_ ( .A(_0564_ ), .B(_1239_ ), .Y(_1240_ ) );
sky130_fd_sc_hd__nor2_1 _2927_ ( .A(_1238_ ), .B(_1240_ ), .Y(_1241_ ) );
sky130_fd_sc_hd__xnor2_1 _2928_ ( .A(\w3\[0\] ), .B(_1241_ ), .Y(_1548_ ) );
sky130_fd_sc_hd__and2_0 _2929_ ( .A(\text_in_r\[1\] ), .B(_0562_ ), .X(_1242_ ) );
sky130_fd_sc_hd__xnor3_1 _2930_ ( .A(\us03\/_0015_ ), .B(\us03\/_0008_ ), .C(\us21\/_0009_ ), .X(_1243_ ) );
sky130_fd_sc_hd__xnor3_1 _2931_ ( .A(_0725_ ), .B(_1080_ ), .C(_1243_ ), .X(_1244_ ) );
sky130_fd_sc_hd__nor2_1 _2932_ ( .A(_0564_ ), .B(_1244_ ), .Y(_1245_ ) );
sky130_fd_sc_hd__nor2_1 _2933_ ( .A(_1242_ ), .B(_1245_ ), .Y(_1246_ ) );
sky130_fd_sc_hd__xnor2_1 _2934_ ( .A(\w3\[1\] ), .B(_1246_ ), .Y(_1549_ ) );
sky130_fd_sc_hd__xnor3_1 _2935_ ( .A(\us32\/_0009_ ), .B(\us03\/_0010_ ), .C(_0724_ ), .X(_1247_ ) );
sky130_fd_sc_hd__xor3_1 _2936_ ( .A(\us03\/_0009_ ), .B(\us10\/_0010_ ), .C(_1247_ ), .X(_1248_ ) );
sky130_fd_sc_hd__nand2_1 _2937_ ( .A(_1248_ ), .B(_0537_ ), .Y(_1249_ ) );
sky130_fd_sc_hd__nand2_1 _2938_ ( .A(\text_in_r\[2\] ), .B(_0555_ ), .Y(_1250_ ) );
sky130_fd_sc_hd__nand2_1 _2939_ ( .A(_1249_ ), .B(_1250_ ), .Y(_1251_ ) );
sky130_fd_sc_hd__xor2_1 _2940_ ( .A(\w3\[2\] ), .B(_1251_ ), .X(_1550_ ) );
sky130_fd_sc_hd__xnor2_1 _2941_ ( .A(\us32\/_0010_ ), .B(\us32\/_0015_ ), .Y(_1252_ ) );
sky130_fd_sc_hd__xor2_1 _2942_ ( .A(\us21\/_0011_ ), .B(_0732_ ), .X(_1253_ ) );
sky130_fd_sc_hd__xor3_1 _2943_ ( .A(_1094_ ), .B(_1252_ ), .C(_1253_ ), .X(_1254_ ) );
sky130_fd_sc_hd__nand2_1 _2944_ ( .A(_1254_ ), .B(_0547_ ), .Y(_1255_ ) );
sky130_fd_sc_hd__or2b_1 _2945_ ( .A(\text_in_r\[3\] ), .B_N(_0536_ ), .X(_1256_ ) );
sky130_fd_sc_hd__nand2_1 _2946_ ( .A(_1255_ ), .B(_1256_ ), .Y(_1257_ ) );
sky130_fd_sc_hd__xnor2_1 _2947_ ( .A(\w3\[3\] ), .B(_1257_ ), .Y(_1551_ ) );
sky130_fd_sc_hd__xor2_1 _2948_ ( .A(\us32\/_0011_ ), .B(\us32\/_0015_ ), .X(_1258_ ) );
sky130_fd_sc_hd__xor2_1 _2949_ ( .A(\us21\/_0012_ ), .B(_0738_ ), .X(_1259_ ) );
sky130_fd_sc_hd__xnor3_1 _2950_ ( .A(_0747_ ), .B(_1258_ ), .C(_1259_ ), .X(_1260_ ) );
sky130_fd_sc_hd__nand2_1 _2951_ ( .A(_1260_ ), .B(_0547_ ), .Y(_1261_ ) );
sky130_fd_sc_hd__or2b_1 _2952_ ( .A(\text_in_r\[4\] ), .B_N(_0536_ ), .X(_1262_ ) );
sky130_fd_sc_hd__nand2_1 _2953_ ( .A(_1261_ ), .B(_1262_ ), .Y(_1263_ ) );
sky130_fd_sc_hd__xnor2_1 _2954_ ( .A(\w3\[4\] ), .B(_1263_ ), .Y(_1552_ ) );
sky130_fd_sc_hd__and2b_1 _2955_ ( .A_N(\text_in_r\[5\] ), .B(_0549_ ), .X(_1264_ ) );
sky130_fd_sc_hd__xnor3_1 _2956_ ( .A(\us32\/_0012_ ), .B(\us21\/_0013_ ), .C(\us03\/_0013_ ), .X(_1265_ ) );
sky130_fd_sc_hd__xnor3_1 _2957_ ( .A(\us03\/_0012_ ), .B(\us10\/_0013_ ), .C(_1265_ ), .X(_1266_ ) );
sky130_fd_sc_hd__nor2_1 _2958_ ( .A(ld_r ), .B(_1266_ ), .Y(_1267_ ) );
sky130_fd_sc_hd__nor2_1 _2959_ ( .A(_1264_ ), .B(_1267_ ), .Y(_1268_ ) );
sky130_fd_sc_hd__xor2_1 _2960_ ( .A(\w3\[5\] ), .B(_1268_ ), .X(_1553_ ) );
sky130_fd_sc_hd__xnor3_1 _2961_ ( .A(\us32\/_0013_ ), .B(\us21\/_0014_ ), .C(\us03\/_0014_ ), .X(_1269_ ) );
sky130_fd_sc_hd__xnor3_1 _2962_ ( .A(\us03\/_0013_ ), .B(\us10\/_0014_ ), .C(_1269_ ), .X(_1270_ ) );
sky130_fd_sc_hd__nand2_1 _2963_ ( .A(_1270_ ), .B(_0537_ ), .Y(_1271_ ) );
sky130_fd_sc_hd__nand2_1 _2964_ ( .A(\text_in_r\[6\] ), .B(_0555_ ), .Y(_1272_ ) );
sky130_fd_sc_hd__nand2_1 _2965_ ( .A(_1271_ ), .B(_1272_ ), .Y(_1273_ ) );
sky130_fd_sc_hd__xor2_1 _2966_ ( .A(\w3\[6\] ), .B(_1273_ ), .X(_1554_ ) );
sky130_fd_sc_hd__and2_0 _2967_ ( .A(\text_in_r\[7\] ), .B(_0562_ ), .X(_1274_ ) );
sky130_fd_sc_hd__xor3_1 _2968_ ( .A(\us32\/_0014_ ), .B(_0759_ ), .C(_1114_ ), .X(_1275_ ) );
sky130_fd_sc_hd__nor2_1 _2969_ ( .A(_0564_ ), .B(_1275_ ), .Y(_1276_ ) );
sky130_fd_sc_hd__nor2_1 _2970_ ( .A(_1274_ ), .B(_1276_ ), .Y(_1277_ ) );
sky130_fd_sc_hd__xnor2_1 _2971_ ( .A(\w3\[7\] ), .B(_1277_ ), .Y(_1555_ ) );
sky130_fd_sc_hd__xor2_1 _2972_ ( .A(\w0\[24\] ), .B(\us00\/_0008_ ), .X(_0418_ ) );
sky130_fd_sc_hd__xor2_1 _2973_ ( .A(\w0\[25\] ), .B(\us00\/_0009_ ), .X(_0419_ ) );
sky130_fd_sc_hd__xor2_1 _2974_ ( .A(\w0\[26\] ), .B(\us00\/_0010_ ), .X(_0420_ ) );
sky130_fd_sc_hd__xor2_1 _2975_ ( .A(\w0\[27\] ), .B(\us00\/_0011_ ), .X(_0421_ ) );
sky130_fd_sc_hd__xor2_1 _2976_ ( .A(\w0\[28\] ), .B(\us00\/_0012_ ), .X(_0422_ ) );
sky130_fd_sc_hd__xor2_1 _2977_ ( .A(\w0\[29\] ), .B(\us00\/_0013_ ), .X(_0423_ ) );
sky130_fd_sc_hd__xor2_1 _2978_ ( .A(\w0\[30\] ), .B(\us00\/_0014_ ), .X(_0424_ ) );
sky130_fd_sc_hd__xor2_1 _2979_ ( .A(\us00\/_0015_ ), .B(\w0\[31\] ), .X(_0425_ ) );
sky130_fd_sc_hd__xor2_1 _2980_ ( .A(\w1\[24\] ), .B(\us01\/_0008_ ), .X(_0514_ ) );
sky130_fd_sc_hd__xor2_1 _2981_ ( .A(\w1\[25\] ), .B(\us01\/_0009_ ), .X(_0515_ ) );
sky130_fd_sc_hd__xor2_1 _2982_ ( .A(\w1\[26\] ), .B(\us01\/_0010_ ), .X(_0516_ ) );
sky130_fd_sc_hd__xor2_1 _2983_ ( .A(\w1\[27\] ), .B(\us01\/_0011_ ), .X(_0517_ ) );
sky130_fd_sc_hd__xor2_1 _2984_ ( .A(\w1\[28\] ), .B(\us01\/_0012_ ), .X(_0518_ ) );
sky130_fd_sc_hd__xor2_1 _2985_ ( .A(\w1\[29\] ), .B(\us01\/_0013_ ), .X(_0519_ ) );
sky130_fd_sc_hd__xor2_1 _2986_ ( .A(\w1\[30\] ), .B(\us01\/_0014_ ), .X(_0520_ ) );
sky130_fd_sc_hd__xor2_1 _2987_ ( .A(\us01\/_0015_ ), .B(\w1\[31\] ), .X(_0521_ ) );
sky130_fd_sc_hd__xor2_1 _2988_ ( .A(\w2\[24\] ), .B(\us02\/_0008_ ), .X(_0474_ ) );
sky130_fd_sc_hd__xor2_1 _2989_ ( .A(\w2\[25\] ), .B(\us02\/_0009_ ), .X(_0475_ ) );
sky130_fd_sc_hd__xor2_1 _2990_ ( .A(\w2\[26\] ), .B(\us02\/_0010_ ), .X(_0476_ ) );
sky130_fd_sc_hd__xor2_1 _2991_ ( .A(\w2\[27\] ), .B(\us02\/_0011_ ), .X(_0477_ ) );
sky130_fd_sc_hd__xor2_1 _2992_ ( .A(\w2\[28\] ), .B(\us02\/_0012_ ), .X(_0478_ ) );
sky130_fd_sc_hd__xor2_1 _2993_ ( .A(\w2\[29\] ), .B(\us02\/_0013_ ), .X(_0479_ ) );
sky130_fd_sc_hd__xor2_1 _2994_ ( .A(\w2\[30\] ), .B(\us02\/_0014_ ), .X(_0480_ ) );
sky130_fd_sc_hd__xor2_1 _2995_ ( .A(\us02\/_0015_ ), .B(\w2\[31\] ), .X(_0481_ ) );
sky130_fd_sc_hd__xor2_1 _2996_ ( .A(\w3\[24\] ), .B(\us03\/_0008_ ), .X(_0442_ ) );
sky130_fd_sc_hd__xor2_1 _2997_ ( .A(\w3\[25\] ), .B(\us03\/_0009_ ), .X(_0443_ ) );
sky130_fd_sc_hd__xor2_1 _2998_ ( .A(\w3\[26\] ), .B(\us03\/_0010_ ), .X(_0444_ ) );
sky130_fd_sc_hd__xor2_1 _2999_ ( .A(\w3\[27\] ), .B(\us03\/_0011_ ), .X(_0445_ ) );
sky130_fd_sc_hd__xor2_1 _3000_ ( .A(\w3\[28\] ), .B(\us03\/_0012_ ), .X(_0446_ ) );
sky130_fd_sc_hd__xor2_1 _3001_ ( .A(\w3\[29\] ), .B(\us03\/_0013_ ), .X(_0447_ ) );
sky130_fd_sc_hd__xor2_1 _3002_ ( .A(\w3\[30\] ), .B(\us03\/_0014_ ), .X(_0448_ ) );
sky130_fd_sc_hd__xor2_1 _3003_ ( .A(\us03\/_0015_ ), .B(\u0\/_0842_ ), .X(_0449_ ) );
sky130_fd_sc_hd__xor2_1 _3004_ ( .A(\us11\/_0008_ ), .B(\w0\[16\] ), .X(_0410_ ) );
sky130_fd_sc_hd__xor2_1 _3005_ ( .A(_1373_ ), .B(\w0\[17\] ), .X(_0411_ ) );
sky130_fd_sc_hd__xor2_1 _3006_ ( .A(\us11\/_0010_ ), .B(\w0\[18\] ), .X(_0412_ ) );
sky130_fd_sc_hd__xor2_1 _3007_ ( .A(\us11\/_0011_ ), .B(\w0\[19\] ), .X(_0413_ ) );
sky130_fd_sc_hd__xor2_1 _3008_ ( .A(\us11\/_0012_ ), .B(\w0\[20\] ), .X(_0414_ ) );
sky130_fd_sc_hd__xor2_1 _3009_ ( .A(_1377_ ), .B(\w0\[21\] ), .X(_0415_ ) );
sky130_fd_sc_hd__xor2_1 _3010_ ( .A(\us11\/_0014_ ), .B(\w0\[22\] ), .X(_0416_ ) );
sky130_fd_sc_hd__xor2_1 _3011_ ( .A(_1379_ ), .B(\w0\[23\] ), .X(_0417_ ) );
sky130_fd_sc_hd__xor2_1 _3012_ ( .A(\us12\/_0008_ ), .B(\w1\[16\] ), .X(_0506_ ) );
sky130_fd_sc_hd__xor2_1 _3013_ ( .A(\us12\/_0009_ ), .B(\w1\[17\] ), .X(_0507_ ) );
sky130_fd_sc_hd__xor2_1 _3014_ ( .A(\us12\/_0010_ ), .B(\w1\[18\] ), .X(_0508_ ) );
sky130_fd_sc_hd__xor2_1 _3015_ ( .A(\us12\/_0011_ ), .B(\w1\[19\] ), .X(_0509_ ) );
sky130_fd_sc_hd__xor2_1 _3016_ ( .A(\us12\/_0012_ ), .B(\w1\[20\] ), .X(_0510_ ) );
sky130_fd_sc_hd__xor2_1 _3017_ ( .A(\us12\/_0013_ ), .B(\w1\[21\] ), .X(_0511_ ) );
sky130_fd_sc_hd__xor2_1 _3018_ ( .A(\us12\/_0014_ ), .B(\w1\[22\] ), .X(_0512_ ) );
sky130_fd_sc_hd__xor2_1 _3019_ ( .A(\us12\/_0015_ ), .B(\w1\[23\] ), .X(_0513_ ) );
sky130_fd_sc_hd__xor2_1 _3020_ ( .A(\us13\/_0008_ ), .B(\w2\[16\] ), .X(_0466_ ) );
sky130_fd_sc_hd__xor2_1 _3021_ ( .A(\us13\/_0009_ ), .B(\w2\[17\] ), .X(_0467_ ) );
sky130_fd_sc_hd__xor2_1 _3022_ ( .A(\us13\/_0010_ ), .B(\w2\[18\] ), .X(_0468_ ) );
sky130_fd_sc_hd__xor2_1 _3023_ ( .A(\us13\/_0011_ ), .B(\w2\[19\] ), .X(_0469_ ) );
sky130_fd_sc_hd__xor2_1 _3024_ ( .A(\us13\/_0012_ ), .B(\w2\[20\] ), .X(_0470_ ) );
sky130_fd_sc_hd__xor2_1 _3025_ ( .A(\us13\/_0013_ ), .B(\w2\[21\] ), .X(_0471_ ) );
sky130_fd_sc_hd__xor2_1 _3026_ ( .A(\us13\/_0014_ ), .B(\w2\[22\] ), .X(_0472_ ) );
sky130_fd_sc_hd__xor2_1 _3027_ ( .A(_1419_ ), .B(\w2\[23\] ), .X(_0473_ ) );
sky130_fd_sc_hd__xor2_1 _3028_ ( .A(\us10\/_0008_ ), .B(\w3\[16\] ), .X(_0434_ ) );
sky130_fd_sc_hd__xor2_1 _3029_ ( .A(\us10\/_0009_ ), .B(\w3\[17\] ), .X(_0435_ ) );
sky130_fd_sc_hd__xor2_1 _3030_ ( .A(\us10\/_0010_ ), .B(\w3\[18\] ), .X(_0436_ ) );
sky130_fd_sc_hd__xor2_1 _3031_ ( .A(\us10\/_0011_ ), .B(\w3\[19\] ), .X(_0437_ ) );
sky130_fd_sc_hd__xor2_1 _3032_ ( .A(\us10\/_0012_ ), .B(\w3\[20\] ), .X(_0438_ ) );
sky130_fd_sc_hd__xor2_1 _3033_ ( .A(\us10\/_0013_ ), .B(\w3\[21\] ), .X(_0439_ ) );
sky130_fd_sc_hd__xor2_1 _3034_ ( .A(\us10\/_0014_ ), .B(\w3\[22\] ), .X(_0440_ ) );
sky130_fd_sc_hd__xor2_1 _3035_ ( .A(_1387_ ), .B(\w3\[23\] ), .X(_0441_ ) );
sky130_fd_sc_hd__xor2_1 _3036_ ( .A(\us22\/_0008_ ), .B(\w0\[8\] ), .X(_0402_ ) );
sky130_fd_sc_hd__xor2_1 _3037_ ( .A(\us22\/_0009_ ), .B(\w0\[9\] ), .X(_0403_ ) );
sky130_fd_sc_hd__xor2_1 _3038_ ( .A(\us22\/_0010_ ), .B(\w0\[10\] ), .X(_0404_ ) );
sky130_fd_sc_hd__xor2_1 _3039_ ( .A(\us22\/_0011_ ), .B(\w0\[11\] ), .X(_0405_ ) );
sky130_fd_sc_hd__xor2_2 _3040_ ( .A(\us22\/_0012_ ), .B(\w0\[12\] ), .X(_0406_ ) );
sky130_fd_sc_hd__xor2_1 _3041_ ( .A(\us22\/_0013_ ), .B(\w0\[13\] ), .X(_0407_ ) );
sky130_fd_sc_hd__xor2_1 _3042_ ( .A(\us22\/_0014_ ), .B(\w0\[14\] ), .X(_0408_ ) );
sky130_fd_sc_hd__xor2_1 _3043_ ( .A(\us22\/_0015_ ), .B(\w0\[15\] ), .X(_0409_ ) );
sky130_fd_sc_hd__xor2_1 _3044_ ( .A(\us23\/_0008_ ), .B(\w1\[8\] ), .X(_0490_ ) );
sky130_fd_sc_hd__xor2_1 _3045_ ( .A(\us23\/_0009_ ), .B(\w1\[9\] ), .X(_0491_ ) );
sky130_fd_sc_hd__xor2_1 _3046_ ( .A(\us23\/_0010_ ), .B(\w1\[10\] ), .X(_0492_ ) );
sky130_fd_sc_hd__xor2_1 _3047_ ( .A(\us23\/_0011_ ), .B(\w1\[11\] ), .X(_0493_ ) );
sky130_fd_sc_hd__xor2_1 _3048_ ( .A(\us23\/_0012_ ), .B(\w1\[12\] ), .X(_0494_ ) );
sky130_fd_sc_hd__xor2_1 _3049_ ( .A(\us23\/_0013_ ), .B(\w1\[13\] ), .X(_0495_ ) );
sky130_fd_sc_hd__xor2_1 _3050_ ( .A(\us23\/_0014_ ), .B(\w1\[14\] ), .X(_0496_ ) );
sky130_fd_sc_hd__xor2_1 _3051_ ( .A(\us23\/_0015_ ), .B(\w1\[15\] ), .X(_0497_ ) );
sky130_fd_sc_hd__xor2_1 _3052_ ( .A(\us20\/_0008_ ), .B(\w2\[8\] ), .X(_0458_ ) );
sky130_fd_sc_hd__xor2_1 _3053_ ( .A(\us20\/_0009_ ), .B(\w2\[9\] ), .X(_0459_ ) );
sky130_fd_sc_hd__xor2_1 _3054_ ( .A(\us20\/_0010_ ), .B(\w2\[10\] ), .X(_0460_ ) );
sky130_fd_sc_hd__xor2_1 _3055_ ( .A(\us20\/_0011_ ), .B(\w2\[11\] ), .X(_0461_ ) );
sky130_fd_sc_hd__xor2_2 _3056_ ( .A(\us20\/_0012_ ), .B(\w2\[12\] ), .X(_0462_ ) );
sky130_fd_sc_hd__xor2_1 _3057_ ( .A(\us20\/_0013_ ), .B(\w2\[13\] ), .X(_0463_ ) );
sky130_fd_sc_hd__xor2_1 _3058_ ( .A(\us20\/_0014_ ), .B(\w2\[14\] ), .X(_0464_ ) );
sky130_fd_sc_hd__xor2_1 _3059_ ( .A(_1451_ ), .B(\w2\[15\] ), .X(_0465_ ) );
sky130_fd_sc_hd__xor2_1 _3060_ ( .A(\us21\/_0008_ ), .B(\w3\[8\] ), .X(_0426_ ) );
sky130_fd_sc_hd__xor2_1 _3061_ ( .A(\us21\/_0009_ ), .B(\w3\[9\] ), .X(_0427_ ) );
sky130_fd_sc_hd__xor2_1 _3062_ ( .A(\us21\/_0010_ ), .B(\w3\[10\] ), .X(_0428_ ) );
sky130_fd_sc_hd__xor2_1 _3063_ ( .A(\us21\/_0011_ ), .B(\w3\[11\] ), .X(_0429_ ) );
sky130_fd_sc_hd__xor2_1 _3064_ ( .A(\us21\/_0012_ ), .B(\w3\[12\] ), .X(_0430_ ) );
sky130_fd_sc_hd__xor2_1 _3065_ ( .A(\us21\/_0013_ ), .B(\w3\[13\] ), .X(_0431_ ) );
sky130_fd_sc_hd__xor2_1 _3066_ ( .A(\us21\/_0014_ ), .B(\w3\[14\] ), .X(_0432_ ) );
sky130_fd_sc_hd__xor2_1 _3067_ ( .A(\us21\/_0015_ ), .B(\w3\[15\] ), .X(_0433_ ) );
sky130_fd_sc_hd__xor2_1 _3068_ ( .A(\us33\/_0008_ ), .B(\w0\[0\] ), .X(_0394_ ) );
sky130_fd_sc_hd__xor2_1 _3069_ ( .A(\us33\/_0009_ ), .B(\w0\[1\] ), .X(_0395_ ) );
sky130_fd_sc_hd__xor2_1 _3070_ ( .A(\us33\/_0010_ ), .B(\w0\[2\] ), .X(_0396_ ) );
sky130_fd_sc_hd__xor2_1 _3071_ ( .A(\us33\/_0011_ ), .B(\w0\[3\] ), .X(_0397_ ) );
sky130_fd_sc_hd__xor2_1 _3072_ ( .A(\us33\/_0012_ ), .B(\w0\[4\] ), .X(_0398_ ) );
sky130_fd_sc_hd__xor2_1 _3073_ ( .A(\us33\/_0013_ ), .B(\w0\[5\] ), .X(_0399_ ) );
sky130_fd_sc_hd__xor2_1 _3074_ ( .A(\us33\/_0014_ ), .B(\w0\[6\] ), .X(_0400_ ) );
sky130_fd_sc_hd__xor2_2 _3075_ ( .A(\us33\/_0015_ ), .B(\w0\[7\] ), .X(_0401_ ) );
sky130_fd_sc_hd__xor2_1 _3076_ ( .A(\us30\/_0008_ ), .B(\w1\[0\] ), .X(_0482_ ) );
sky130_fd_sc_hd__xor2_1 _3077_ ( .A(\us30\/_0009_ ), .B(\w1\[1\] ), .X(_0483_ ) );
sky130_fd_sc_hd__xor2_1 _3078_ ( .A(\us30\/_0010_ ), .B(\w1\[2\] ), .X(_0484_ ) );
sky130_fd_sc_hd__xor2_1 _3079_ ( .A(\us30\/_0011_ ), .B(\w1\[3\] ), .X(_0485_ ) );
sky130_fd_sc_hd__xor2_1 _3080_ ( .A(\us30\/_0012_ ), .B(\w1\[4\] ), .X(_0486_ ) );
sky130_fd_sc_hd__xor2_1 _3081_ ( .A(\us30\/_0013_ ), .B(\w1\[5\] ), .X(_0487_ ) );
sky130_fd_sc_hd__xor2_1 _3082_ ( .A(\us30\/_0014_ ), .B(\w1\[6\] ), .X(_0488_ ) );
sky130_fd_sc_hd__xor2_1 _3083_ ( .A(_0646_ ), .B(\w1\[7\] ), .X(_0489_ ) );
sky130_fd_sc_hd__xor2_1 _3084_ ( .A(\us31\/_0008_ ), .B(\w2\[0\] ), .X(_0450_ ) );
sky130_fd_sc_hd__xor2_1 _3085_ ( .A(\us31\/_0009_ ), .B(\w2\[1\] ), .X(_0451_ ) );
sky130_fd_sc_hd__xor2_1 _3086_ ( .A(\us31\/_0010_ ), .B(\w2\[2\] ), .X(_0452_ ) );
sky130_fd_sc_hd__xor2_1 _3087_ ( .A(\us31\/_0011_ ), .B(\w2\[3\] ), .X(_0453_ ) );
sky130_fd_sc_hd__xor2_1 _3088_ ( .A(\us31\/_0012_ ), .B(\w2\[4\] ), .X(_0454_ ) );
sky130_fd_sc_hd__xor2_1 _3089_ ( .A(\us31\/_0013_ ), .B(\w2\[5\] ), .X(_0455_ ) );
sky130_fd_sc_hd__xor2_1 _3090_ ( .A(\us31\/_0014_ ), .B(\w2\[6\] ), .X(_0456_ ) );
sky130_fd_sc_hd__xor2_1 _3091_ ( .A(\us31\/_0015_ ), .B(\w2\[7\] ), .X(_0457_ ) );
sky130_fd_sc_hd__xor2_1 _3092_ ( .A(\us32\/_0008_ ), .B(\w3\[0\] ), .X(_0498_ ) );
sky130_fd_sc_hd__xor2_1 _3093_ ( .A(\us32\/_0009_ ), .B(\w3\[1\] ), .X(_0499_ ) );
sky130_fd_sc_hd__xor2_1 _3094_ ( .A(\us32\/_0010_ ), .B(\w3\[2\] ), .X(_0500_ ) );
sky130_fd_sc_hd__xor2_1 _3095_ ( .A(\us32\/_0011_ ), .B(\w3\[3\] ), .X(_0501_ ) );
sky130_fd_sc_hd__xor2_1 _3096_ ( .A(\us32\/_0012_ ), .B(\w3\[4\] ), .X(_0502_ ) );
sky130_fd_sc_hd__xor2_1 _3097_ ( .A(\us32\/_0013_ ), .B(\w3\[5\] ), .X(_0503_ ) );
sky130_fd_sc_hd__xor2_1 _3098_ ( .A(\us32\/_0014_ ), .B(\w3\[6\] ), .X(_0504_ ) );
sky130_fd_sc_hd__xor2_1 _3099_ ( .A(\us32\/_0015_ ), .B(\w3\[7\] ), .X(_0505_ ) );
sky130_fd_sc_hd__conb_1 _34 ( .HI( ), .LO(net34 ) );
sky130_fd_sc_hd__clkbuf_1 _3495_ ( .A(\us11\/_0015_ ), .X(_1379_ ) );
sky130_fd_sc_hd__conb_1 _34_35 ( .HI( ), .LO(net35 ) );
sky130_fd_sc_hd__conb_1 _34_36 ( .HI( ), .LO(net36 ) );
sky130_fd_sc_hd__conb_1 _34_37 ( .HI( ), .LO(net37 ) );
sky130_fd_sc_hd__conb_1 _34_38 ( .HI( ), .LO(net38 ) );
sky130_fd_sc_hd__conb_1 _34_39 ( .HI( ), .LO(net39 ) );
sky130_fd_sc_hd__conb_1 _34_40 ( .HI( ), .LO(net40 ) );
sky130_fd_sc_hd__conb_1 _34_41 ( .HI( ), .LO(net41 ) );
sky130_fd_sc_hd__conb_1 _34_42 ( .HI( ), .LO(net42 ) );
sky130_fd_sc_hd__conb_1 _34_43 ( .HI( ), .LO(net43 ) );
sky130_fd_sc_hd__conb_1 _34_44 ( .HI( ), .LO(net44 ) );
sky130_fd_sc_hd__conb_1 _34_45 ( .HI( ), .LO(net45 ) );
sky130_fd_sc_hd__conb_1 _34_46 ( .HI( ), .LO(net46 ) );
sky130_fd_sc_hd__conb_1 _34_47 ( .HI( ), .LO(net47 ) );
sky130_fd_sc_hd__conb_1 _34_48 ( .HI( ), .LO(net48 ) );
sky130_fd_sc_hd__clkbuf_1 _3504_ ( .A(\us11\/_0009_ ), .X(_1373_ ) );
sky130_fd_sc_hd__clkbuf_1 _3528_ ( .A(\us11\/_0013_ ), .X(_1377_ ) );
sky130_fd_sc_hd__clkbuf_1 _3592_ ( .A(\us13\/_0015_ ), .X(_1419_ ) );
sky130_fd_sc_hd__clkbuf_1 _3636_ ( .A(\us20\/_0015_ ), .X(_1451_ ) );
sky130_fd_sc_hd__clkbuf_1 _3640_ ( .A(\us10\/_0015_ ), .X(_1387_ ) );
sky130_fd_sc_hd__clkbuf_1 _3887_ ( .A(_0425_ ), .X(_0164_ ) );
sky130_fd_sc_hd__dfxtp_1 _4008_ ( .D(_0261_ ), .Q(\dcnt\[0\] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_1 _4009_ ( .D(_0262_ ), .Q(\dcnt\[1\] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_1 _4010_ ( .D(_0263_ ), .Q(\dcnt\[2\] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_1 _4011_ ( .D(_0264_ ), .Q(\dcnt\[3\] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_1 _4012_ ( .D(_0265_ ), .Q(done ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4013_ ( .D(_0266_ ), .Q(\text_in_r\[0\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4014_ ( .D(_0305_ ), .Q(\text_in_r\[1\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4015_ ( .D(_0316_ ), .Q(\text_in_r\[2\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4016_ ( .D(_0327_ ), .Q(\text_in_r\[3\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4017_ ( .D(_0338_ ), .Q(\text_in_r\[4\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4018_ ( .D(_0349_ ), .Q(\text_in_r\[5\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4019_ ( .D(_0360_ ), .Q(\text_in_r\[6\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4020_ ( .D(_0371_ ), .Q(\text_in_r\[7\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4021_ ( .D(_0382_ ), .Q(\text_in_r\[8\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4022_ ( .D(_0393_ ), .Q(\text_in_r\[9\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4023_ ( .D(_0277_ ), .Q(\text_in_r\[10\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4024_ ( .D(_0288_ ), .Q(\text_in_r\[11\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4025_ ( .D(_0297_ ), .Q(\text_in_r\[12\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4026_ ( .D(_0298_ ), .Q(\text_in_r\[13\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4027_ ( .D(_0299_ ), .Q(\text_in_r\[14\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4028_ ( .D(_0300_ ), .Q(\text_in_r\[15\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4029_ ( .D(_0301_ ), .Q(\text_in_r\[16\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4030_ ( .D(_0302_ ), .Q(\text_in_r\[17\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4031_ ( .D(_0303_ ), .Q(\text_in_r\[18\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4032_ ( .D(_0304_ ), .Q(\text_in_r\[19\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4033_ ( .D(_0306_ ), .Q(\text_in_r\[20\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4034_ ( .D(_0307_ ), .Q(\text_in_r\[21\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4035_ ( .D(_0308_ ), .Q(\text_in_r\[22\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4036_ ( .D(_0309_ ), .Q(\text_in_r\[23\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4037_ ( .D(_0310_ ), .Q(\text_in_r\[24\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4038_ ( .D(_0311_ ), .Q(\text_in_r\[25\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4039_ ( .D(_0312_ ), .Q(\text_in_r\[26\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4040_ ( .D(_0313_ ), .Q(\text_in_r\[27\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4041_ ( .D(_0314_ ), .Q(\text_in_r\[28\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4042_ ( .D(_0315_ ), .Q(\text_in_r\[29\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4043_ ( .D(_0317_ ), .Q(\text_in_r\[30\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4044_ ( .D(_0318_ ), .Q(\text_in_r\[31\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4045_ ( .D(_0319_ ), .Q(\text_in_r\[32\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4046_ ( .D(_0320_ ), .Q(\text_in_r\[33\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4047_ ( .D(_0321_ ), .Q(\text_in_r\[34\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4048_ ( .D(_0322_ ), .Q(\text_in_r\[35\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4049_ ( .D(_0323_ ), .Q(\text_in_r\[36\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4050_ ( .D(_0324_ ), .Q(\text_in_r\[37\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4051_ ( .D(_0325_ ), .Q(\text_in_r\[38\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4052_ ( .D(_0326_ ), .Q(\text_in_r\[39\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4053_ ( .D(_0328_ ), .Q(\text_in_r\[40\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4054_ ( .D(_0329_ ), .Q(\text_in_r\[41\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4055_ ( .D(_0330_ ), .Q(\text_in_r\[42\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4056_ ( .D(_0331_ ), .Q(\text_in_r\[43\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4057_ ( .D(_0332_ ), .Q(\text_in_r\[44\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4058_ ( .D(_0333_ ), .Q(\text_in_r\[45\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4059_ ( .D(_0334_ ), .Q(\text_in_r\[46\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4060_ ( .D(_0335_ ), .Q(\text_in_r\[47\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4061_ ( .D(_0336_ ), .Q(\text_in_r\[48\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4062_ ( .D(_0337_ ), .Q(\text_in_r\[49\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4063_ ( .D(_0339_ ), .Q(\text_in_r\[50\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4064_ ( .D(_0340_ ), .Q(\text_in_r\[51\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4065_ ( .D(_0341_ ), .Q(\text_in_r\[52\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4066_ ( .D(_0342_ ), .Q(\text_in_r\[53\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4067_ ( .D(_0343_ ), .Q(\text_in_r\[54\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4068_ ( .D(_0344_ ), .Q(\text_in_r\[55\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4069_ ( .D(_0345_ ), .Q(\text_in_r\[56\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4070_ ( .D(_0346_ ), .Q(\text_in_r\[57\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4071_ ( .D(_0347_ ), .Q(\text_in_r\[58\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4072_ ( .D(_0348_ ), .Q(\text_in_r\[59\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4073_ ( .D(_0350_ ), .Q(\text_in_r\[60\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4074_ ( .D(_0351_ ), .Q(\text_in_r\[61\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4075_ ( .D(_0352_ ), .Q(\text_in_r\[62\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4076_ ( .D(_0353_ ), .Q(\text_in_r\[63\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4077_ ( .D(_0354_ ), .Q(\text_in_r\[64\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4078_ ( .D(_0355_ ), .Q(\text_in_r\[65\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4079_ ( .D(_0356_ ), .Q(\text_in_r\[66\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4080_ ( .D(_0357_ ), .Q(\text_in_r\[67\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4081_ ( .D(_0358_ ), .Q(\text_in_r\[68\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4082_ ( .D(_0359_ ), .Q(\text_in_r\[69\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4083_ ( .D(_0361_ ), .Q(\text_in_r\[70\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4084_ ( .D(_0362_ ), .Q(\text_in_r\[71\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4085_ ( .D(_0363_ ), .Q(\text_in_r\[72\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4086_ ( .D(_0364_ ), .Q(\text_in_r\[73\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4087_ ( .D(_0365_ ), .Q(\text_in_r\[74\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4088_ ( .D(_0366_ ), .Q(\text_in_r\[75\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4089_ ( .D(_0367_ ), .Q(\text_in_r\[76\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4090_ ( .D(_0368_ ), .Q(\text_in_r\[77\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4091_ ( .D(_0369_ ), .Q(\text_in_r\[78\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4092_ ( .D(_0370_ ), .Q(\text_in_r\[79\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4093_ ( .D(_0372_ ), .Q(\text_in_r\[80\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4094_ ( .D(_0373_ ), .Q(\text_in_r\[81\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4095_ ( .D(_0374_ ), .Q(\text_in_r\[82\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4096_ ( .D(_0375_ ), .Q(\text_in_r\[83\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4097_ ( .D(_0376_ ), .Q(\text_in_r\[84\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4098_ ( .D(_0377_ ), .Q(\text_in_r\[85\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4099_ ( .D(_0378_ ), .Q(\text_in_r\[86\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4100_ ( .D(_0379_ ), .Q(\text_in_r\[87\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4101_ ( .D(_0380_ ), .Q(\text_in_r\[88\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4102_ ( .D(_0381_ ), .Q(\text_in_r\[89\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4103_ ( .D(_0383_ ), .Q(\text_in_r\[90\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4104_ ( .D(_0384_ ), .Q(\text_in_r\[91\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4105_ ( .D(_0385_ ), .Q(\text_in_r\[92\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4106_ ( .D(_0386_ ), .Q(\text_in_r\[93\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4107_ ( .D(_0387_ ), .Q(\text_in_r\[94\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4108_ ( .D(_0388_ ), .Q(\text_in_r\[95\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4109_ ( .D(_0389_ ), .Q(\text_in_r\[96\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4110_ ( .D(_0390_ ), .Q(\text_in_r\[97\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4111_ ( .D(_0391_ ), .Q(\text_in_r\[98\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4112_ ( .D(_0392_ ), .Q(\text_in_r\[99\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4113_ ( .D(_0267_ ), .Q(\text_in_r\[100\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4114_ ( .D(_0268_ ), .Q(\text_in_r\[101\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4115_ ( .D(_0269_ ), .Q(\text_in_r\[102\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4116_ ( .D(_0270_ ), .Q(\text_in_r\[103\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4117_ ( .D(_0271_ ), .Q(\text_in_r\[104\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4118_ ( .D(_0272_ ), .Q(\text_in_r\[105\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4119_ ( .D(_0273_ ), .Q(\text_in_r\[106\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4120_ ( .D(_0274_ ), .Q(\text_in_r\[107\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4121_ ( .D(_0275_ ), .Q(\text_in_r\[108\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4122_ ( .D(_0276_ ), .Q(\text_in_r\[109\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4123_ ( .D(_0278_ ), .Q(\text_in_r\[110\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4124_ ( .D(_0279_ ), .Q(\text_in_r\[111\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4125_ ( .D(_0280_ ), .Q(\text_in_r\[112\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4126_ ( .D(_0281_ ), .Q(\text_in_r\[113\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4127_ ( .D(_0282_ ), .Q(\text_in_r\[114\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4128_ ( .D(_0283_ ), .Q(\text_in_r\[115\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4129_ ( .D(_0284_ ), .Q(\text_in_r\[116\] ), .CLK(CTS_5 ) );
sky130_fd_sc_hd__dfxtp_1 _4130_ ( .D(_0285_ ), .Q(\text_in_r\[117\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4131_ ( .D(_0286_ ), .Q(\text_in_r\[118\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4132_ ( .D(_0287_ ), .Q(\text_in_r\[119\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4133_ ( .D(_0289_ ), .Q(\text_in_r\[120\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4134_ ( .D(_0290_ ), .Q(\text_in_r\[121\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4135_ ( .D(_0291_ ), .Q(\text_in_r\[122\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4136_ ( .D(_0292_ ), .Q(\text_in_r\[123\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4137_ ( .D(_0293_ ), .Q(\text_in_r\[124\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4138_ ( .D(_0294_ ), .Q(\text_in_r\[125\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4139_ ( .D(_0295_ ), .Q(\text_in_r\[126\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4140_ ( .D(_0296_ ), .Q(\text_in_r\[127\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4141_ ( .D(ld ), .Q(ld_r ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4142_ ( .D(_1548_ ), .Q(\sa33\[0\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4143_ ( .D(_1549_ ), .Q(\sa33\[1\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4144_ ( .D(_1550_ ), .Q(\sa33\[2\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4145_ ( .D(_1551_ ), .Q(\sa33\[3\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4146_ ( .D(_1552_ ), .Q(\sa33\[4\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4147_ ( .D(_1553_ ), .Q(\sa33\[5\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4148_ ( .D(_1554_ ), .Q(\sa33\[6\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4149_ ( .D(_1555_ ), .Q(\sa33\[7\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4150_ ( .D(_1484_ ), .Q(\sa23\[0\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4151_ ( .D(_1485_ ), .Q(\sa23\[1\] ), .CLK(CTS_11 ) );
sky130_fd_sc_hd__dfxtp_1 _4152_ ( .D(_1486_ ), .Q(\sa23\[2\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4153_ ( .D(_1487_ ), .Q(\sa23\[3\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4154_ ( .D(_1488_ ), .Q(\sa23\[4\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4155_ ( .D(_1489_ ), .Q(\sa23\[5\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4156_ ( .D(_1490_ ), .Q(\sa23\[6\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4157_ ( .D(_1491_ ), .Q(\sa23\[7\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4158_ ( .D(_1420_ ), .Q(\sa13\[0\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4159_ ( .D(_1421_ ), .Q(\sa13\[1\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4160_ ( .D(_1422_ ), .Q(\sa13\[2\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4161_ ( .D(_1423_ ), .Q(\sa13\[3\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4162_ ( .D(_1424_ ), .Q(\sa13\[4\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4163_ ( .D(_1425_ ), .Q(\sa13\[5\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4164_ ( .D(_1426_ ), .Q(\sa13\[6\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4165_ ( .D(_1427_ ), .Q(\sa13\[7\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4166_ ( .D(_1348_ ), .Q(\sa03\[0\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4167_ ( .D(_1349_ ), .Q(\sa03\[1\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4168_ ( .D(_1350_ ), .Q(\sa03\[2\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4169_ ( .D(_1351_ ), .Q(\sa03\[3\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4170_ ( .D(_1352_ ), .Q(\sa03\[4\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4171_ ( .D(_1353_ ), .Q(\sa03\[5\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4172_ ( .D(_1354_ ), .Q(\sa03\[6\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4173_ ( .D(_1355_ ), .Q(\sa03\[7\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4174_ ( .D(_1532_ ), .Q(\sa32\[0\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4175_ ( .D(_1533_ ), .Q(\sa32\[1\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4176_ ( .D(_1534_ ), .Q(\sa32\[2\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4177_ ( .D(_1535_ ), .Q(\sa32\[3\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4178_ ( .D(_1536_ ), .Q(\sa32\[4\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4179_ ( .D(_1537_ ), .Q(\sa32\[5\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4180_ ( .D(_1538_ ), .Q(\sa32\[6\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4181_ ( .D(_1539_ ), .Q(\sa32\[7\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4182_ ( .D(_1476_ ), .Q(\sa22\[0\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4183_ ( .D(_1477_ ), .Q(\sa22\[1\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4184_ ( .D(_1478_ ), .Q(\sa22\[2\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4185_ ( .D(_1479_ ), .Q(\sa22\[3\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4186_ ( .D(_1480_ ), .Q(\sa22\[4\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4187_ ( .D(_1481_ ), .Q(\sa22\[5\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4188_ ( .D(_1482_ ), .Q(\sa22\[6\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4189_ ( .D(_1483_ ), .Q(\sa22\[7\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4190_ ( .D(_1404_ ), .Q(\sa12\[0\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4191_ ( .D(_1405_ ), .Q(\sa12\[1\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4192_ ( .D(_1406_ ), .Q(\sa12\[2\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4193_ ( .D(_1407_ ), .Q(\sa12\[3\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4194_ ( .D(_1408_ ), .Q(\sa12\[4\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4195_ ( .D(_1409_ ), .Q(\sa12\[5\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4196_ ( .D(_1410_ ), .Q(\sa12\[6\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4197_ ( .D(_1411_ ), .Q(\sa12\[7\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4198_ ( .D(_1332_ ), .Q(\sa02\[0\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4199_ ( .D(_1333_ ), .Q(\sa02\[1\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4200_ ( .D(_1334_ ), .Q(\sa02\[2\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4201_ ( .D(_1335_ ), .Q(\sa02\[3\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4202_ ( .D(_1336_ ), .Q(\sa02\[4\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4203_ ( .D(_1337_ ), .Q(\sa02\[5\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4204_ ( .D(_1338_ ), .Q(\sa02\[6\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4205_ ( .D(_1339_ ), .Q(\sa02\[7\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4206_ ( .D(_1516_ ), .Q(\sa31\[0\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4207_ ( .D(_1517_ ), .Q(\sa31\[1\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4208_ ( .D(_1518_ ), .Q(\sa31\[2\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4209_ ( .D(_1519_ ), .Q(\sa31\[3\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4210_ ( .D(_1520_ ), .Q(\sa31\[4\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4211_ ( .D(_1521_ ), .Q(\sa31\[5\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4212_ ( .D(_1522_ ), .Q(\sa31\[6\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4213_ ( .D(_1523_ ), .Q(\sa31\[7\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4214_ ( .D(_1452_ ), .Q(\sa21\[0\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4215_ ( .D(_1453_ ), .Q(\sa21\[1\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4216_ ( .D(_1454_ ), .Q(\sa21\[2\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4217_ ( .D(_1455_ ), .Q(\sa21\[3\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4218_ ( .D(_1456_ ), .Q(\sa21\[4\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4219_ ( .D(_1457_ ), .Q(\sa21\[5\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4220_ ( .D(_1458_ ), .Q(\sa21\[6\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4221_ ( .D(_1459_ ), .Q(\sa21\[7\] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4222_ ( .D(_1388_ ), .Q(\sa11\[0\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4223_ ( .D(_1389_ ), .Q(\sa11\[1\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4224_ ( .D(_1390_ ), .Q(\sa11\[2\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4225_ ( .D(_1391_ ), .Q(\sa11\[3\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4226_ ( .D(_1392_ ), .Q(\sa11\[4\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4227_ ( .D(_1393_ ), .Q(\sa11\[5\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4228_ ( .D(_1394_ ), .Q(\sa11\[6\] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4229_ ( .D(_1395_ ), .Q(\sa11\[7\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4230_ ( .D(_1316_ ), .Q(\sa01\[0\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4231_ ( .D(_1317_ ), .Q(\sa01\[1\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4232_ ( .D(_1318_ ), .Q(\sa01\[2\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4233_ ( .D(_1319_ ), .Q(\sa01\[3\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4234_ ( .D(_1320_ ), .Q(\sa01\[4\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4235_ ( .D(_1321_ ), .Q(\sa01\[5\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4236_ ( .D(_1322_ ), .Q(\sa01\[6\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4237_ ( .D(_1323_ ), .Q(\sa01\[7\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4238_ ( .D(_1492_ ), .Q(\sa30\[0\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4239_ ( .D(_1493_ ), .Q(\sa30\[1\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4240_ ( .D(_1494_ ), .Q(\sa30\[2\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4241_ ( .D(_1495_ ), .Q(\sa30\[3\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4242_ ( .D(_1496_ ), .Q(\sa30\[4\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4243_ ( .D(_1497_ ), .Q(\sa30\[5\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4244_ ( .D(_1498_ ), .Q(\sa30\[6\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4245_ ( .D(_1499_ ), .Q(\sa30\[7\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4246_ ( .D(_1428_ ), .Q(\sa20\[0\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4247_ ( .D(_1429_ ), .Q(\sa20\[1\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4248_ ( .D(_1430_ ), .Q(\sa20\[2\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4249_ ( .D(_1431_ ), .Q(\sa20\[3\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4250_ ( .D(_1432_ ), .Q(\sa20\[4\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4251_ ( .D(_1433_ ), .Q(\sa20\[5\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4252_ ( .D(_1434_ ), .Q(\sa20\[6\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4253_ ( .D(_1435_ ), .Q(\sa20\[7\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4254_ ( .D(_1364_ ), .Q(\sa10\[0\] ), .CLK(CTS_5 ) );
sky130_fd_sc_hd__dfxtp_1 _4255_ ( .D(_1365_ ), .Q(\sa10\[1\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4256_ ( .D(_1366_ ), .Q(\sa10\[2\] ), .CLK(CTS_5 ) );
sky130_fd_sc_hd__dfxtp_1 _4257_ ( .D(_1367_ ), .Q(\sa10\[3\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4258_ ( .D(_1368_ ), .Q(\sa10\[4\] ), .CLK(CTS_5 ) );
sky130_fd_sc_hd__dfxtp_1 _4259_ ( .D(_1369_ ), .Q(\sa10\[5\] ), .CLK(CTS_5 ) );
sky130_fd_sc_hd__dfxtp_1 _4260_ ( .D(_1370_ ), .Q(\sa10\[6\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4261_ ( .D(_1371_ ), .Q(\sa10\[7\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4262_ ( .D(_1300_ ), .Q(\sa00\[0\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4263_ ( .D(_1301_ ), .Q(\sa00\[1\] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_1 _4264_ ( .D(_1302_ ), .Q(\sa00\[2\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4265_ ( .D(_1303_ ), .Q(\sa00\[3\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4266_ ( .D(_1304_ ), .Q(\sa00\[4\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4267_ ( .D(_1305_ ), .Q(\sa00\[5\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4268_ ( .D(_1306_ ), .Q(\sa00\[6\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4269_ ( .D(_1307_ ), .Q(\sa00\[7\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4270_ ( .D(_0418_ ), .Q(\text_out[120] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4271_ ( .D(_0419_ ), .Q(\text_out[121] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_1 _4272_ ( .D(_0420_ ), .Q(\text_out[122] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4273_ ( .D(_0421_ ), .Q(\text_out[123] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4274_ ( .D(_0422_ ), .Q(\text_out[124] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_2 _4275_ ( .D(_0423_ ), .Q(\text_out[125] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4276_ ( .D(_0424_ ), .Q(\text_out[126] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4277_ ( .D(_0164_ ), .Q(\text_out[127] ), .CLK(CTS_5 ) );
sky130_fd_sc_hd__dfxtp_1 _4278_ ( .D(_0514_ ), .Q(\text_out[88] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4279_ ( .D(_0515_ ), .Q(\text_out[89] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4280_ ( .D(_0516_ ), .Q(\text_out[90] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4281_ ( .D(_0517_ ), .Q(\text_out[91] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4282_ ( .D(_0518_ ), .Q(\text_out[92] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4283_ ( .D(_0519_ ), .Q(\text_out[93] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4284_ ( .D(_0520_ ), .Q(\text_out[94] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4285_ ( .D(_0521_ ), .Q(\text_out[95] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4286_ ( .D(_0474_ ), .Q(\text_out[56] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4287_ ( .D(_0475_ ), .Q(\text_out[57] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4288_ ( .D(_0476_ ), .Q(\text_out[58] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4289_ ( .D(_0477_ ), .Q(\text_out[59] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4290_ ( .D(_0478_ ), .Q(\text_out[60] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4291_ ( .D(_0479_ ), .Q(\text_out[61] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4292_ ( .D(_0480_ ), .Q(\text_out[62] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4293_ ( .D(_0481_ ), .Q(\text_out[63] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4294_ ( .D(_0442_ ), .Q(\text_out[24] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4295_ ( .D(_0443_ ), .Q(\text_out[25] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4296_ ( .D(_0444_ ), .Q(\text_out[26] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4297_ ( .D(_0445_ ), .Q(\text_out[27] ), .CLK(CTS_11 ) );
sky130_fd_sc_hd__dfxtp_1 _4298_ ( .D(_0446_ ), .Q(\text_out[28] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4299_ ( .D(_0447_ ), .Q(\text_out[29] ), .CLK(CTS_11 ) );
sky130_fd_sc_hd__dfxtp_1 _4300_ ( .D(_0448_ ), .Q(\text_out[30] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4301_ ( .D(_0449_ ), .Q(\text_out[31] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4302_ ( .D(_0410_ ), .Q(\text_out[112] ), .CLK(CTS_5 ) );
sky130_fd_sc_hd__dfxtp_1 _4303_ ( .D(_0411_ ), .Q(\text_out[113] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4304_ ( .D(_0412_ ), .Q(\text_out[114] ), .CLK(CTS_5 ) );
sky130_fd_sc_hd__dfxtp_1 _4305_ ( .D(_0413_ ), .Q(\text_out[115] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4306_ ( .D(_0414_ ), .Q(\text_out[116] ), .CLK(CTS_5 ) );
sky130_fd_sc_hd__dfxtp_1 _4307_ ( .D(_0415_ ), .Q(\text_out[117] ), .CLK(CTS_5 ) );
sky130_fd_sc_hd__dfxtp_1 _4308_ ( .D(_0416_ ), .Q(\text_out[118] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4309_ ( .D(_0417_ ), .Q(\text_out[119] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4310_ ( .D(_0506_ ), .Q(FE_OFN0_text_out_80 ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4311_ ( .D(_0507_ ), .Q(\text_out[81] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4312_ ( .D(_0508_ ), .Q(\text_out[82] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4313_ ( .D(_0509_ ), .Q(\text_out[83] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4314_ ( .D(_0510_ ), .Q(\text_out[84] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4315_ ( .D(_0511_ ), .Q(\text_out[85] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4316_ ( .D(_0512_ ), .Q(\text_out[86] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_2 _4317_ ( .D(_0513_ ), .Q(\text_out[87] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4318_ ( .D(_0466_ ), .Q(\text_out[48] ), .CLK(CTS_5 ) );
sky130_fd_sc_hd__dfxtp_2 _4319_ ( .D(_0467_ ), .Q(\text_out[49] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4320_ ( .D(_0468_ ), .Q(\text_out[50] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4321_ ( .D(_0469_ ), .Q(\text_out[51] ), .CLK(CTS_11 ) );
sky130_fd_sc_hd__dfxtp_1 _4322_ ( .D(_0470_ ), .Q(\text_out[52] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4323_ ( .D(_0471_ ), .Q(\text_out[53] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4324_ ( .D(_0472_ ), .Q(\text_out[54] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4325_ ( .D(_0473_ ), .Q(\text_out[55] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4326_ ( .D(_0434_ ), .Q(\text_out[16] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4327_ ( .D(_0435_ ), .Q(\text_out[17] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_2 _4328_ ( .D(_0436_ ), .Q(\text_out[18] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4329_ ( .D(_0437_ ), .Q(\text_out[19] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4330_ ( .D(_0438_ ), .Q(\text_out[20] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4331_ ( .D(_0439_ ), .Q(\text_out[21] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4332_ ( .D(_0440_ ), .Q(\text_out[22] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4333_ ( .D(_0441_ ), .Q(\text_out[23] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4334_ ( .D(_0402_ ), .Q(\text_out[104] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_1 _4335_ ( .D(_0403_ ), .Q(\text_out[105] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_1 _4336_ ( .D(_0404_ ), .Q(\text_out[106] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4337_ ( .D(_0405_ ), .Q(\text_out[107] ), .CLK(CTS_11 ) );
sky130_fd_sc_hd__dfxtp_1 _4338_ ( .D(_0406_ ), .Q(\text_out[108] ), .CLK(CTS_5 ) );
sky130_fd_sc_hd__dfxtp_1 _4339_ ( .D(_0407_ ), .Q(\text_out[109] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_1 _4340_ ( .D(_0408_ ), .Q(\text_out[110] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4341_ ( .D(_0409_ ), .Q(\text_out[111] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_1 _4342_ ( .D(_0490_ ), .Q(\text_out[72] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4343_ ( .D(_0491_ ), .Q(\text_out[73] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 _4344_ ( .D(_0492_ ), .Q(\text_out[74] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4345_ ( .D(_0493_ ), .Q(\text_out[75] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4346_ ( .D(_0494_ ), .Q(\text_out[76] ), .CLK(CTS_11 ) );
sky130_fd_sc_hd__dfxtp_1 _4347_ ( .D(_0495_ ), .Q(\text_out[77] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4348_ ( .D(_0496_ ), .Q(\text_out[78] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4349_ ( .D(_0497_ ), .Q(\text_out[79] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4350_ ( .D(_0458_ ), .Q(\text_out[40] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4351_ ( .D(_0459_ ), .Q(\text_out[41] ), .CLK(CTS_11 ) );
sky130_fd_sc_hd__dfxtp_1 _4352_ ( .D(_0460_ ), .Q(\text_out[42] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4353_ ( .D(_0461_ ), .Q(\text_out[43] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4354_ ( .D(_0462_ ), .Q(\text_out[44] ), .CLK(CTS_5 ) );
sky130_fd_sc_hd__dfxtp_2 _4355_ ( .D(_0463_ ), .Q(\text_out[45] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 _4356_ ( .D(_0464_ ), .Q(\text_out[46] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4357_ ( .D(_0465_ ), .Q(\text_out[47] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4358_ ( .D(_0426_ ), .Q(\text_out[8] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4359_ ( .D(_0427_ ), .Q(\text_out[9] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4360_ ( .D(_0428_ ), .Q(\text_out[10] ), .CLK(CTS_11 ) );
sky130_fd_sc_hd__dfxtp_1 _4361_ ( .D(_0429_ ), .Q(\text_out[11] ), .CLK(CTS_11 ) );
sky130_fd_sc_hd__dfxtp_1 _4362_ ( .D(_0430_ ), .Q(\text_out[12] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4363_ ( .D(_0431_ ), .Q(\text_out[13] ), .CLK(CTS_11 ) );
sky130_fd_sc_hd__dfxtp_1 _4364_ ( .D(_0432_ ), .Q(\text_out[14] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 _4365_ ( .D(_0433_ ), .Q(\text_out[15] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4366_ ( .D(_0394_ ), .Q(\text_out[96] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_1 _4367_ ( .D(_0395_ ), .Q(\text_out[97] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4368_ ( .D(_0396_ ), .Q(\text_out[98] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4369_ ( .D(_0397_ ), .Q(\text_out[99] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4370_ ( .D(_0398_ ), .Q(\text_out[100] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4371_ ( .D(_0399_ ), .Q(\text_out[101] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_1 _4372_ ( .D(_0400_ ), .Q(\text_out[102] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4373_ ( .D(_0401_ ), .Q(\text_out[103] ), .CLK(CTS_5 ) );
sky130_fd_sc_hd__dfxtp_1 _4374_ ( .D(_0482_ ), .Q(\text_out[64] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4375_ ( .D(_0483_ ), .Q(\text_out[65] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4376_ ( .D(_0484_ ), .Q(\text_out[66] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 _4377_ ( .D(_0485_ ), .Q(\text_out[67] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_2 _4378_ ( .D(_0486_ ), .Q(\text_out[68] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_2 _4379_ ( .D(_0487_ ), .Q(\text_out[69] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_2 _4380_ ( .D(_0488_ ), .Q(\text_out[70] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4381_ ( .D(_0489_ ), .Q(\text_out[71] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4382_ ( .D(_0450_ ), .Q(\text_out[32] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4383_ ( .D(_0451_ ), .Q(\text_out[33] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 _4384_ ( .D(_0452_ ), .Q(\text_out[34] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_2 _4385_ ( .D(_0453_ ), .Q(\text_out[35] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 _4386_ ( .D(_0454_ ), .Q(\text_out[36] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_1 _4387_ ( .D(_0455_ ), .Q(\text_out[37] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4388_ ( .D(_0456_ ), .Q(\text_out[38] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_1 _4389_ ( .D(_0457_ ), .Q(\text_out[39] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4390_ ( .D(_0498_ ), .Q(\text_out[0] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_1 _4391_ ( .D(_0499_ ), .Q(\text_out[1] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 _4392_ ( .D(_0500_ ), .Q(\text_out[2] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 _4393_ ( .D(_0501_ ), .Q(\text_out[3] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 _4394_ ( .D(_0502_ ), .Q(\text_out[4] ), .CLK(CTS_18 ) );
sky130_fd_sc_hd__dfxtp_1 _4395_ ( .D(_0503_ ), .Q(\text_out[5] ), .CLK(CTS_12 ) );
sky130_fd_sc_hd__dfxtp_1 _4396_ ( .D(_0504_ ), .Q(\text_out[6] ), .CLK(CTS_8 ) );
sky130_fd_sc_hd__dfxtp_1 _4397_ ( .D(_0505_ ), .Q(\text_out[7] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__xor2_1 \u0/_0850_ ( .A(\u0\/u3\/_0008_ ), .B(\w0\[0\] ), .X(\u0\/_0385_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0851_ ( .A(\u0\/rcon\[0\] ), .B(\u0\/_0385_ ), .X(\u0\/_0386_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/_0852_ ( .A(ld ), .X(\u0\/_0387_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/_0853_ ( .A(\u0\/_0387_ ), .X(\u0\/_0388_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0854_ ( .A0(\u0\/_0386_ ), .A1(\key[96] ), .S(\u0\/_0388_ ), .X(\u0\/_0128_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0855_ ( .A(\u0\/u3\/_0009_ ), .B(\w0\[1\] ), .X(\u0\/_0389_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0856_ ( .A(\u0\/rcon\[1\] ), .B(\u0\/_0389_ ), .X(\u0\/_0390_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0857_ ( .A0(\u0\/_0390_ ), .A1(\key[97] ), .S(\u0\/_0388_ ), .X(\u0\/_0139_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0858_ ( .A(\u0\/u3\/_0010_ ), .B(\w0\[2\] ), .X(\u0\/_0391_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0859_ ( .A(\u0\/rcon\[2\] ), .B(\u0\/_0391_ ), .X(\u0\/_0392_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0860_ ( .A0(\u0\/_0392_ ), .A1(\key[98] ), .S(\u0\/_0388_ ), .X(\u0\/_0150_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0861_ ( .A(\u0\/u3\/_0011_ ), .B(\w0\[3\] ), .X(\u0\/_0393_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0862_ ( .A(\u0\/rcon\[3\] ), .B(\u0\/_0393_ ), .X(\u0\/_0394_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0863_ ( .A0(\u0\/_0394_ ), .A1(\key[99] ), .S(\u0\/_0388_ ), .X(\u0\/_0153_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0864_ ( .A(\u0\/u3\/_0012_ ), .B(\w0\[4\] ), .X(\u0\/_0395_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0865_ ( .A(\u0\/rcon\[4\] ), .B(\u0\/_0395_ ), .X(\u0\/_0396_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0866_ ( .A0(\u0\/_0396_ ), .A1(\key[100] ), .S(\u0\/_0388_ ), .X(\u0\/_0154_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0867_ ( .A(\u0\/u3\/_0013_ ), .B(\w0\[5\] ), .X(\u0\/_0397_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0868_ ( .A(\u0\/rcon\[5\] ), .B(\u0\/_0397_ ), .X(\u0\/_0398_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0869_ ( .A0(\u0\/_0398_ ), .A1(\key[101] ), .S(\u0\/_0388_ ), .X(\u0\/_0155_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0870_ ( .A(\u0\/u3\/_0014_ ), .B(\w0\[6\] ), .X(\u0\/_0399_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0871_ ( .A(\u0\/rcon\[6\] ), .B(\u0\/_0399_ ), .X(\u0\/_0400_ ) );
sky130_fd_sc_hd__buf_2 \u0/_0872_ ( .A(\u0\/_0387_ ), .X(\u0\/_0401_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0873_ ( .A0(\u0\/_0400_ ), .A1(\key[102] ), .S(\u0\/_0401_ ), .X(\u0\/_0156_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0874_ ( .A(\u0\/u3\/_0015_ ), .B(\w0\[7\] ), .X(\u0\/_0402_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0875_ ( .A(\u0\/rcon\[7\] ), .B(\u0\/_0402_ ), .X(\u0\/_0403_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0876_ ( .A0(\u0\/_0403_ ), .A1(\key[103] ), .S(\u0\/_0401_ ), .X(\u0\/_0157_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0877_ ( .A(\u0\/u2\/_0008_ ), .B(\w0\[8\] ), .X(\u0\/_0404_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0878_ ( .A(\u0\/rcon\[8\] ), .B(\u0\/_0404_ ), .X(\u0\/_0405_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0879_ ( .A0(\u0\/_0405_ ), .A1(\key[104] ), .S(\u0\/_0401_ ), .X(\u0\/_0158_ ) );
sky130_fd_sc_hd__xor2_2 \u0/_0880_ ( .A(\u0\/u2\/_0009_ ), .B(\w0\[9\] ), .X(\u0\/_0406_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0881_ ( .A(\u0\/rcon\[9\] ), .B(\u0\/_0406_ ), .X(\u0\/_0407_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0882_ ( .A0(\u0\/_0407_ ), .A1(\key[105] ), .S(\u0\/_0401_ ), .X(\u0\/_0159_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0883_ ( .A(\u0\/u2\/_0010_ ), .B(\w0\[10\] ), .X(\u0\/_0408_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0884_ ( .A(\u0\/rcon\[10\] ), .B(\u0\/_0408_ ), .X(\u0\/_0409_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0885_ ( .A0(\u0\/_0409_ ), .A1(\key[106] ), .S(\u0\/_0401_ ), .X(\u0\/_0129_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0886_ ( .A(\u0\/u2\/_0011_ ), .B(\w0\[11\] ), .X(\u0\/_0410_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0887_ ( .A(\u0\/rcon\[11\] ), .B(\u0\/_0410_ ), .X(\u0\/_0411_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0888_ ( .A0(\u0\/_0411_ ), .A1(\key[107] ), .S(\u0\/_0401_ ), .X(\u0\/_0130_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0889_ ( .A(\u0\/u2\/_0012_ ), .B(\w0\[12\] ), .X(\u0\/_0412_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0890_ ( .A(\u0\/rcon\[12\] ), .B(\u0\/_0412_ ), .X(\u0\/_0413_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0891_ ( .A0(\u0\/_0413_ ), .A1(\key[108] ), .S(\u0\/_0401_ ), .X(\u0\/_0131_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0892_ ( .A(\u0\/u2\/_0013_ ), .B(\w0\[13\] ), .X(\u0\/_0414_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0893_ ( .A(\u0\/rcon\[13\] ), .B(\u0\/_0414_ ), .X(\u0\/_0415_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0894_ ( .A0(\u0\/_0415_ ), .A1(\key[109] ), .S(\u0\/_0401_ ), .X(\u0\/_0132_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0895_ ( .A(\u0\/u2\/_0014_ ), .B(\w0\[14\] ), .X(\u0\/_0416_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0896_ ( .A(\u0\/rcon\[14\] ), .B(\u0\/_0416_ ), .X(\u0\/_0417_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0897_ ( .A0(\u0\/_0417_ ), .A1(\key[110] ), .S(\u0\/_0401_ ), .X(\u0\/_0133_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0898_ ( .A(\u0\/u2\/_0015_ ), .B(\w0\[15\] ), .X(\u0\/_0418_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0899_ ( .A(\u0\/rcon\[15\] ), .B(\u0\/_0418_ ), .X(\u0\/_0419_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0900_ ( .A0(\u0\/_0419_ ), .A1(\key[111] ), .S(\u0\/_0401_ ), .X(\u0\/_0134_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0901_ ( .A(\u0\/u1\/_0008_ ), .B(\w0\[16\] ), .X(\u0\/_0420_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0902_ ( .A(\u0\/rcon\[16\] ), .B(\u0\/_0420_ ), .X(\u0\/_0421_ ) );
sky130_fd_sc_hd__buf_2 \u0/_0903_ ( .A(\u0\/_0387_ ), .X(\u0\/_0422_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0904_ ( .A0(\u0\/_0421_ ), .A1(\key[112] ), .S(\u0\/_0422_ ), .X(\u0\/_0135_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0905_ ( .A(\u0\/u1\/_0009_ ), .B(\w0\[17\] ), .X(\u0\/_0423_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0906_ ( .A(\u0\/rcon\[17\] ), .B(\u0\/_0423_ ), .X(\u0\/_0424_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0907_ ( .A0(\u0\/_0424_ ), .A1(\key[113] ), .S(\u0\/_0422_ ), .X(\u0\/_0136_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0908_ ( .A(\u0\/u1\/_0010_ ), .B(\w0\[18\] ), .X(\u0\/_0425_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0909_ ( .A(\u0\/rcon\[18\] ), .B(\u0\/_0425_ ), .X(\u0\/_0426_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0910_ ( .A0(\u0\/_0426_ ), .A1(\key[114] ), .S(\u0\/_0422_ ), .X(\u0\/_0137_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0911_ ( .A(\u0\/u1\/_0011_ ), .B(\w0\[19\] ), .X(\u0\/_0427_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0912_ ( .A(\u0\/rcon\[19\] ), .B(\u0\/_0427_ ), .X(\u0\/_0428_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0913_ ( .A0(\u0\/_0428_ ), .A1(\key[115] ), .S(\u0\/_0422_ ), .X(\u0\/_0138_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0914_ ( .A(\u0\/u1\/_0012_ ), .B(\w0\[20\] ), .X(\u0\/_0429_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0915_ ( .A(\u0\/rcon\[20\] ), .B(\u0\/_0429_ ), .X(\u0\/_0430_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0916_ ( .A0(\u0\/_0430_ ), .A1(\key[116] ), .S(\u0\/_0422_ ), .X(\u0\/_0140_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0917_ ( .A(\u0\/u1\/_0013_ ), .B(\w0\[21\] ), .X(\u0\/_0431_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0918_ ( .A(\u0\/rcon\[21\] ), .B(\u0\/_0431_ ), .X(\u0\/_0432_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0919_ ( .A0(\u0\/_0432_ ), .A1(\key[117] ), .S(\u0\/_0422_ ), .X(\u0\/_0141_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0920_ ( .A(\u0\/u1\/_0014_ ), .B(\w0\[22\] ), .X(\u0\/_0433_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0921_ ( .A(\u0\/rcon\[22\] ), .B(\u0\/_0433_ ), .X(\u0\/_0434_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0922_ ( .A0(\u0\/_0434_ ), .A1(\key[118] ), .S(\u0\/_0422_ ), .X(\u0\/_0142_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0923_ ( .A(\u0\/u1\/_0015_ ), .B(\w0\[23\] ), .X(\u0\/_0435_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0924_ ( .A(\u0\/rcon\[23\] ), .B(\u0\/_0435_ ), .X(\u0\/_0436_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0925_ ( .A0(\u0\/_0436_ ), .A1(\key[119] ), .S(\u0\/_0422_ ), .X(\u0\/_0143_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0926_ ( .A(\u0\/u0\/_0008_ ), .B(\w0\[24\] ), .X(\u0\/_0437_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0927_ ( .A(\u0\/rcon\[24\] ), .B(\u0\/_0437_ ), .X(\u0\/_0438_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0928_ ( .A0(\u0\/_0438_ ), .A1(\key[120] ), .S(\u0\/_0422_ ), .X(\u0\/_0144_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0929_ ( .A(\u0\/u0\/_0009_ ), .B(\w0\[25\] ), .X(\u0\/_0439_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0930_ ( .A(\u0\/rcon\[25\] ), .B(\u0\/_0439_ ), .X(\u0\/_0440_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0931_ ( .A0(\u0\/_0440_ ), .A1(\key[121] ), .S(\u0\/_0422_ ), .X(\u0\/_0145_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0932_ ( .A(\u0\/u0\/_0010_ ), .B(\w0\[26\] ), .X(\u0\/_0441_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0933_ ( .A(\u0\/rcon\[26\] ), .B(\u0\/_0441_ ), .X(\u0\/_0442_ ) );
sky130_fd_sc_hd__buf_2 \u0/_0934_ ( .A(\u0\/_0387_ ), .X(\u0\/_0443_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0935_ ( .A0(\u0\/_0442_ ), .A1(\key[122] ), .S(\u0\/_0443_ ), .X(\u0\/_0146_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0936_ ( .A(\u0\/u0\/_0011_ ), .B(\w0\[27\] ), .X(\u0\/_0444_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0937_ ( .A(\u0\/rcon\[27\] ), .B(\u0\/_0444_ ), .X(\u0\/_0445_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0938_ ( .A0(\u0\/_0445_ ), .A1(\key[123] ), .S(\u0\/_0443_ ), .X(\u0\/_0147_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0939_ ( .A(\u0\/u0\/_0012_ ), .B(\w0\[28\] ), .X(\u0\/_0446_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0940_ ( .A(\u0\/rcon\[28\] ), .B(\u0\/_0446_ ), .X(\u0\/_0447_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0941_ ( .A0(\u0\/_0447_ ), .A1(\key[124] ), .S(\u0\/_0443_ ), .X(\u0\/_0148_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0942_ ( .A(\u0\/u0\/_0013_ ), .B(\w0\[29\] ), .X(\u0\/_0448_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0943_ ( .A(\u0\/rcon\[29\] ), .B(\u0\/_0448_ ), .X(\u0\/_0449_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0944_ ( .A0(\u0\/_0449_ ), .A1(\key[125] ), .S(\u0\/_0443_ ), .X(\u0\/_0149_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0945_ ( .A(\u0\/u0\/_0014_ ), .B(\w0\[30\] ), .X(\u0\/_0450_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0946_ ( .A(\u0\/rcon\[30\] ), .B(\u0\/_0450_ ), .X(\u0\/_0451_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0947_ ( .A0(\u0\/_0451_ ), .A1(\key[126] ), .S(\u0\/_0443_ ), .X(\u0\/_0151_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0948_ ( .A(\u0\/u0\/_0015_ ), .B(\w0\[31\] ), .X(\u0\/_0452_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_0949_ ( .A(\u0\/rcon\[31\] ), .B(\u0\/_0452_ ), .X(\u0\/_0453_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_0950_ ( .A0(\u0\/_0453_ ), .A1(\key[127] ), .S(\u0\/_0443_ ), .X(\u0\/_0152_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/_0951_ ( .A(\u0\/_0387_ ), .X(\u0\/_0454_ ) );
sky130_fd_sc_hd__buf_2 \u0/_0952_ ( .A(\u0\/_0454_ ), .X(\u0\/_0455_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_0953_ ( .A1(\w1\[0\] ), .A2(\u0\/_0386_ ), .B1_N(\u0\/_0387_ ), .Y(\u0\/_0456_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_0954_ ( .A1(\w1\[0\] ), .A2(\u0\/_0386_ ), .B1(\u0\/_0456_ ), .X(\u0\/_0457_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_0955_ ( .A1(\u0\/_0455_ ), .A2(\key[64] ), .B1_N(\u0\/_0457_ ), .X(\u0\/_0160_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_0956_ ( .A1(\w1\[1\] ), .A2(\u0\/_0390_ ), .B1_N(\u0\/_0387_ ), .Y(\u0\/_0458_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_0957_ ( .A1(\w1\[1\] ), .A2(\u0\/_0390_ ), .B1(\u0\/_0458_ ), .X(\u0\/_0459_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_0958_ ( .A1(\u0\/_0455_ ), .A2(\key[65] ), .B1_N(\u0\/_0459_ ), .X(\u0\/_0171_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/_0959_ ( .A(ld ), .X(\u0\/_0460_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_0960_ ( .A1(\w1\[2\] ), .A2(\u0\/_0392_ ), .B1_N(\u0\/_0460_ ), .Y(\u0\/_0461_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_0961_ ( .A1(\w1\[2\] ), .A2(\u0\/_0392_ ), .B1(\u0\/_0461_ ), .X(\u0\/_0462_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_0962_ ( .A1(\u0\/_0455_ ), .A2(\key[66] ), .B1_N(\u0\/_0462_ ), .X(\u0\/_0182_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_0963_ ( .A1(\w1\[3\] ), .A2(\u0\/_0394_ ), .B1_N(\u0\/_0460_ ), .Y(\u0\/_0463_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_0964_ ( .A1(\w1\[3\] ), .A2(\u0\/_0394_ ), .B1(\u0\/_0463_ ), .X(\u0\/_0464_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_0965_ ( .A1(\u0\/_0455_ ), .A2(\key[67] ), .B1_N(\u0\/_0464_ ), .X(\u0\/_0185_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_0966_ ( .A1(\w1\[4\] ), .A2(\u0\/_0396_ ), .B1_N(\u0\/_0460_ ), .Y(\u0\/_0465_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_0967_ ( .A1(\w1\[4\] ), .A2(\u0\/_0396_ ), .B1(\u0\/_0465_ ), .X(\u0\/_0466_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_0968_ ( .A1(\u0\/_0455_ ), .A2(\key[68] ), .B1_N(\u0\/_0466_ ), .X(\u0\/_0186_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_0969_ ( .A1(\w1\[5\] ), .A2(\u0\/_0398_ ), .B1_N(\u0\/_0460_ ), .Y(\u0\/_0467_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_0970_ ( .A1(\w1\[5\] ), .A2(\u0\/_0398_ ), .B1(\u0\/_0467_ ), .X(\u0\/_0468_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_0971_ ( .A1(\u0\/_0455_ ), .A2(\key[69] ), .B1_N(\u0\/_0468_ ), .X(\u0\/_0187_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_0972_ ( .A1(\w1\[6\] ), .A2(\u0\/_0400_ ), .B1_N(\u0\/_0460_ ), .Y(\u0\/_0469_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_0973_ ( .A1(\w1\[6\] ), .A2(\u0\/_0400_ ), .B1(\u0\/_0469_ ), .X(\u0\/_0470_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_0974_ ( .A1(\u0\/_0455_ ), .A2(\key[70] ), .B1_N(\u0\/_0470_ ), .X(\u0\/_0188_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_0975_ ( .A1(\w1\[7\] ), .A2(\u0\/_0403_ ), .B1_N(\u0\/_0460_ ), .Y(\u0\/_0471_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_0976_ ( .A1(\w1\[7\] ), .A2(\u0\/_0403_ ), .B1(\u0\/_0471_ ), .X(\u0\/_0472_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_0977_ ( .A1(\u0\/_0455_ ), .A2(\key[71] ), .B1_N(\u0\/_0472_ ), .X(\u0\/_0189_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_0978_ ( .A1(\w1\[8\] ), .A2(\u0\/_0405_ ), .B1_N(\u0\/_0460_ ), .Y(\u0\/_0473_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_0979_ ( .A1(\w1\[8\] ), .A2(\u0\/_0405_ ), .B1(\u0\/_0473_ ), .X(\u0\/_0474_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_0980_ ( .A1(\u0\/_0455_ ), .A2(\key[72] ), .B1_N(\u0\/_0474_ ), .X(\u0\/_0190_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_0981_ ( .A1(\w1\[9\] ), .A2(\u0\/_0407_ ), .B1_N(\u0\/_0460_ ), .Y(\u0\/_0475_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_0982_ ( .A1(\w1\[9\] ), .A2(\u0\/_0407_ ), .B1(\u0\/_0475_ ), .X(\u0\/_0476_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_0983_ ( .A1(\u0\/_0455_ ), .A2(\key[73] ), .B1_N(\u0\/_0476_ ), .X(\u0\/_0191_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_0985_ ( .A1(\w1\[10\] ), .A2(\u0\/_0409_ ), .B1_N(\u0\/_0460_ ), .Y(\u0\/_0478_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_0986_ ( .A1(\w1\[10\] ), .A2(\u0\/_0409_ ), .B1(\u0\/_0478_ ), .X(\u0\/_0479_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_0987_ ( .A1(\u0\/_0455_ ), .A2(\key[74] ), .B1_N(\u0\/_0479_ ), .X(\u0\/_0161_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_0988_ ( .A1(\w1\[11\] ), .A2(\u0\/_0411_ ), .B1_N(\u0\/_0460_ ), .Y(\u0\/_0480_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_0989_ ( .A1(\w1\[11\] ), .A2(\u0\/_0411_ ), .B1(\u0\/_0480_ ), .X(\u0\/_0481_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_0990_ ( .A1(\u0\/_0455_ ), .A2(\key[75] ), .B1_N(\u0\/_0481_ ), .X(\u0\/_0162_ ) );
sky130_fd_sc_hd__buf_2 \u0/_0991_ ( .A(ld ), .X(\u0\/_0482_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_0992_ ( .A1(\w1\[12\] ), .A2(\u0\/_0413_ ), .B1_N(\u0\/_0482_ ), .Y(\u0\/_0483_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_0993_ ( .A1(\w1\[12\] ), .A2(\u0\/_0413_ ), .B1(\u0\/_0483_ ), .X(\u0\/_0484_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_0994_ ( .A1(\u0\/_0455_ ), .A2(\key[76] ), .B1_N(\u0\/_0484_ ), .X(\u0\/_0163_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_0995_ ( .A1(\w1\[13\] ), .A2(\u0\/_0415_ ), .B1_N(\u0\/_0482_ ), .Y(\u0\/_0485_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_0996_ ( .A1(\w1\[13\] ), .A2(\u0\/_0415_ ), .B1(\u0\/_0485_ ), .X(\u0\/_0486_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_0997_ ( .A1(\u0\/_0455_ ), .A2(\key[77] ), .B1_N(\u0\/_0486_ ), .X(\u0\/_0164_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_0998_ ( .A1(\w1\[14\] ), .A2(\u0\/_0417_ ), .B1_N(\u0\/_0482_ ), .Y(\u0\/_0487_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_0999_ ( .A1(\w1\[14\] ), .A2(\u0\/_0417_ ), .B1(\u0\/_0487_ ), .X(\u0\/_0488_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1000_ ( .A1(\u0\/_0455_ ), .A2(\key[78] ), .B1_N(\u0\/_0488_ ), .X(\u0\/_0165_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1001_ ( .A1(\w1\[15\] ), .A2(\u0\/_0419_ ), .B1_N(\u0\/_0482_ ), .Y(\u0\/_0489_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1002_ ( .A1(\w1\[15\] ), .A2(\u0\/_0419_ ), .B1(\u0\/_0489_ ), .X(\u0\/_0490_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1003_ ( .A1(\u0\/_0455_ ), .A2(\key[79] ), .B1_N(\u0\/_0490_ ), .X(\u0\/_0166_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1004_ ( .A1(\w1\[16\] ), .A2(\u0\/_0421_ ), .B1_N(\u0\/_0482_ ), .Y(\u0\/_0491_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1005_ ( .A1(\w1\[16\] ), .A2(\u0\/_0421_ ), .B1(\u0\/_0491_ ), .X(\u0\/_0492_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1006_ ( .A1(\u0\/_0455_ ), .A2(\key[80] ), .B1_N(\u0\/_0492_ ), .X(\u0\/_0167_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1007_ ( .A1(\w1\[17\] ), .A2(\u0\/_0424_ ), .B1_N(\u0\/_0482_ ), .Y(\u0\/_0493_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1008_ ( .A1(\w1\[17\] ), .A2(\u0\/_0424_ ), .B1(\u0\/_0493_ ), .X(\u0\/_0494_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1009_ ( .A1(\u0\/_0455_ ), .A2(\key[81] ), .B1_N(\u0\/_0494_ ), .X(\u0\/_0168_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1010_ ( .A1(\w1\[18\] ), .A2(\u0\/_0426_ ), .B1_N(\u0\/_0482_ ), .Y(\u0\/_0495_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1011_ ( .A1(\w1\[18\] ), .A2(\u0\/_0426_ ), .B1(\u0\/_0495_ ), .X(\u0\/_0496_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1012_ ( .A1(\u0\/_0455_ ), .A2(\key[82] ), .B1_N(\u0\/_0496_ ), .X(\u0\/_0169_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1013_ ( .A1(\w1\[19\] ), .A2(\u0\/_0428_ ), .B1_N(\u0\/_0482_ ), .Y(\u0\/_0497_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1014_ ( .A1(\w1\[19\] ), .A2(\u0\/_0428_ ), .B1(\u0\/_0497_ ), .X(\u0\/_0498_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1015_ ( .A1(\u0\/_0455_ ), .A2(\key[83] ), .B1_N(\u0\/_0498_ ), .X(\u0\/_0170_ ) );
sky130_fd_sc_hd__buf_2 \u0/_1016_ ( .A(\u0\/_0387_ ), .X(\u0\/_0499_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1017_ ( .A1(\w1\[20\] ), .A2(\u0\/_0430_ ), .B1_N(\u0\/_0482_ ), .Y(\u0\/_0500_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1018_ ( .A1(\w1\[20\] ), .A2(\u0\/_0430_ ), .B1(\u0\/_0500_ ), .X(\u0\/_0501_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1019_ ( .A1(\u0\/_0499_ ), .A2(\key[84] ), .B1_N(\u0\/_0501_ ), .X(\u0\/_0172_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1020_ ( .A1(\w1\[21\] ), .A2(\u0\/_0432_ ), .B1_N(\u0\/_0482_ ), .Y(\u0\/_0502_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1021_ ( .A1(\w1\[21\] ), .A2(\u0\/_0432_ ), .B1(\u0\/_0502_ ), .X(\u0\/_0503_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1022_ ( .A1(\u0\/_0499_ ), .A2(\key[85] ), .B1_N(\u0\/_0503_ ), .X(\u0\/_0173_ ) );
sky130_fd_sc_hd__buf_2 \u0/_1023_ ( .A(ld ), .X(\u0\/_0504_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1024_ ( .A1(\w1\[22\] ), .A2(\u0\/_0434_ ), .B1_N(\u0\/_0504_ ), .Y(\u0\/_0505_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1025_ ( .A1(\w1\[22\] ), .A2(\u0\/_0434_ ), .B1(\u0\/_0505_ ), .X(\u0\/_0506_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1026_ ( .A1(\u0\/_0499_ ), .A2(\key[86] ), .B1_N(\u0\/_0506_ ), .X(\u0\/_0174_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1027_ ( .A1(\w1\[23\] ), .A2(\u0\/_0436_ ), .B1_N(\u0\/_0504_ ), .Y(\u0\/_0507_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1028_ ( .A1(\w1\[23\] ), .A2(\u0\/_0436_ ), .B1(\u0\/_0507_ ), .X(\u0\/_0508_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1029_ ( .A1(\u0\/_0499_ ), .A2(\key[87] ), .B1_N(\u0\/_0508_ ), .X(\u0\/_0175_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1030_ ( .A1(\w1\[24\] ), .A2(\u0\/_0438_ ), .B1_N(\u0\/_0504_ ), .Y(\u0\/_0509_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1031_ ( .A1(\w1\[24\] ), .A2(\u0\/_0438_ ), .B1(\u0\/_0509_ ), .X(\u0\/_0510_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1032_ ( .A1(\u0\/_0499_ ), .A2(\key[88] ), .B1_N(\u0\/_0510_ ), .X(\u0\/_0176_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1033_ ( .A1(\w1\[25\] ), .A2(\u0\/_0440_ ), .B1_N(\u0\/_0504_ ), .Y(\u0\/_0511_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1034_ ( .A1(\w1\[25\] ), .A2(\u0\/_0440_ ), .B1(\u0\/_0511_ ), .X(\u0\/_0512_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1035_ ( .A1(\u0\/_0499_ ), .A2(\key[89] ), .B1_N(\u0\/_0512_ ), .X(\u0\/_0177_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1036_ ( .A1(\w1\[26\] ), .A2(\u0\/_0442_ ), .B1_N(\u0\/_0504_ ), .Y(\u0\/_0513_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1037_ ( .A1(\w1\[26\] ), .A2(\u0\/_0442_ ), .B1(\u0\/_0513_ ), .X(\u0\/_0514_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1038_ ( .A1(\u0\/_0499_ ), .A2(\key[90] ), .B1_N(\u0\/_0514_ ), .X(\u0\/_0178_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1039_ ( .A1(\w1\[27\] ), .A2(\u0\/_0445_ ), .B1_N(\u0\/_0504_ ), .Y(\u0\/_0515_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1040_ ( .A1(\w1\[27\] ), .A2(\u0\/_0445_ ), .B1(\u0\/_0515_ ), .X(\u0\/_0516_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1041_ ( .A1(\u0\/_0499_ ), .A2(\key[91] ), .B1_N(\u0\/_0516_ ), .X(\u0\/_0179_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1042_ ( .A1(\w1\[28\] ), .A2(\u0\/_0447_ ), .B1_N(\u0\/_0504_ ), .Y(\u0\/_0517_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1043_ ( .A1(\w1\[28\] ), .A2(\u0\/_0447_ ), .B1(\u0\/_0517_ ), .X(\u0\/_0518_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1044_ ( .A1(\u0\/_0499_ ), .A2(\key[92] ), .B1_N(\u0\/_0518_ ), .X(\u0\/_0180_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1045_ ( .A1(\w1\[29\] ), .A2(\u0\/_0449_ ), .B1_N(\u0\/_0504_ ), .Y(\u0\/_0519_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1046_ ( .A1(\w1\[29\] ), .A2(\u0\/_0449_ ), .B1(\u0\/_0519_ ), .X(\u0\/_0520_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1047_ ( .A1(\u0\/_0499_ ), .A2(\key[93] ), .B1_N(\u0\/_0520_ ), .X(\u0\/_0181_ ) );
sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 \u0/_1048_ ( .A(ld ), .X(\u0\/_0521_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1049_ ( .A1(\w1\[30\] ), .A2(\u0\/_0451_ ), .B1_N(\u0\/_0504_ ), .Y(\u0\/_0522_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1050_ ( .A1(\w1\[30\] ), .A2(\u0\/_0451_ ), .B1(\u0\/_0522_ ), .X(\u0\/_0523_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1051_ ( .A1(\u0\/_0521_ ), .A2(\key[94] ), .B1_N(\u0\/_0523_ ), .X(\u0\/_0183_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/_1052_ ( .A1(\w1\[31\] ), .A2(\u0\/_0453_ ), .B1_N(\u0\/_0504_ ), .Y(\u0\/_0524_ ) );
sky130_fd_sc_hd__a21o_1 \u0/_1053_ ( .A1(\w1\[31\] ), .A2(\u0\/_0453_ ), .B1(\u0\/_0524_ ), .X(\u0\/_0525_ ) );
sky130_fd_sc_hd__a21bo_1 \u0/_1054_ ( .A1(\u0\/_0521_ ), .A2(\key[95] ), .B1_N(\u0\/_0525_ ), .X(\u0\/_0184_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1055_ ( .A0(\w2\[0\] ), .A1(\key[32] ), .S(\u0\/_0521_ ), .Y(\u0\/_0526_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1056_ ( .A0(\w2\[0\] ), .A1(\u0\/_0526_ ), .S(\u0\/_0457_ ), .Y(\u0\/_0192_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1057_ ( .A0(\w2\[1\] ), .A1(\key[33] ), .S(\u0\/_0521_ ), .Y(\u0\/_0527_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1058_ ( .A0(\w2\[1\] ), .A1(\u0\/_0527_ ), .S(\u0\/_0459_ ), .Y(\u0\/_0203_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1059_ ( .A0(\w2\[2\] ), .A1(\key[34] ), .S(\u0\/_0521_ ), .Y(\u0\/_0528_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1060_ ( .A0(\w2\[2\] ), .A1(\u0\/_0528_ ), .S(\u0\/_0462_ ), .Y(\u0\/_0214_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1061_ ( .A0(\w2\[3\] ), .A1(\key[35] ), .S(\u0\/_0521_ ), .Y(\u0\/_0529_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1062_ ( .A0(\w2\[3\] ), .A1(\u0\/_0529_ ), .S(\u0\/_0464_ ), .Y(\u0\/_0217_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1063_ ( .A0(\w2\[4\] ), .A1(\key[36] ), .S(\u0\/_0521_ ), .Y(\u0\/_0530_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1064_ ( .A0(\w2\[4\] ), .A1(\u0\/_0530_ ), .S(\u0\/_0466_ ), .Y(\u0\/_0218_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1065_ ( .A0(\w2\[5\] ), .A1(\key[37] ), .S(\u0\/_0521_ ), .Y(\u0\/_0531_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1066_ ( .A0(\w2\[5\] ), .A1(\u0\/_0531_ ), .S(\u0\/_0468_ ), .Y(\u0\/_0219_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1067_ ( .A0(\w2\[6\] ), .A1(\key[38] ), .S(\u0\/_0521_ ), .Y(\u0\/_0532_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1068_ ( .A0(\w2\[6\] ), .A1(\u0\/_0532_ ), .S(\u0\/_0470_ ), .Y(\u0\/_0220_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1069_ ( .A0(\w2\[7\] ), .A1(\key[39] ), .S(\u0\/_0521_ ), .Y(\u0\/_0533_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1070_ ( .A0(\w2\[7\] ), .A1(\u0\/_0533_ ), .S(\u0\/_0472_ ), .Y(\u0\/_0221_ ) );
sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 \u0/_1071_ ( .A(ld ), .X(\u0\/_0534_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1072_ ( .A0(\w2\[8\] ), .A1(\key[40] ), .S(\u0\/_0534_ ), .Y(\u0\/_0535_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1073_ ( .A0(\w2\[8\] ), .A1(\u0\/_0535_ ), .S(\u0\/_0474_ ), .Y(\u0\/_0222_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1074_ ( .A0(\w2\[9\] ), .A1(\key[41] ), .S(\u0\/_0534_ ), .Y(\u0\/_0536_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1075_ ( .A0(\w2\[9\] ), .A1(\u0\/_0536_ ), .S(\u0\/_0476_ ), .Y(\u0\/_0223_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1076_ ( .A0(\w2\[10\] ), .A1(\key[42] ), .S(\u0\/_0534_ ), .Y(\u0\/_0537_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1077_ ( .A0(\w2\[10\] ), .A1(\u0\/_0537_ ), .S(\u0\/_0479_ ), .Y(\u0\/_0193_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1078_ ( .A0(\w2\[11\] ), .A1(\key[43] ), .S(\u0\/_0534_ ), .Y(\u0\/_0538_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1079_ ( .A0(\w2\[11\] ), .A1(\u0\/_0538_ ), .S(\u0\/_0481_ ), .Y(\u0\/_0194_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1080_ ( .A0(\w2\[12\] ), .A1(\key[44] ), .S(\u0\/_0534_ ), .Y(\u0\/_0539_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1081_ ( .A0(\w2\[12\] ), .A1(\u0\/_0539_ ), .S(\u0\/_0484_ ), .Y(\u0\/_0195_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1082_ ( .A0(\w2\[13\] ), .A1(\key[45] ), .S(\u0\/_0534_ ), .Y(\u0\/_0540_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1083_ ( .A0(\w2\[13\] ), .A1(\u0\/_0540_ ), .S(\u0\/_0486_ ), .Y(\u0\/_0196_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1084_ ( .A0(\w2\[14\] ), .A1(\key[46] ), .S(\u0\/_0534_ ), .Y(\u0\/_0541_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1085_ ( .A0(\w2\[14\] ), .A1(\u0\/_0541_ ), .S(\u0\/_0488_ ), .Y(\u0\/_0197_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1086_ ( .A0(\w2\[15\] ), .A1(\key[47] ), .S(\u0\/_0534_ ), .Y(\u0\/_0542_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1087_ ( .A0(\w2\[15\] ), .A1(\u0\/_0542_ ), .S(\u0\/_0490_ ), .Y(\u0\/_0198_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1088_ ( .A0(\w2\[16\] ), .A1(\key[48] ), .S(\u0\/_0534_ ), .Y(\u0\/_0543_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1089_ ( .A0(\w2\[16\] ), .A1(\u0\/_0543_ ), .S(\u0\/_0492_ ), .Y(\u0\/_0199_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1090_ ( .A0(\w2\[17\] ), .A1(\key[49] ), .S(\u0\/_0534_ ), .Y(\u0\/_0544_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1091_ ( .A0(\w2\[17\] ), .A1(\u0\/_0544_ ), .S(\u0\/_0494_ ), .Y(\u0\/_0200_ ) );
sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 \u0/_1092_ ( .A(ld ), .X(\u0\/_0545_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1093_ ( .A0(\w2\[18\] ), .A1(\key[50] ), .S(\u0\/_0545_ ), .Y(\u0\/_0546_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1094_ ( .A0(\w2\[18\] ), .A1(\u0\/_0546_ ), .S(\u0\/_0496_ ), .Y(\u0\/_0201_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1095_ ( .A0(\w2\[19\] ), .A1(\key[51] ), .S(\u0\/_0545_ ), .Y(\u0\/_0547_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1096_ ( .A0(\w2\[19\] ), .A1(\u0\/_0547_ ), .S(\u0\/_0498_ ), .Y(\u0\/_0202_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1097_ ( .A0(\w2\[20\] ), .A1(\key[52] ), .S(\u0\/_0545_ ), .Y(\u0\/_0548_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1098_ ( .A0(\w2\[20\] ), .A1(\u0\/_0548_ ), .S(\u0\/_0501_ ), .Y(\u0\/_0204_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1099_ ( .A0(\w2\[21\] ), .A1(\key[53] ), .S(\u0\/_0545_ ), .Y(\u0\/_0549_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1100_ ( .A0(\w2\[21\] ), .A1(\u0\/_0549_ ), .S(\u0\/_0503_ ), .Y(\u0\/_0205_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1101_ ( .A0(\w2\[22\] ), .A1(\key[54] ), .S(\u0\/_0545_ ), .Y(\u0\/_0550_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1102_ ( .A0(\w2\[22\] ), .A1(\u0\/_0550_ ), .S(\u0\/_0506_ ), .Y(\u0\/_0206_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1103_ ( .A0(\w2\[23\] ), .A1(\key[55] ), .S(\u0\/_0545_ ), .Y(\u0\/_0551_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1104_ ( .A0(\w2\[23\] ), .A1(\u0\/_0551_ ), .S(\u0\/_0508_ ), .Y(\u0\/_0207_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1105_ ( .A0(\w2\[24\] ), .A1(\key[56] ), .S(\u0\/_0545_ ), .Y(\u0\/_0552_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1106_ ( .A0(\w2\[24\] ), .A1(\u0\/_0552_ ), .S(\u0\/_0510_ ), .Y(\u0\/_0208_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1107_ ( .A0(\w2\[25\] ), .A1(\key[57] ), .S(\u0\/_0545_ ), .Y(\u0\/_0553_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1108_ ( .A0(\w2\[25\] ), .A1(\u0\/_0553_ ), .S(\u0\/_0512_ ), .Y(\u0\/_0209_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1109_ ( .A0(\w2\[26\] ), .A1(\key[58] ), .S(\u0\/_0545_ ), .Y(\u0\/_0554_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1110_ ( .A0(\w2\[26\] ), .A1(\u0\/_0554_ ), .S(\u0\/_0514_ ), .Y(\u0\/_0210_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1111_ ( .A0(\w2\[27\] ), .A1(\key[59] ), .S(\u0\/_0545_ ), .Y(\u0\/_0555_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1112_ ( .A0(\w2\[27\] ), .A1(\u0\/_0555_ ), .S(\u0\/_0516_ ), .Y(\u0\/_0211_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1113_ ( .A0(\w2\[28\] ), .A1(\key[60] ), .S(\u0\/_0388_ ), .Y(\u0\/_0556_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1114_ ( .A0(\w2\[28\] ), .A1(\u0\/_0556_ ), .S(\u0\/_0518_ ), .Y(\u0\/_0212_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1115_ ( .A0(\w2\[29\] ), .A1(\key[61] ), .S(\u0\/_0388_ ), .Y(\u0\/_0557_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1116_ ( .A0(\w2\[29\] ), .A1(\u0\/_0557_ ), .S(\u0\/_0520_ ), .Y(\u0\/_0213_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1117_ ( .A0(\w2\[30\] ), .A1(\key[62] ), .S(\u0\/_0388_ ), .Y(\u0\/_0558_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1118_ ( .A0(\w2\[30\] ), .A1(\u0\/_0558_ ), .S(\u0\/_0523_ ), .Y(\u0\/_0215_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1119_ ( .A0(\w2\[31\] ), .A1(\key[63] ), .S(\u0\/_0388_ ), .Y(\u0\/_0559_ ) );
sky130_fd_sc_hd__mux2i_1 \u0/_1120_ ( .A0(\w2\[31\] ), .A1(\u0\/_0559_ ), .S(\u0\/_0525_ ), .Y(\u0\/_0216_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1121_ ( .A(\u0\/rcon\[0\] ), .B(\w1\[0\] ), .Y(\u0\/_0560_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1122_ ( .A(\w2\[0\] ), .B(\w3\[0\] ), .X(\u0\/_0561_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1123_ ( .A(\u0\/_0560_ ), .B(\u0\/_0385_ ), .C(\u0\/_0561_ ), .X(\u0\/_0562_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1124_ ( .A0(\u0\/_0562_ ), .A1(\key[0] ), .S(\u0\/_0443_ ), .X(\u0\/_0224_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1125_ ( .A(\u0\/rcon\[1\] ), .B(\w1\[1\] ), .Y(\u0\/_0563_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1126_ ( .A(\w2\[1\] ), .B(\w3\[1\] ), .X(\u0\/_0564_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1127_ ( .A(\u0\/_0563_ ), .B(\u0\/_0389_ ), .C(\u0\/_0564_ ), .X(\u0\/_0565_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1128_ ( .A0(\u0\/_0565_ ), .A1(\key[1] ), .S(\u0\/_0443_ ), .X(\u0\/_0235_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1129_ ( .A(\u0\/rcon\[2\] ), .B(\w1\[2\] ), .Y(\u0\/_0566_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1130_ ( .A(\w2\[2\] ), .B(\w3\[2\] ), .X(\u0\/_0567_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1131_ ( .A(\u0\/_0566_ ), .B(\u0\/_0391_ ), .C(\u0\/_0567_ ), .X(\u0\/_0568_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1132_ ( .A0(\u0\/_0568_ ), .A1(\key[2] ), .S(\u0\/_0443_ ), .X(\u0\/_0246_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1133_ ( .A(\u0\/rcon\[3\] ), .B(\w1\[3\] ), .Y(\u0\/_0569_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1134_ ( .A(\w2\[3\] ), .B(\w3\[3\] ), .X(\u0\/_0570_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1135_ ( .A(\u0\/_0569_ ), .B(\u0\/_0393_ ), .C(\u0\/_0570_ ), .X(\u0\/_0571_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1136_ ( .A0(\u0\/_0571_ ), .A1(\key[3] ), .S(\u0\/_0443_ ), .X(\u0\/_0249_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1137_ ( .A(\u0\/rcon\[4\] ), .B(\w1\[4\] ), .Y(\u0\/_0572_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1138_ ( .A(\w2\[4\] ), .B(\w3\[4\] ), .X(\u0\/_0573_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1139_ ( .A(\u0\/_0572_ ), .B(\u0\/_0395_ ), .C(\u0\/_0573_ ), .X(\u0\/_0574_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1141_ ( .A0(\u0\/_0574_ ), .A1(\key[4] ), .S(\u0\/_0443_ ), .X(\u0\/_0250_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1142_ ( .A(\u0\/rcon\[5\] ), .B(\w1\[5\] ), .Y(\u0\/_0576_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1143_ ( .A(\w2\[5\] ), .B(\w3\[5\] ), .X(\u0\/_0577_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1144_ ( .A(\u0\/_0576_ ), .B(\u0\/_0397_ ), .C(\u0\/_0577_ ), .X(\u0\/_0578_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1145_ ( .A0(\u0\/_0578_ ), .A1(\key[5] ), .S(\u0\/_0443_ ), .X(\u0\/_0251_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1146_ ( .A(\u0\/rcon\[6\] ), .B(\w1\[6\] ), .Y(\u0\/_0579_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1147_ ( .A(\w2\[6\] ), .B(\w3\[6\] ), .X(\u0\/_0580_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1148_ ( .A(\u0\/_0579_ ), .B(\u0\/_0399_ ), .C(\u0\/_0580_ ), .X(\u0\/_0581_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1149_ ( .A0(\u0\/_0581_ ), .A1(\key[6] ), .S(\u0\/_0443_ ), .X(\u0\/_0252_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1150_ ( .A(\u0\/rcon\[7\] ), .B(\w1\[7\] ), .Y(\u0\/_0582_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1151_ ( .A(\w2\[7\] ), .B(\w3\[7\] ), .X(\u0\/_0583_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1152_ ( .A(\u0\/_0582_ ), .B(\u0\/_0402_ ), .C(\u0\/_0583_ ), .X(\u0\/_0584_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1153_ ( .A0(\u0\/_0584_ ), .A1(\key[7] ), .S(\u0\/_0443_ ), .X(\u0\/_0253_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1154_ ( .A(\u0\/rcon\[8\] ), .B(\w1\[8\] ), .Y(\u0\/_0585_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1155_ ( .A(\w2\[8\] ), .B(\w3\[8\] ), .X(\u0\/_0586_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1156_ ( .A(\u0\/_0585_ ), .B(\u0\/_0404_ ), .C(\u0\/_0586_ ), .X(\u0\/_0587_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1157_ ( .A0(\u0\/_0587_ ), .A1(\key[8] ), .S(\u0\/_0443_ ), .X(\u0\/_0254_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1158_ ( .A(\u0\/rcon\[9\] ), .B(\w1\[9\] ), .Y(\u0\/_0588_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1159_ ( .A(\w2\[9\] ), .B(\w3\[9\] ), .X(\u0\/_0589_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1160_ ( .A(\u0\/_0588_ ), .B(\u0\/_0406_ ), .C(\u0\/_0589_ ), .X(\u0\/_0590_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1161_ ( .A0(\u0\/_0590_ ), .A1(\key[9] ), .S(\u0\/_0443_ ), .X(\u0\/_0255_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1162_ ( .A(\u0\/rcon\[10\] ), .B(\w1\[10\] ), .Y(\u0\/_0591_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1163_ ( .A(\w2\[10\] ), .B(\w3\[10\] ), .X(\u0\/_0592_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1164_ ( .A(\u0\/_0591_ ), .B(\u0\/_0408_ ), .C(\u0\/_0592_ ), .X(\u0\/_0593_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1165_ ( .A0(\u0\/_0593_ ), .A1(\key[10] ), .S(\u0\/_0443_ ), .X(\u0\/_0225_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1166_ ( .A(\u0\/rcon\[11\] ), .B(\w1\[11\] ), .Y(\u0\/_0594_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1167_ ( .A(\w2\[11\] ), .B(\w3\[11\] ), .X(\u0\/_0595_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1168_ ( .A(\u0\/_0594_ ), .B(\u0\/_0410_ ), .C(\u0\/_0595_ ), .X(\u0\/_0596_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1169_ ( .A0(\u0\/_0596_ ), .A1(\key[11] ), .S(\u0\/_0443_ ), .X(\u0\/_0226_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1170_ ( .A(\u0\/rcon\[12\] ), .B(\w1\[12\] ), .Y(\u0\/_0597_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1171_ ( .A(\w2\[12\] ), .B(\w3\[12\] ), .X(\u0\/_0598_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1172_ ( .A(\u0\/_0597_ ), .B(\u0\/_0412_ ), .C(\u0\/_0598_ ), .X(\u0\/_0599_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1173_ ( .A0(\u0\/_0599_ ), .A1(\key[12] ), .S(\u0\/_0443_ ), .X(\u0\/_0227_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1174_ ( .A(\u0\/rcon\[13\] ), .B(\w1\[13\] ), .Y(\u0\/_0600_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1175_ ( .A(\w2\[13\] ), .B(\w3\[13\] ), .X(\u0\/_0601_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1176_ ( .A(\u0\/_0600_ ), .B(\u0\/_0414_ ), .C(\u0\/_0601_ ), .X(\u0\/_0602_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1177_ ( .A0(\u0\/_0602_ ), .A1(\key[13] ), .S(\u0\/_0443_ ), .X(\u0\/_0228_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1178_ ( .A(\u0\/rcon\[14\] ), .B(\w1\[14\] ), .Y(\u0\/_0603_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1179_ ( .A(\w2\[14\] ), .B(\w3\[14\] ), .X(\u0\/_0604_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1180_ ( .A(\u0\/_0603_ ), .B(\u0\/_0416_ ), .C(\u0\/_0604_ ), .X(\u0\/_0605_ ) );
sky130_fd_sc_hd__buf_2 \u0/_1181_ ( .A(\u0\/_0387_ ), .X(\u0\/_0606_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1182_ ( .A0(\u0\/_0605_ ), .A1(\key[14] ), .S(\u0\/_0606_ ), .X(\u0\/_0229_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1183_ ( .A(\u0\/rcon\[15\] ), .B(\w1\[15\] ), .Y(\u0\/_0607_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1184_ ( .A(\w2\[15\] ), .B(\w3\[15\] ), .X(\u0\/_0608_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1185_ ( .A(\u0\/_0607_ ), .B(\u0\/_0418_ ), .C(\u0\/_0608_ ), .X(\u0\/_0609_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1186_ ( .A0(\u0\/_0609_ ), .A1(\key[15] ), .S(\u0\/_0606_ ), .X(\u0\/_0230_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1187_ ( .A(\u0\/rcon\[16\] ), .B(\w1\[16\] ), .Y(\u0\/_0610_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1188_ ( .A(\w2\[16\] ), .B(\w3\[16\] ), .X(\u0\/_0611_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1189_ ( .A(\u0\/_0610_ ), .B(\u0\/_0420_ ), .C(\u0\/_0611_ ), .X(\u0\/_0612_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1190_ ( .A0(\u0\/_0612_ ), .A1(\key[16] ), .S(\u0\/_0606_ ), .X(\u0\/_0231_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1191_ ( .A(\u0\/rcon\[17\] ), .B(\w1\[17\] ), .Y(\u0\/_0613_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1192_ ( .A(\w2\[17\] ), .B(\w3\[17\] ), .X(\u0\/_0614_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1193_ ( .A(\u0\/_0613_ ), .B(\u0\/_0423_ ), .C(\u0\/_0614_ ), .X(\u0\/_0615_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1194_ ( .A0(\u0\/_0615_ ), .A1(\key[17] ), .S(\u0\/_0606_ ), .X(\u0\/_0232_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1195_ ( .A(\u0\/rcon\[18\] ), .B(\w1\[18\] ), .Y(\u0\/_0616_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1196_ ( .A(\w2\[18\] ), .B(\w3\[18\] ), .X(\u0\/_0617_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1197_ ( .A(\u0\/_0616_ ), .B(\u0\/_0425_ ), .C(\u0\/_0617_ ), .X(\u0\/_0618_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1198_ ( .A0(\u0\/_0618_ ), .A1(\key[18] ), .S(\u0\/_0606_ ), .X(\u0\/_0233_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1199_ ( .A(\u0\/rcon\[19\] ), .B(\w1\[19\] ), .Y(\u0\/_0619_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1200_ ( .A(\w2\[19\] ), .B(\w3\[19\] ), .X(\u0\/_0620_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1201_ ( .A(\u0\/_0619_ ), .B(\u0\/_0427_ ), .C(\u0\/_0620_ ), .X(\u0\/_0621_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1202_ ( .A0(\u0\/_0621_ ), .A1(\key[19] ), .S(\u0\/_0606_ ), .X(\u0\/_0234_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1203_ ( .A(\u0\/rcon\[20\] ), .B(\w1\[20\] ), .Y(\u0\/_0622_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1204_ ( .A(\w2\[20\] ), .B(\w3\[20\] ), .X(\u0\/_0623_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1205_ ( .A(\u0\/_0622_ ), .B(\u0\/_0429_ ), .C(\u0\/_0623_ ), .X(\u0\/_0624_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1206_ ( .A0(\u0\/_0624_ ), .A1(\key[20] ), .S(\u0\/_0606_ ), .X(\u0\/_0236_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1207_ ( .A(\u0\/rcon\[21\] ), .B(\w1\[21\] ), .Y(\u0\/_0625_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1208_ ( .A(\w2\[21\] ), .B(\w3\[21\] ), .X(\u0\/_0626_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1209_ ( .A(\u0\/_0625_ ), .B(\u0\/_0431_ ), .C(\u0\/_0626_ ), .X(\u0\/_0627_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1210_ ( .A0(\u0\/_0627_ ), .A1(\key[21] ), .S(\u0\/_0606_ ), .X(\u0\/_0237_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1211_ ( .A(\u0\/rcon\[22\] ), .B(\w1\[22\] ), .Y(\u0\/_0628_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1212_ ( .A(\w2\[22\] ), .B(\w3\[22\] ), .X(\u0\/_0629_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1213_ ( .A(\u0\/_0628_ ), .B(\u0\/_0433_ ), .C(\u0\/_0629_ ), .X(\u0\/_0630_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1214_ ( .A0(\u0\/_0630_ ), .A1(\key[22] ), .S(\u0\/_0606_ ), .X(\u0\/_0238_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1215_ ( .A(\u0\/rcon\[23\] ), .B(\w1\[23\] ), .Y(\u0\/_0631_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1216_ ( .A(\w2\[23\] ), .B(\w3\[23\] ), .X(\u0\/_0632_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1217_ ( .A(\u0\/_0631_ ), .B(\u0\/_0435_ ), .C(\u0\/_0632_ ), .X(\u0\/_0633_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1218_ ( .A0(\u0\/_0633_ ), .A1(\key[23] ), .S(\u0\/_0606_ ), .X(\u0\/_0239_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1219_ ( .A(\u0\/rcon\[24\] ), .B(\w1\[24\] ), .Y(\u0\/_0634_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1220_ ( .A(\w2\[24\] ), .B(\w3\[24\] ), .X(\u0\/_0635_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1221_ ( .A(\u0\/_0634_ ), .B(\u0\/_0437_ ), .C(\u0\/_0635_ ), .X(\u0\/_0636_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1222_ ( .A0(\u0\/_0636_ ), .A1(\key[24] ), .S(\u0\/_0454_ ), .X(\u0\/_0240_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1223_ ( .A(\u0\/rcon\[25\] ), .B(\w1\[25\] ), .Y(\u0\/_0637_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1224_ ( .A(\w2\[25\] ), .B(\w3\[25\] ), .X(\u0\/_0638_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1225_ ( .A(\u0\/_0637_ ), .B(\u0\/_0439_ ), .C(\u0\/_0638_ ), .X(\u0\/_0639_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1226_ ( .A0(\u0\/_0639_ ), .A1(\key[25] ), .S(\u0\/_0454_ ), .X(\u0\/_0241_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1227_ ( .A(\u0\/rcon\[26\] ), .B(\w1\[26\] ), .Y(\u0\/_0640_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1228_ ( .A(\w2\[26\] ), .B(\w3\[26\] ), .X(\u0\/_0641_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1229_ ( .A(\u0\/_0640_ ), .B(\u0\/_0441_ ), .C(\u0\/_0641_ ), .X(\u0\/_0642_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1230_ ( .A0(\u0\/_0642_ ), .A1(\key[26] ), .S(\u0\/_0454_ ), .X(\u0\/_0242_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1231_ ( .A(\u0\/rcon\[27\] ), .B(\w1\[27\] ), .Y(\u0\/_0643_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1232_ ( .A(\w2\[27\] ), .B(\w3\[27\] ), .X(\u0\/_0644_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1233_ ( .A(\u0\/_0643_ ), .B(\u0\/_0444_ ), .C(\u0\/_0644_ ), .X(\u0\/_0645_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1234_ ( .A0(\u0\/_0645_ ), .A1(\key[27] ), .S(\u0\/_0454_ ), .X(\u0\/_0243_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1235_ ( .A(\u0\/rcon\[28\] ), .B(\w1\[28\] ), .Y(\u0\/_0646_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1236_ ( .A(\w2\[28\] ), .B(\w3\[28\] ), .X(\u0\/_0647_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1237_ ( .A(\u0\/_0646_ ), .B(\u0\/_0446_ ), .C(\u0\/_0647_ ), .X(\u0\/_0648_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1238_ ( .A0(\u0\/_0648_ ), .A1(\key[28] ), .S(\u0\/_0454_ ), .X(\u0\/_0244_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1239_ ( .A(\u0\/rcon\[29\] ), .B(\w1\[29\] ), .Y(\u0\/_0649_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1240_ ( .A(\w2\[29\] ), .B(\w3\[29\] ), .X(\u0\/_0650_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1241_ ( .A(\u0\/_0649_ ), .B(\u0\/_0448_ ), .C(\u0\/_0650_ ), .X(\u0\/_0651_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1242_ ( .A0(\u0\/_0651_ ), .A1(\key[29] ), .S(\u0\/_0454_ ), .X(\u0\/_0245_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1243_ ( .A(\u0\/rcon\[30\] ), .B(\w1\[30\] ), .Y(\u0\/_0652_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1244_ ( .A(\w2\[30\] ), .B(\w3\[30\] ), .X(\u0\/_0653_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1245_ ( .A(\u0\/_0652_ ), .B(\u0\/_0450_ ), .C(\u0\/_0653_ ), .X(\u0\/_0654_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1246_ ( .A0(\u0\/_0654_ ), .A1(\key[30] ), .S(\u0\/_0454_ ), .X(\u0\/_0247_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/_1247_ ( .A(\u0\/rcon\[31\] ), .B(\w1\[31\] ), .Y(\u0\/_0655_ ) );
sky130_fd_sc_hd__xor2_1 \u0/_1248_ ( .A(\w2\[31\] ), .B(\u0\/_0842_ ), .X(\u0\/_0656_ ) );
sky130_fd_sc_hd__xnor3_1 \u0/_1249_ ( .A(\u0\/_0655_ ), .B(\u0\/_0452_ ), .C(\u0\/_0656_ ), .X(\u0\/_0657_ ) );
sky130_fd_sc_hd__mux2_1 \u0/_1250_ ( .A0(\u0\/_0657_ ), .A1(\key[31] ), .S(\u0\/_0454_ ), .X(\u0\/_0248_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/_1697_ ( .A(\w3\[31\] ), .X(\u0\/_0842_ ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1700_ ( .D(\u0\/_0128_ ), .Q(\w0\[0\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1701_ ( .D(\u0\/_0139_ ), .Q(\w0\[1\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1702_ ( .D(\u0\/_0150_ ), .Q(\w0\[2\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1703_ ( .D(\u0\/_0153_ ), .Q(\w0\[3\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1704_ ( .D(\u0\/_0154_ ), .Q(\w0\[4\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1705_ ( .D(\u0\/_0155_ ), .Q(\w0\[5\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1706_ ( .D(\u0\/_0156_ ), .Q(\w0\[6\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1707_ ( .D(\u0\/_0157_ ), .Q(\w0\[7\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1708_ ( .D(\u0\/_0158_ ), .Q(\w0\[8\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1709_ ( .D(\u0\/_0159_ ), .Q(\w0\[9\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1710_ ( .D(\u0\/_0129_ ), .Q(\w0\[10\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1711_ ( .D(\u0\/_0130_ ), .Q(\w0\[11\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1712_ ( .D(\u0\/_0131_ ), .Q(\w0\[12\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1713_ ( .D(\u0\/_0132_ ), .Q(\w0\[13\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1714_ ( .D(\u0\/_0133_ ), .Q(\w0\[14\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1715_ ( .D(\u0\/_0134_ ), .Q(\w0\[15\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1716_ ( .D(\u0\/_0135_ ), .Q(\w0\[16\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1717_ ( .D(\u0\/_0136_ ), .Q(\w0\[17\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1718_ ( .D(\u0\/_0137_ ), .Q(\w0\[18\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1719_ ( .D(\u0\/_0138_ ), .Q(\w0\[19\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1720_ ( .D(\u0\/_0140_ ), .Q(\w0\[20\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1721_ ( .D(\u0\/_0141_ ), .Q(\w0\[21\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1722_ ( .D(\u0\/_0142_ ), .Q(\w0\[22\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1723_ ( .D(\u0\/_0143_ ), .Q(\w0\[23\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1724_ ( .D(\u0\/_0144_ ), .Q(\w0\[24\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1725_ ( .D(\u0\/_0145_ ), .Q(\w0\[25\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1726_ ( .D(\u0\/_0146_ ), .Q(\w0\[26\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1727_ ( .D(\u0\/_0147_ ), .Q(\w0\[27\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1728_ ( .D(\u0\/_0148_ ), .Q(\w0\[28\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1729_ ( .D(\u0\/_0149_ ), .Q(\w0\[29\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1730_ ( .D(\u0\/_0151_ ), .Q(\w0\[30\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1731_ ( .D(\u0\/_0152_ ), .Q(\w0\[31\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1732_ ( .D(\u0\/_0160_ ), .Q(\w1\[0\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1733_ ( .D(\u0\/_0171_ ), .Q(\w1\[1\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1734_ ( .D(\u0\/_0182_ ), .Q(\w1\[2\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1735_ ( .D(\u0\/_0185_ ), .Q(\w1\[3\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1736_ ( .D(\u0\/_0186_ ), .Q(\w1\[4\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1737_ ( .D(\u0\/_0187_ ), .Q(\w1\[5\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1738_ ( .D(\u0\/_0188_ ), .Q(\w1\[6\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1739_ ( .D(\u0\/_0189_ ), .Q(\w1\[7\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1740_ ( .D(\u0\/_0190_ ), .Q(\w1\[8\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1741_ ( .D(\u0\/_0191_ ), .Q(\w1\[9\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1742_ ( .D(\u0\/_0161_ ), .Q(\w1\[10\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1743_ ( .D(\u0\/_0162_ ), .Q(\w1\[11\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1744_ ( .D(\u0\/_0163_ ), .Q(\w1\[12\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1745_ ( .D(\u0\/_0164_ ), .Q(\w1\[13\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1746_ ( .D(\u0\/_0165_ ), .Q(\w1\[14\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1747_ ( .D(\u0\/_0166_ ), .Q(\w1\[15\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1748_ ( .D(\u0\/_0167_ ), .Q(\w1\[16\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1749_ ( .D(\u0\/_0168_ ), .Q(\w1\[17\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1750_ ( .D(\u0\/_0169_ ), .Q(\w1\[18\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1751_ ( .D(\u0\/_0170_ ), .Q(\w1\[19\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1752_ ( .D(\u0\/_0172_ ), .Q(\w1\[20\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1753_ ( .D(\u0\/_0173_ ), .Q(\w1\[21\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1754_ ( .D(\u0\/_0174_ ), .Q(\w1\[22\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1755_ ( .D(\u0\/_0175_ ), .Q(\w1\[23\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1756_ ( .D(\u0\/_0176_ ), .Q(\w1\[24\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1757_ ( .D(\u0\/_0177_ ), .Q(\w1\[25\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1758_ ( .D(\u0\/_0178_ ), .Q(\w1\[26\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1759_ ( .D(\u0\/_0179_ ), .Q(\w1\[27\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1760_ ( .D(\u0\/_0180_ ), .Q(\w1\[28\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1761_ ( .D(\u0\/_0181_ ), .Q(\w1\[29\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1762_ ( .D(\u0\/_0183_ ), .Q(\w1\[30\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1763_ ( .D(\u0\/_0184_ ), .Q(\w1\[31\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1764_ ( .D(\u0\/_0192_ ), .Q(\w2\[0\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1765_ ( .D(\u0\/_0203_ ), .Q(\w2\[1\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1766_ ( .D(\u0\/_0214_ ), .Q(\w2\[2\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1767_ ( .D(\u0\/_0217_ ), .Q(\w2\[3\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1768_ ( .D(\u0\/_0218_ ), .Q(\w2\[4\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1769_ ( .D(\u0\/_0219_ ), .Q(\w2\[5\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1770_ ( .D(\u0\/_0220_ ), .Q(\w2\[6\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1771_ ( .D(\u0\/_0221_ ), .Q(\w2\[7\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1772_ ( .D(\u0\/_0222_ ), .Q(\w2\[8\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1773_ ( .D(\u0\/_0223_ ), .Q(\w2\[9\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1774_ ( .D(\u0\/_0193_ ), .Q(\w2\[10\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1775_ ( .D(\u0\/_0194_ ), .Q(\w2\[11\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1776_ ( .D(\u0\/_0195_ ), .Q(\w2\[12\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1777_ ( .D(\u0\/_0196_ ), .Q(\w2\[13\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1778_ ( .D(\u0\/_0197_ ), .Q(\w2\[14\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1779_ ( .D(\u0\/_0198_ ), .Q(\w2\[15\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1780_ ( .D(\u0\/_0199_ ), .Q(\w2\[16\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1781_ ( .D(\u0\/_0200_ ), .Q(\w2\[17\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1782_ ( .D(\u0\/_0201_ ), .Q(\w2\[18\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1783_ ( .D(\u0\/_0202_ ), .Q(\w2\[19\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1784_ ( .D(\u0\/_0204_ ), .Q(\w2\[20\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1785_ ( .D(\u0\/_0205_ ), .Q(\w2\[21\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1786_ ( .D(\u0\/_0206_ ), .Q(\w2\[22\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1787_ ( .D(\u0\/_0207_ ), .Q(\w2\[23\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1788_ ( .D(\u0\/_0208_ ), .Q(\w2\[24\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1789_ ( .D(\u0\/_0209_ ), .Q(\w2\[25\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1790_ ( .D(\u0\/_0210_ ), .Q(\w2\[26\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1791_ ( .D(\u0\/_0211_ ), .Q(\w2\[27\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1792_ ( .D(\u0\/_0212_ ), .Q(\w2\[28\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1793_ ( .D(\u0\/_0213_ ), .Q(\w2\[29\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1794_ ( .D(\u0\/_0215_ ), .Q(\w2\[30\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1795_ ( .D(\u0\/_0216_ ), .Q(\w2\[31\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_2 \u0/_1796_ ( .D(\u0\/_0224_ ), .Q(\w3\[0\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_2 \u0/_1797_ ( .D(\u0\/_0235_ ), .Q(\w3\[1\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_2 \u0/_1798_ ( .D(\u0\/_0246_ ), .Q(\w3\[2\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_2 \u0/_1799_ ( .D(\u0\/_0249_ ), .Q(\w3\[3\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1800_ ( .D(\u0\/_0250_ ), .Q(\w3\[4\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1801_ ( .D(\u0\/_0251_ ), .Q(\w3\[5\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1802_ ( .D(\u0\/_0252_ ), .Q(\w3\[6\] ), .CLK(CTS_14 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1803_ ( .D(\u0\/_0253_ ), .Q(\w3\[7\] ), .CLK(CTS_20 ) );
sky130_fd_sc_hd__dfxtp_2 \u0/_1804_ ( .D(\u0\/_0254_ ), .Q(\w3\[8\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_2 \u0/_1805_ ( .D(\u0\/_0255_ ), .Q(\w3\[9\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1806_ ( .D(\u0\/_0225_ ), .Q(\w3\[10\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1807_ ( .D(\u0\/_0226_ ), .Q(\w3\[11\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1808_ ( .D(\u0\/_0227_ ), .Q(\w3\[12\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1809_ ( .D(\u0\/_0228_ ), .Q(\w3\[13\] ), .CLK(CTS_21 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1810_ ( .D(\u0\/_0229_ ), .Q(\w3\[14\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1811_ ( .D(\u0\/_0230_ ), .Q(\w3\[15\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_2 \u0/_1812_ ( .D(\u0\/_0231_ ), .Q(\w3\[16\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1813_ ( .D(\u0\/_0232_ ), .Q(\w3\[17\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_2 \u0/_1814_ ( .D(\u0\/_0233_ ), .Q(\w3\[18\] ), .CLK(CTS_7 ) );
sky130_fd_sc_hd__dfxtp_2 \u0/_1815_ ( .D(\u0\/_0234_ ), .Q(\w3\[19\] ), .CLK(CTS_1 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1816_ ( .D(\u0\/_0236_ ), .Q(\w3\[20\] ), .CLK(CTS_4 ) );
sky130_fd_sc_hd__dfxtp_2 \u0/_1817_ ( .D(\u0\/_0237_ ), .Q(\w3\[21\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_2 \u0/_1818_ ( .D(\u0\/_0238_ ), .Q(\w3\[22\] ), .CLK(CTS_9 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1819_ ( .D(\u0\/_0239_ ), .Q(\w3\[23\] ), .CLK(CTS_3 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1820_ ( .D(\u0\/_0240_ ), .Q(\w3\[24\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_2 \u0/_1821_ ( .D(\u0\/_0241_ ), .Q(\w3\[25\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1822_ ( .D(\u0\/_0242_ ), .Q(\w3\[26\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_2 \u0/_1823_ ( .D(\u0\/_0243_ ), .Q(\w3\[27\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1824_ ( .D(\u0\/_0244_ ), .Q(\w3\[28\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1825_ ( .D(\u0\/_0245_ ), .Q(\w3\[29\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1826_ ( .D(\u0\/_0247_ ), .Q(\w3\[30\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/_1827_ ( .D(\u0\/_0248_ ), .Q(\w3\[31\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_072_ ( .A(ld ), .X(\u0\/r0\/_049_ ) );
sky130_fd_sc_hd__a31o_1 \u0/r0/_073_ ( .A1(\u0\/r0\/rcnt\[0\] ), .A2(\u0\/r0\/rcnt\[1\] ), .A3(\u0\/r0\/rcnt\[2\] ), .B1(\u0\/r0\/_049_ ), .X(\u0\/r0\/_036_ ) );
sky130_fd_sc_hd__nand3b_1 \u0/r0/_074_ ( .A_N(\u0\/r0\/rcnt\[3\] ), .B(\u0\/r0\/rcnt\[0\] ), .C(\u0\/r0\/rcnt\[1\] ), .Y(\u0\/r0\/_050_ ) );
sky130_fd_sc_hd__or2b_1 \u0/r0/_075_ ( .A(\u0\/r0\/_050_ ), .B_N(\u0\/r0\/rcnt\[2\] ), .X(\u0\/r0\/_051_ ) );
sky130_fd_sc_hd__nor2_1 \u0/r0/_076_ ( .A(\u0\/r0\/rcnt\[0\] ), .B(ld ), .Y(\u0\/r0\/_044_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/r0/_077_ ( .A(\u0\/r0\/rcnt\[1\] ), .B(\u0\/r0\/rcnt\[2\] ), .C_N(\u0\/r0\/_044_ ), .Y(\u0\/r0\/_052_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/r0/_078_ ( .A1(\u0\/r0\/_049_ ), .A2(\u0\/r0\/_051_ ), .B1_N(\u0\/r0\/_052_ ), .Y(\u0\/r0\/_037_ ) );
sky130_fd_sc_hd__or2b_1 \u0/r0/_079_ ( .A(\u0\/r0\/rcnt\[1\] ), .B_N(\u0\/r0\/rcnt\[0\] ), .X(\u0\/r0\/_053_ ) );
sky130_fd_sc_hd__and2_1 \u0/r0/_080_ ( .A(\u0\/r0\/rcnt\[0\] ), .B(\u0\/r0\/rcnt\[1\] ), .X(\u0\/r0\/_054_ ) );
sky130_fd_sc_hd__xor2_1 \u0/r0/_081_ ( .A(\u0\/r0\/rcnt\[2\] ), .B(\u0\/r0\/_054_ ), .X(\u0\/r0\/_055_ ) );
sky130_fd_sc_hd__inv_1 \u0/r0/_082_ ( .A(\u0\/r0\/rcnt\[3\] ), .Y(\u0\/r0\/_056_ ) );
sky130_fd_sc_hd__and2_0 \u0/r0/_083_ ( .A(\u0\/r0\/_054_ ), .B(\u0\/r0\/rcnt\[2\] ), .X(\u0\/r0\/_057_ ) );
sky130_fd_sc_hd__xor2_1 \u0/r0/_084_ ( .A(\u0\/r0\/_056_ ), .B(\u0\/r0\/_057_ ), .X(\u0\/r0\/_058_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/r0/_085_ ( .A_N(\u0\/r0\/_055_ ), .B(\u0\/r0\/_058_ ), .Y(\u0\/r0\/_059_ ) );
sky130_fd_sc_hd__and2b_1 \u0/r0/_086_ ( .A_N(\u0\/r0\/rcnt\[2\] ), .B(\u0\/r0\/rcnt\[3\] ), .X(\u0\/r0\/_060_ ) );
sky130_fd_sc_hd__nand3b_1 \u0/r0/_087_ ( .A_N(\u0\/r0\/rcnt\[1\] ), .B(\u0\/r0\/_060_ ), .C(\u0\/r0\/_044_ ), .Y(\u0\/r0\/_061_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/r0/_088_ ( .A1(\u0\/r0\/_049_ ), .A2(\u0\/r0\/_053_ ), .A3(\u0\/r0\/_059_ ), .B1(\u0\/r0\/_061_ ), .Y(\u0\/r0\/_038_ ) );
sky130_fd_sc_hd__nand2_1 \u0/r0/_089_ ( .A(\u0\/r0\/_044_ ), .B(\u0\/r0\/rcnt\[1\] ), .Y(\u0\/r0\/_062_ ) );
sky130_fd_sc_hd__o22ai_1 \u0/r0/_090_ ( .A1(\u0\/r0\/_049_ ), .A2(\u0\/r0\/_051_ ), .B1(\u0\/r0\/_062_ ), .B2(\u0\/r0\/_059_ ), .Y(\u0\/r0\/_039_ ) );
sky130_fd_sc_hd__nor2_1 \u0/r0/_091_ ( .A(\u0\/r0\/rcnt\[0\] ), .B(\u0\/r0\/rcnt\[1\] ), .Y(\u0\/r0\/_063_ ) );
sky130_fd_sc_hd__nand2_1 \u0/r0/_092_ ( .A(\u0\/r0\/_060_ ), .B(\u0\/r0\/_063_ ), .Y(\u0\/r0\/_064_ ) );
sky130_fd_sc_hd__a21oi_1 \u0/r0/_093_ ( .A1(\u0\/r0\/_064_ ), .A2(\u0\/r0\/_050_ ), .B1(\u0\/r0\/_049_ ), .Y(\u0\/r0\/_040_ ) );
sky130_fd_sc_hd__nand2_1 \u0/r0/_094_ ( .A(\u0\/r0\/_055_ ), .B(\u0\/r0\/_056_ ), .Y(\u0\/r0\/_065_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/r0/_095_ ( .A(\u0\/r0\/_049_ ), .B(\u0\/r0\/_065_ ), .C_N(\u0\/r0\/_063_ ), .Y(\u0\/r0\/_066_ ) );
sky130_fd_sc_hd__o21bai_1 \u0/r0/_096_ ( .A1(\u0\/r0\/_049_ ), .A2(\u0\/r0\/_064_ ), .B1_N(\u0\/r0\/_066_ ), .Y(\u0\/r0\/_041_ ) );
sky130_fd_sc_hd__nor3_1 \u0/r0/_097_ ( .A(\u0\/r0\/_049_ ), .B(\u0\/r0\/_053_ ), .C(\u0\/r0\/_065_ ), .Y(\u0\/r0\/_042_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/r0/_098_ ( .A(\u0\/r0\/rcnt\[3\] ), .B(\u0\/r0\/_062_ ), .C_N(\u0\/r0\/_055_ ), .Y(\u0\/r0\/_043_ ) );
sky130_fd_sc_hd__nor3_1 \u0/r0/_099_ ( .A(\u0\/r0\/_049_ ), .B(\u0\/r0\/_063_ ), .C(\u0\/r0\/_054_ ), .Y(\u0\/r0\/_045_ ) );
sky130_fd_sc_hd__o21ba_1 \u0/r0/_100_ ( .A1(\u0\/r0\/rcnt\[2\] ), .A2(\u0\/r0\/_054_ ), .B1_N(\u0\/r0\/_036_ ), .X(\u0\/r0\/_046_ ) );
sky130_fd_sc_hd__nor2_1 \u0/r0/_101_ ( .A(\u0\/r0\/_049_ ), .B(\u0\/r0\/_058_ ), .Y(\u0\/r0\/_047_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_127_ ( .A(net25 ), .X(\u0\/rcon\[0\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_128_ ( .A(net26 ), .X(\u0\/rcon\[1\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_129_ ( .A(net27 ), .X(\u0\/rcon\[2\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_130_ ( .A(net28 ), .X(\u0\/rcon\[3\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_131_ ( .A(net29 ), .X(\u0\/rcon\[4\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_132_ ( .A(net30 ), .X(\u0\/rcon\[5\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_133_ ( .A(net31 ), .X(\u0\/rcon\[6\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_134_ ( .A(net32 ), .X(\u0\/rcon\[7\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_135_ ( .A(net33 ), .X(\u0\/rcon\[8\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_136_ ( .A(net34 ), .X(\u0\/rcon\[9\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_137_ ( .A(net35 ), .X(\u0\/rcon\[10\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_138_ ( .A(net36 ), .X(\u0\/rcon\[11\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_139_ ( .A(net37 ), .X(\u0\/rcon\[12\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_140_ ( .A(net38 ), .X(\u0\/rcon\[13\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_141_ ( .A(net39 ), .X(\u0\/rcon\[14\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_142_ ( .A(net40 ), .X(\u0\/rcon\[15\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_143_ ( .A(net41 ), .X(\u0\/rcon\[16\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_144_ ( .A(net42 ), .X(\u0\/rcon\[17\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_145_ ( .A(net43 ), .X(\u0\/rcon\[18\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_146_ ( .A(net44 ), .X(\u0\/rcon\[19\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_147_ ( .A(net45 ), .X(\u0\/rcon\[20\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_148_ ( .A(net46 ), .X(\u0\/rcon\[21\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_149_ ( .A(net47 ), .X(\u0\/rcon\[22\] ) );
sky130_fd_sc_hd__clkbuf_1 \u0/r0/_150_ ( .A(net48 ), .X(\u0\/rcon\[23\] ) );
sky130_fd_sc_hd__dfxtp_1 \u0/r0/_168_ ( .D(\u0\/r0\/_036_ ), .Q(\u0\/rcon\[24\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/r0/_169_ ( .D(\u0\/r0\/_037_ ), .Q(\u0\/rcon\[25\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/r0/_170_ ( .D(\u0\/r0\/_038_ ), .Q(\u0\/rcon\[26\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/r0/_171_ ( .D(\u0\/r0\/_039_ ), .Q(\u0\/rcon\[27\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/r0/_172_ ( .D(\u0\/r0\/_040_ ), .Q(\u0\/rcon\[28\] ), .CLK(CTS_17 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/r0/_173_ ( .D(\u0\/r0\/_041_ ), .Q(\u0\/rcon\[29\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/r0/_174_ ( .D(\u0\/r0\/_042_ ), .Q(\u0\/rcon\[30\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/r0/_175_ ( .D(\u0\/r0\/_043_ ), .Q(\u0\/rcon\[31\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/r0/_176_ ( .D(\u0\/r0\/_044_ ), .Q(\u0\/r0\/rcnt\[0\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/r0/_177_ ( .D(\u0\/r0\/_045_ ), .Q(\u0\/r0\/rcnt\[1\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/r0/_178_ ( .D(\u0\/r0\/_046_ ), .Q(\u0\/r0\/rcnt\[2\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__dfxtp_1 \u0/r0/_179_ ( .D(\u0\/r0\/_047_ ), .Q(\u0\/r0\/rcnt\[3\] ), .CLK(CTS_16 ) );
sky130_fd_sc_hd__nor2b_1 \u0/u0/_0753_ ( .A(\w3\[18\] ), .B_N(\w3\[19\] ), .Y(\u0\/u0\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \u0/u0/_0755_ ( .A(\u0\/u0\/_0001_ ), .B(\w3\[16\] ), .X(\u0\/u0\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \u0/u0/_0756_ ( .A(\u0\/u0\/_0096_ ), .B(\u0\/u0\/_0118_ ), .X(\u0\/u0\/_0129_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0757_ ( .A(\w3\[23\] ), .B(\w3\[22\] ), .X(\u0\/u0\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_0758_ ( .A(\w3\[20\] ), .B(\w3\[21\] ), .Y(\u0\/u0\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0759_ ( .A(\u0\/u0\/_0140_ ), .B(\u0\/u0\/_0151_ ), .X(\u0\/u0\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0761_ ( .A(\u0\/u0\/_0129_ ), .B(\u0\/u0\/_0162_ ), .X(\u0\/u0\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0762_ ( .A(\u0\/u0\/_0096_ ), .X(\u0\/u0\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u0/_0763_ ( .A(\u0\/u0\/_0001_ ), .B_N(\w3\[16\] ), .Y(\u0\/u0\/_0205_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0764_ ( .A(\u0\/u0\/_0205_ ), .X(\u0\/u0\/_0216_ ) );
sky130_fd_sc_hd__and3_1 \u0/u0/_0765_ ( .A(\u0\/u0\/_0162_ ), .B(\u0\/u0\/_0194_ ), .C(\u0\/u0\/_0216_ ), .X(\u0\/u0\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \u0/u0/_0766_ ( .A(\u0\/u0\/_0183_ ), .SLEEP(\u0\/u0\/_0227_ ), .X(\u0\/u0\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u0/_0767_ ( .A(\w3\[16\] ), .B_N(\u0\/u0\/_0001_ ), .Y(\u0\/u0\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_0768_ ( .A(\w3\[18\] ), .B(\w3\[19\] ), .Y(\u0\/u0\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0769_ ( .A(\u0\/u0\/_0249_ ), .B(\u0\/u0\/_0260_ ), .X(\u0\/u0\/_0271_ ) );
sky130_fd_sc_hd__buf_2 \u0/u0/_0771_ ( .A(\u0\/u0\/_0271_ ), .X(\u0\/u0\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0772_ ( .A(\u0\/u0\/_0162_ ), .X(\u0\/u0\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_0773_ ( .A(\u0\/u0\/_0293_ ), .B(\u0\/u0\/_0304_ ), .Y(\u0\/u0\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \u0/u0/_0774_ ( .A(\u0\/u0\/_0001_ ), .Y(\u0\/u0\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \u0/u0/_0776_ ( .A(\w3\[16\] ), .Y(\u0\/u0\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0777_ ( .A(\w3\[18\] ), .B(\w3\[19\] ), .X(\u0\/u0\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0779_ ( .A(\u0\/u0\/_0358_ ), .X(\u0\/u0\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_0780_ ( .A1(\u0\/u0\/_0325_ ), .A2(\u0\/u0\/_0347_ ), .B1(\u0\/u0\/_0380_ ), .C1(\u0\/u0\/_0304_ ), .Y(\u0\/u0\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u0/_0781_ ( .A_N(\u0\/u0\/_0238_ ), .B(\u0\/u0\/_0314_ ), .C(\u0\/u0\/_0391_ ), .X(\u0\/u0\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u0/_0782_ ( .A(\w3\[19\] ), .B_N(\w3\[18\] ), .Y(\u0\/u0\/_0412_ ) );
sky130_fd_sc_hd__buf_2 \u0/u0/_0783_ ( .A(\u0\/u0\/_0412_ ), .X(\u0\/u0\/_0423_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0784_ ( .A(\u0\/u0\/_0423_ ), .B(\u0\/u0\/_0205_ ), .X(\u0\/u0\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u0/_0787_ ( .A(\w3\[21\] ), .B_N(\w3\[20\] ), .Y(\u0\/u0\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0788_ ( .A(\u0\/u0\/_0467_ ), .B(\u0\/u0\/_0140_ ), .X(\u0\/u0\/_0478_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_0791_ ( .A(\u0\/u0\/_0134_ ), .B(\u0\/u0\/_0218_ ), .Y(\u0\/u0\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_0792_ ( .A(\u0\/u0\/_0478_ ), .B(\u0\/u0\/_0271_ ), .Y(\u0\/u0\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0793_ ( .A(\u0\/u0\/_0194_ ), .X(\u0\/u0\/_0532_ ) );
sky130_fd_sc_hd__buf_2 \u0/u0/_0794_ ( .A(\u0\/u0\/_0249_ ), .X(\u0\/u0\/_0543_ ) );
sky130_fd_sc_hd__and2_1 \u0/u0/_0795_ ( .A(\u0\/u0\/_0543_ ), .B(\u0\/u0\/_0358_ ), .X(\u0\/u0\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0797_ ( .A(\u0\/u0\/_0554_ ), .X(\u0\/u0\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \u0/u0/_0798_ ( .A(\u0\/u0\/_0216_ ), .B(\u0\/u0\/_0358_ ), .X(\u0\/u0\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0800_ ( .A(\u0\/u0\/_0586_ ), .X(\u0\/u0\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_0801_ ( .A1(\u0\/u0\/_0532_ ), .A2(\u0\/u0\/_0575_ ), .A3(\u0\/u0\/_0608_ ), .B1(\u0\/u0\/_0218_ ), .Y(\u0\/u0\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_0802_ ( .A(\u0\/u0\/_0401_ ), .B(\u0\/u0\/_0510_ ), .C(\u0\/u0\/_0521_ ), .D(\u0\/u0\/_0619_ ), .X(\u0\/u0\/_0629_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0803_ ( .A(\u0\/u0\/_0358_ ), .B(\u0\/u0\/_0001_ ), .X(\u0\/u0\/_0640_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0804_ ( .A(\u0\/u0\/_0640_ ), .X(\u0\/u0\/_0651_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0805_ ( .A(\u0\/u0\/_0205_ ), .B(\u0\/u0\/_0260_ ), .X(\u0\/u0\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0806_ ( .A(\u0\/u0\/_0662_ ), .X(\u0\/u0\/_0672_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0807_ ( .A(\u0\/u0\/_0672_ ), .X(\u0\/u0\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u0/_0808_ ( .A(\w3\[22\] ), .B_N(\w3\[23\] ), .Y(\u0\/u0\/_0694_ ) );
sky130_fd_sc_hd__and2_2 \u0/u0/_0809_ ( .A(\u0\/u0\/_0467_ ), .B(\u0\/u0\/_0694_ ), .X(\u0\/u0\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0811_ ( .A(\u0\/u0\/_0705_ ), .X(\u0\/u0\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_0812_ ( .A1(\u0\/u0\/_0651_ ), .A2(\u0\/u0\/_0293_ ), .A3(\u0\/u0\/_0683_ ), .B1(\u0\/u0\/_0727_ ), .Y(\u0\/u0\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_0813_ ( .A(\u0\/u0\/_0001_ ), .B(\w3\[16\] ), .Y(\u0\/u0\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0814_ ( .A(\u0\/u0\/_0730_ ), .B(\u0\/u0\/_0260_ ), .X(\u0\/u0\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0815_ ( .A(\u0\/u0\/_0731_ ), .X(\u0\/u0\/_0732_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0816_ ( .A(\u0\/u0\/_0732_ ), .X(\u0\/u0\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0817_ ( .A(\w3\[16\] ), .X(\u0\/u0\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u0/_0818_ ( .A1(\u0\/u0\/_0325_ ), .A2(\u0\/u0\/_0734_ ), .B1(\u0\/u0\/_0423_ ), .X(\u0\/u0\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0819_ ( .A(\u0\/u0\/_0694_ ), .B(\u0\/u0\/_0151_ ), .X(\u0\/u0\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0821_ ( .A(\u0\/u0\/_0736_ ), .X(\u0\/u0\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0822_ ( .A(\u0\/u0\/_0738_ ), .X(\u0\/u0\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_0823_ ( .A1(\u0\/u0\/_0733_ ), .A2(\u0\/u0\/_0735_ ), .A3(\u0\/u0\/_0293_ ), .B1(\u0\/u0\/_0739_ ), .Y(\u0\/u0\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u0/_0824_ ( .A(\u0\/u0\/_0730_ ), .B_N(\u0\/u0\/_0358_ ), .Y(\u0\/u0\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_0825_ ( .A(\u0\/u0\/_0741_ ), .B(\u0\/u0\/_0739_ ), .Y(\u0\/u0\/_0742_ ) );
sky130_fd_sc_hd__buf_2 \u0/u0/_0826_ ( .A(\u0\/u0\/_0118_ ), .X(\u0\/u0\/_0743_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_0827_ ( .A1(\u0\/u0\/_0743_ ), .A2(\u0\/u0\/_0216_ ), .B1(\u0\/u0\/_0532_ ), .C1(\u0\/u0\/_0739_ ), .Y(\u0\/u0\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_0828_ ( .A(\u0\/u0\/_0729_ ), .B(\u0\/u0\/_0740_ ), .C(\u0\/u0\/_0742_ ), .D(\u0\/u0\/_0744_ ), .X(\u0\/u0\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0829_ ( .A(\u0\/u0\/_0423_ ), .B(\u0\/u0\/_0730_ ), .X(\u0\/u0\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0830_ ( .A(\u0\/u0\/_0746_ ), .X(\u0\/u0\/_0747_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0831_ ( .A(\u0\/u0\/_0747_ ), .X(\u0\/u0\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u0/_0832_ ( .A(\w3\[20\] ), .B_N(\w3\[21\] ), .Y(\u0\/u0\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0833_ ( .A(\u0\/u0\/_0749_ ), .B(\u0\/u0\/_0694_ ), .X(\u0\/u0\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0835_ ( .A(\u0\/u0\/_0750_ ), .X(\u0\/u0\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0836_ ( .A(\u0\/u0\/_0752_ ), .X(\u0\/u0\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0837_ ( .A(\u0\/u0\/_0118_ ), .B(\u0\/u0\/_0358_ ), .X(\u0\/u0\/_0017_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0838_ ( .A(\u0\/u0\/_0017_ ), .X(\u0\/u0\/_0018_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0839_ ( .A(\u0\/u0\/_0752_ ), .B(\u0\/u0\/_0018_ ), .X(\u0\/u0\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0840_ ( .A(\u0\/u0\/_0358_ ), .B(\u0\/u0\/_0325_ ), .X(\u0\/u0\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0842_ ( .A(\u0\/u0\/_0096_ ), .B(\u0\/u0\/_0205_ ), .X(\u0\/u0\/_0022_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0843_ ( .A(\u0\/u0\/_0022_ ), .X(\u0\/u0\/_0023_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u0/_0844_ ( .A1(\u0\/u0\/_0020_ ), .A2(\u0\/u0\/_0023_ ), .B1(\u0\/u0\/_0752_ ), .X(\u0\/u0\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_0845_ ( .A1(\u0\/u0\/_0748_ ), .A2(\u0\/u0\/_0016_ ), .B1(\u0\/u0\/_0019_ ), .C1(\u0\/u0\/_0024_ ), .Y(\u0\/u0\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \u0/u0/_0846_ ( .A(\w3\[20\] ), .B(\w3\[21\] ), .X(\u0\/u0\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0847_ ( .A(\u0\/u0\/_0694_ ), .B(\u0\/u0\/_0026_ ), .X(\u0\/u0\/_0027_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0850_ ( .A(\u0\/u0\/_0358_ ), .B(\u0\/u0\/_0730_ ), .X(\u0\/u0\/_0030_ ) );
sky130_fd_sc_hd__buf_2 \u0/u0/_0852_ ( .A(\u0\/u0\/_0030_ ), .X(\u0\/u0\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_0853_ ( .A(\u0\/u0\/_0247_ ), .B(\u0\/u0\/_0032_ ), .Y(\u0\/u0\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_0854_ ( .A(\u0\/u0\/_0247_ ), .B(\u0\/u0\/_0735_ ), .Y(\u0\/u0\/_0034_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0855_ ( .A(\u0\/u0\/_0118_ ), .B(\u0\/u0\/_0260_ ), .X(\u0\/u0\/_0035_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0856_ ( .A(\u0\/u0\/_0035_ ), .X(\u0\/u0\/_0036_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0857_ ( .A(\u0\/u0\/_0027_ ), .B(\u0\/u0\/_0036_ ), .X(\u0\/u0\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0858_ ( .A(\u0\/u0\/_0260_ ), .X(\u0\/u0\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_0859_ ( .A(\u0\/u0\/_0038_ ), .B(\u0\/u0\/_0347_ ), .Y(\u0\/u0\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u0/_0860_ ( .A_N(\u0\/u0\/_0039_ ), .B(\u0\/u0\/_0027_ ), .X(\u0\/u0\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_0861_ ( .A(\u0\/u0\/_0037_ ), .B(\u0\/u0\/_0040_ ), .Y(\u0\/u0\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_0862_ ( .A(\u0\/u0\/_0025_ ), .B(\u0\/u0\/_0033_ ), .C(\u0\/u0\/_0034_ ), .D(\u0\/u0\/_0041_ ), .X(\u0\/u0\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0863_ ( .A(\u0\/u0\/_0749_ ), .B(\u0\/u0\/_0140_ ), .X(\u0\/u0\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \u0/u0/_0865_ ( .A(\w3\[16\] ), .B(\w3\[18\] ), .C(\w3\[19\] ), .X(\u0\/u0\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0866_ ( .A(\u0\/u0\/_0043_ ), .B(\u0\/u0\/_0045_ ), .X(\u0\/u0\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0867_ ( .A(\u0\/u0\/_0096_ ), .B(\u0\/u0\/_0543_ ), .X(\u0\/u0\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0869_ ( .A(\u0\/u0\/_0047_ ), .B(\u0\/u0\/_0043_ ), .X(\u0\/u0\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0870_ ( .A(\u0\/u0\/_0730_ ), .X(\u0\/u0\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0871_ ( .A(\u0\/u0\/_0043_ ), .X(\u0\/u0\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_0872_ ( .A1(\u0\/u0\/_0743_ ), .A2(\u0\/u0\/_0050_ ), .B1(\u0\/u0\/_0194_ ), .C1(\u0\/u0\/_0051_ ), .Y(\u0\/u0\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u0/_0873_ ( .A(\u0\/u0\/_0046_ ), .B(\u0\/u0\/_0049_ ), .C_N(\u0\/u0\/_0052_ ), .Y(\u0\/u0\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0874_ ( .A(\u0\/u0\/_0026_ ), .B(\u0\/u0\/_0140_ ), .X(\u0\/u0\/_0054_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0876_ ( .A(\u0\/u0\/_0054_ ), .X(\u0\/u0\/_0056_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_0877_ ( .A1(\u0\/u0\/_0532_ ), .A2(\u0\/u0\/_0575_ ), .B1(\u0\/u0\/_0056_ ), .Y(\u0\/u0\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0878_ ( .A(\u0\/u0\/_0423_ ), .B(\u0\/u0\/_0325_ ), .X(\u0\/u0\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0880_ ( .A(\u0\/u0\/_0051_ ), .X(\u0\/u0\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_0881_ ( .A1(\u0\/u0\/_0732_ ), .A2(\u0\/u0\/_0036_ ), .A3(\u0\/u0\/_0058_ ), .B1(\u0\/u0\/_0060_ ), .Y(\u0\/u0\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0882_ ( .A(\u0\/u0\/_0260_ ), .B(\u0\/u0\/_0001_ ), .X(\u0\/u0\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0884_ ( .A(\u0\/u0\/_0062_ ), .X(\u0\/u0\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_0885_ ( .A1(\u0\/u0\/_0064_ ), .A2(\u0\/u0\/_0748_ ), .A3(\u0\/u0\/_0683_ ), .B1(\u0\/u0\/_0056_ ), .Y(\u0\/u0\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_0886_ ( .A(\u0\/u0\/_0053_ ), .B(\u0\/u0\/_0057_ ), .C(\u0\/u0\/_0061_ ), .D(\u0\/u0\/_0065_ ), .X(\u0\/u0\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_0887_ ( .A(\u0\/u0\/_0629_ ), .B(\u0\/u0\/_0745_ ), .C(\u0\/u0\/_0042_ ), .D(\u0\/u0\/_0066_ ), .X(\u0\/u0\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u0/_0889_ ( .A(\w3\[23\] ), .B_N(\w3\[22\] ), .Y(\u0\/u0\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0890_ ( .A(\u0\/u0\/_0069_ ), .B(\u0\/u0\/_0151_ ), .X(\u0\/u0\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0892_ ( .A(\u0\/u0\/_0070_ ), .X(\u0\/u0\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_0893_ ( .A1(\u0\/u0\/_0129_ ), .A2(\u0\/u0\/_0586_ ), .B1(\u0\/u0\/_0072_ ), .Y(\u0\/u0\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_0894_ ( .A1(\u0\/u0\/_0380_ ), .A2(\u0\/u0\/_0347_ ), .B1(\u0\/u0\/_0194_ ), .B2(\u0\/u0\/_0216_ ), .Y(\u0\/u0\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u0/_0895_ ( .A(\u0\/u0\/_0074_ ), .B_N(\u0\/u0\/_0070_ ), .Y(\u0\/u0\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u0/_0896_ ( .A(\u0\/u0\/_0073_ ), .SLEEP(\u0\/u0\/_0075_ ), .X(\u0\/u0\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \u0/u0/_0897_ ( .A(\u0\/u0\/_0467_ ), .B(\u0\/u0\/_0069_ ), .X(\u0\/u0\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0898_ ( .A(\u0\/u0\/_0077_ ), .X(\u0\/u0\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0899_ ( .A(\u0\/u0\/_0412_ ), .B(\u0\/u0\/_0118_ ), .X(\u0\/u0\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0901_ ( .A(\u0\/u0\/_0078_ ), .B(\u0\/u0\/_0079_ ), .X(\u0\/u0\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0902_ ( .A(\u0\/u0\/_0412_ ), .B(\u0\/u0\/_0249_ ), .X(\u0\/u0\/_0082_ ) );
sky130_fd_sc_hd__buf_2 \u0/u0/_0904_ ( .A(\u0\/u0\/_0082_ ), .X(\u0\/u0\/_0084_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0905_ ( .A(\u0\/u0\/_0084_ ), .B(\u0\/u0\/_0078_ ), .X(\u0\/u0\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u0/_0906_ ( .A1(\w3\[16\] ), .A2(\u0\/u0\/_0325_ ), .B1(\u0\/u0\/_0260_ ), .Y(\u0\/u0\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u0/_0907_ ( .A_N(\u0\/u0\/_0086_ ), .B(\u0\/u0\/_0078_ ), .X(\u0\/u0\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u0/_0908_ ( .A(\u0\/u0\/_0081_ ), .B(\u0\/u0\/_0085_ ), .C(\u0\/u0\/_0087_ ), .Y(\u0\/u0\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0909_ ( .A(\u0\/u0\/_0072_ ), .X(\u0\/u0\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_0910_ ( .A1(\u0\/u0\/_0733_ ), .A2(\u0\/u0\/_0748_ ), .A3(\u0\/u0\/_0683_ ), .B1(\u0\/u0\/_0089_ ), .Y(\u0\/u0\/_0090_ ) );
sky130_fd_sc_hd__buf_2 \u0/u0/_0911_ ( .A(\u0\/u0\/_0129_ ), .X(\u0\/u0\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0912_ ( .A(\u0\/u0\/_0018_ ), .X(\u0\/u0\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0913_ ( .A(\u0\/u0\/_0023_ ), .X(\u0\/u0\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0914_ ( .A(\u0\/u0\/_0078_ ), .X(\u0\/u0\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_0915_ ( .A1(\u0\/u0\/_0091_ ), .A2(\u0\/u0\/_0092_ ), .A3(\u0\/u0\/_0093_ ), .B1(\u0\/u0\/_0094_ ), .Y(\u0\/u0\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_0916_ ( .A(\u0\/u0\/_0076_ ), .B(\u0\/u0\/_0088_ ), .C(\u0\/u0\/_0090_ ), .D(\u0\/u0\/_0095_ ), .X(\u0\/u0\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \u0/u0/_0917_ ( .A(\u0\/u0\/_0069_ ), .B(\u0\/u0\/_0026_ ), .X(\u0\/u0\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \u0/u0/_0918_ ( .A(\u0\/u0\/_0098_ ), .X(\u0\/u0\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0919_ ( .A(\u0\/u0\/_0434_ ), .B(\u0\/u0\/_0099_ ), .X(\u0\/u0\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0920_ ( .A(\u0\/u0\/_0079_ ), .B(\u0\/u0\/_0098_ ), .X(\u0\/u0\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0921_ ( .A(\u0\/u0\/_0325_ ), .X(\u0\/u0\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_0922_ ( .A1(\u0\/u0\/_0102_ ), .A2(\u0\/u0\/_0734_ ), .B1(\u0\/u0\/_0038_ ), .C1(\u0\/u0\/_0099_ ), .Y(\u0\/u0\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u0/_0923_ ( .A(\u0\/u0\/_0100_ ), .B(\u0\/u0\/_0101_ ), .C_N(\u0\/u0\/_0103_ ), .Y(\u0\/u0\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_0924_ ( .A1(\u0\/u0\/_0554_ ), .A2(\u0\/u0\/_0586_ ), .B1(\u0\/u0\/_0099_ ), .Y(\u0\/u0\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_0925_ ( .A(\u0\/u0\/_0129_ ), .B(\u0\/u0\/_0099_ ), .Y(\u0\/u0\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0926_ ( .A(\u0\/u0\/_0105_ ), .B(\u0\/u0\/_0106_ ), .X(\u0\/u0\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0927_ ( .A(\u0\/u0\/_0423_ ), .X(\u0\/u0\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \u0/u0/_0928_ ( .A(\u0\/u0\/_0260_ ), .B(\w3\[16\] ), .X(\u0\/u0\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0929_ ( .A(\u0\/u0\/_0069_ ), .B(\u0\/u0\/_0749_ ), .X(\u0\/u0\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0931_ ( .A(\u0\/u0\/_0111_ ), .X(\u0\/u0\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0932_ ( .A(\u0\/u0\/_0113_ ), .X(\u0\/u0\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_0933_ ( .A1(\u0\/u0\/_0109_ ), .A2(\u0\/u0\/_0110_ ), .B1(\u0\/u0\/_0114_ ), .Y(\u0\/u0\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_0934_ ( .A(\u0\/u0\/_0023_ ), .Y(\u0\/u0\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_0935_ ( .A(\u0\/u0\/_0554_ ), .Y(\u0\/u0\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u0/_0936_ ( .A1(\u0\/u0\/_0050_ ), .A2(\u0\/u0\/_0743_ ), .B1(\u0\/u0\/_0194_ ), .Y(\u0\/u0\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_0937_ ( .A(\u0\/u0\/_0113_ ), .Y(\u0\/u0\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \u0/u0/_0938_ ( .A1(\u0\/u0\/_0116_ ), .A2(\u0\/u0\/_0117_ ), .A3(\u0\/u0\/_0119_ ), .B1(\u0\/u0\/_0120_ ), .X(\u0\/u0\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_0939_ ( .A(\u0\/u0\/_0104_ ), .B(\u0\/u0\/_0108_ ), .C(\u0\/u0\/_0115_ ), .D(\u0\/u0\/_0121_ ), .X(\u0\/u0\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_0940_ ( .A(\w3\[23\] ), .B(\w3\[22\] ), .Y(\u0\/u0\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0941_ ( .A(\u0\/u0\/_0749_ ), .B(\u0\/u0\/_0123_ ), .X(\u0\/u0\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0943_ ( .A(\u0\/u0\/_0082_ ), .B(\u0\/u0\/_0124_ ), .X(\u0\/u0\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_0944_ ( .A(\u0\/u0\/_0271_ ), .B(\u0\/u0\/_0124_ ), .Y(\u0\/u0\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0945_ ( .A(\u0\/u0\/_0124_ ), .X(\u0\/u0\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0946_ ( .A(\u0\/u0\/_0260_ ), .B(\u0\/u0\/_0325_ ), .X(\u0\/u0\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_0948_ ( .A(\u0\/u0\/_0128_ ), .B(\u0\/u0\/_0130_ ), .Y(\u0\/u0\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_0949_ ( .A(\u0\/u0\/_0127_ ), .B(\u0\/u0\/_0132_ ), .Y(\u0\/u0\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \u0/u0/_0950_ ( .A(\u0\/u0\/_0434_ ), .X(\u0\/u0\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_0951_ ( .A(\u0\/u0\/_0134_ ), .B(\u0\/u0\/_0128_ ), .Y(\u0\/u0\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u0/_0952_ ( .A(\u0\/u0\/_0126_ ), .B(\u0\/u0\/_0133_ ), .C_N(\u0\/u0\/_0135_ ), .Y(\u0\/u0\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \u0/u0/_0953_ ( .A(\u0\/u0\/_0026_ ), .B(\u0\/u0\/_0123_ ), .X(\u0\/u0\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0955_ ( .A(\u0\/u0\/_0137_ ), .X(\u0\/u0\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_0956_ ( .A1(\u0\/u0\/_0110_ ), .A2(\u0\/u0\/_0293_ ), .A3(\u0\/u0\/_0084_ ), .B1(\u0\/u0\/_0139_ ), .Y(\u0\/u0\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0957_ ( .A(\u0\/u0\/_0096_ ), .B(\u0\/u0\/_0730_ ), .X(\u0\/u0\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0959_ ( .A(\u0\/u0\/_0142_ ), .X(\u0\/u0\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_0960_ ( .A1(\u0\/u0\/_0020_ ), .A2(\u0\/u0\/_0144_ ), .A3(\u0\/u0\/_0018_ ), .B1(\u0\/u0\/_0139_ ), .Y(\u0\/u0\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u0/_0961_ ( .A(\w3\[18\] ), .B(\u0\/u0\/_0050_ ), .C_N(\w3\[19\] ), .Y(\u0\/u0\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0962_ ( .A(\u0\/u0\/_0128_ ), .X(\u0\/u0\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_0963_ ( .A1(\u0\/u0\/_0146_ ), .A2(\u0\/u0\/_0032_ ), .A3(\u0\/u0\/_0651_ ), .B1(\u0\/u0\/_0147_ ), .Y(\u0\/u0\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_0964_ ( .A(\u0\/u0\/_0136_ ), .B(\u0\/u0\/_0141_ ), .C(\u0\/u0\/_0145_ ), .D(\u0\/u0\/_0148_ ), .X(\u0\/u0\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0965_ ( .A(\u0\/u0\/_0123_ ), .B(\u0\/u0\/_0151_ ), .X(\u0\/u0\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_0967_ ( .A(\u0\/u0\/_0150_ ), .X(\u0\/u0\/_0153_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0968_ ( .A(\u0\/u0\/_0150_ ), .B(\u0\/u0\/_0062_ ), .X(\u0\/u0\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_0969_ ( .A(\u0\/u0\/_0079_ ), .B(\u0\/u0\/_0150_ ), .Y(\u0\/u0\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u0/_0970_ ( .A(\u0\/u0\/_0150_ ), .B(\u0\/u0\/_0423_ ), .C(\u0\/u0\/_0543_ ), .Y(\u0\/u0\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_0971_ ( .A(\u0\/u0\/_0155_ ), .B(\u0\/u0\/_0156_ ), .Y(\u0\/u0\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_0972_ ( .A1(\u0\/u0\/_0153_ ), .A2(\u0\/u0\/_0134_ ), .B1(\u0\/u0\/_0154_ ), .C1(\u0\/u0\/_0157_ ), .Y(\u0\/u0\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0973_ ( .A(\u0\/u0\/_0467_ ), .B(\u0\/u0\/_0123_ ), .X(\u0\/u0\/_0159_ ) );
sky130_fd_sc_hd__buf_2 \u0/u0/_0975_ ( .A(\u0\/u0\/_0159_ ), .X(\u0\/u0\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u0/_0976_ ( .A_N(\u0\/u0\/_0119_ ), .B(\u0\/u0\/_0161_ ), .X(\u0\/u0\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_0977_ ( .A(\u0\/u0\/_0163_ ), .Y(\u0\/u0\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_0978_ ( .A1(\u0\/u0\/_0146_ ), .A2(\u0\/u0\/_0575_ ), .A3(\u0\/u0\/_0608_ ), .B1(\u0\/u0\/_0153_ ), .Y(\u0\/u0\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_0979_ ( .A1(\u0\/u0\/_0062_ ), .A2(\u0\/u0\/_0084_ ), .A3(\u0\/u0\/_0134_ ), .B1(\u0\/u0\/_0161_ ), .Y(\u0\/u0\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_0980_ ( .A(\u0\/u0\/_0158_ ), .B(\u0\/u0\/_0164_ ), .C(\u0\/u0\/_0165_ ), .D(\u0\/u0\/_0166_ ), .X(\u0\/u0\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_0981_ ( .A(\u0\/u0\/_0097_ ), .B(\u0\/u0\/_0122_ ), .C(\u0\/u0\/_0149_ ), .D(\u0\/u0\/_0167_ ), .X(\u0\/u0\/_0168_ ) );
sky130_fd_sc_hd__and2_1 \u0/u0/_0982_ ( .A(\u0\/u0\/_0672_ ), .B(\u0\/u0\/_0150_ ), .X(\u0\/u0\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_0983_ ( .A(\u0\/u0\/_0154_ ), .B(\u0\/u0\/_0169_ ), .Y(\u0\/u0\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \u0/u0/_0984_ ( .A(\u0\/u0\/_0123_ ), .B(\u0\/u0\/_0151_ ), .C(\u0\/u0\/_0038_ ), .X(\u0\/u0\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0985_ ( .A(\u0\/u0\/_0170_ ), .B(\u0\/u0\/_0171_ ), .X(\u0\/u0\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_0986_ ( .A(\u0\/u0\/_0172_ ), .Y(\u0\/u0\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u0/_0987_ ( .A(\u0\/u0\/_0067_ ), .B(\u0\/u0\/_0168_ ), .C(\u0\/u0\/_0174_ ), .Y(\u0\/u0\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/u0/_0988_ ( .A(\u0\/u0\/_0001_ ), .B(\w3\[16\] ), .Y(\u0\/u0\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \u0/u0/_0989_ ( .A(\u0\/u0\/_0175_ ), .B(\u0\/u0\/_0358_ ), .X(\u0\/u0\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0990_ ( .A(\u0\/u0\/_0176_ ), .B(\u0\/u0\/_0478_ ), .X(\u0\/u0\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_0991_ ( .A(\u0\/u0\/_0084_ ), .B(\u0\/u0\/_0113_ ), .Y(\u0\/u0\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0992_ ( .A(\u0\/u0\/_0111_ ), .B(\u0\/u0\/_0062_ ), .X(\u0\/u0\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0993_ ( .A(\u0\/u0\/_0111_ ), .B(\u0\/u0\/_0672_ ), .X(\u0\/u0\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_0994_ ( .A(\u0\/u0\/_0179_ ), .B(\u0\/u0\/_0180_ ), .Y(\u0\/u0\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0995_ ( .A(\u0\/u0\/_0054_ ), .B(\u0\/u0\/_0058_ ), .X(\u0\/u0\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_0996_ ( .A(\u0\/u0\/_0182_ ), .Y(\u0\/u0\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u0/_0997_ ( .A_N(\u0\/u0\/_0177_ ), .B(\u0\/u0\/_0178_ ), .C(\u0\/u0\/_0181_ ), .D(\u0\/u0\/_0184_ ), .X(\u0\/u0\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0998_ ( .A(\u0\/u0\/_0098_ ), .B(\u0\/u0\/_0741_ ), .X(\u0\/u0\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_0999_ ( .A(\u0\/u0\/_0047_ ), .B(\u0\/u0\/_0098_ ), .X(\u0\/u0\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \u0/u0/_1000_ ( .A(\u0\/u0\/_0186_ ), .B(\u0\/u0\/_0187_ ), .X(\u0\/u0\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1001_ ( .A(\u0\/u0\/_0188_ ), .Y(\u0\/u0\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1002_ ( .A(\u0\/u0\/_0738_ ), .B(\u0\/u0\/_0735_ ), .X(\u0\/u0\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1003_ ( .A(\u0\/u0\/_0271_ ), .B(\u0\/u0\/_0736_ ), .X(\u0\/u0\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_1004_ ( .A(\u0\/u0\/_0190_ ), .B(\u0\/u0\/_0191_ ), .Y(\u0\/u0\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \u0/u0/_1005_ ( .A(\u0\/u0\/_0096_ ), .B(\u0\/u0\/_0325_ ), .X(\u0\/u0\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1006_ ( .A1(\u0\/u0\/_0193_ ), .A2(\u0\/u0\/_0176_ ), .B1(\u0\/u0\/_0043_ ), .Y(\u0\/u0\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1007_ ( .A(\u0\/u0\/_0185_ ), .B(\u0\/u0\/_0189_ ), .C(\u0\/u0\/_0192_ ), .D(\u0\/u0\/_0195_ ), .X(\u0\/u0\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u0/_1008_ ( .A_N(\w3\[19\] ), .B(\u0\/u0\/_0734_ ), .C(\w3\[18\] ), .X(\u0\/u0\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1009_ ( .A(\u0\/u0\/_0137_ ), .B(\u0\/u0\/_0197_ ), .X(\u0\/u0\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_1010_ ( .A(\u0\/u0\/_0198_ ), .B(\u0\/u0\/_0040_ ), .Y(\u0\/u0\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1011_ ( .A(\u0\/u0\/_0293_ ), .B(\u0\/u0\/_0137_ ), .X(\u0\/u0\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1012_ ( .A(\u0\/u0\/_0200_ ), .Y(\u0\/u0\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1013_ ( .A(\u0\/u0\/_0137_ ), .B(\u0\/u0\/_0110_ ), .Y(\u0\/u0\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1014_ ( .A(\u0\/u0\/_0139_ ), .B(\u0\/u0\/_0020_ ), .Y(\u0\/u0\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1015_ ( .A(\u0\/u0\/_0199_ ), .B(\u0\/u0\/_0201_ ), .C(\u0\/u0\/_0202_ ), .D(\u0\/u0\/_0203_ ), .X(\u0\/u0\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u0/_1016_ ( .A1(\u0\/u0\/_0532_ ), .A2(\u0\/u0\/_0109_ ), .B1(\u0\/u0\/_0102_ ), .C1(\u0\/u0\/_0727_ ), .X(\u0\/u0\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1017_ ( .A(\u0\/u0\/_0023_ ), .B(\u0\/u0\/_0078_ ), .Y(\u0\/u0\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1018_ ( .A(\u0\/u0\/_0078_ ), .B(\u0\/u0\/_0142_ ), .Y(\u0\/u0\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1019_ ( .A(\u0\/u0\/_0207_ ), .B(\u0\/u0\/_0208_ ), .Y(\u0\/u0\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1020_ ( .A1(\u0\/u0\/_0094_ ), .A2(\u0\/u0\/_0176_ ), .B1(\u0\/u0\/_0206_ ), .C1(\u0\/u0\/_0209_ ), .Y(\u0\/u0\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1021_ ( .A(\u0\/u0\/_0662_ ), .B(\u0\/u0\/_0070_ ), .X(\u0\/u0\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u0/_1022_ ( .A(\u0\/u0\/_0732_ ), .B(\u0\/u0\/_0123_ ), .C(\u0\/u0\/_0749_ ), .Y(\u0\/u0\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u0/_1023_ ( .A(\u0\/u0\/_0732_ ), .B(\u0\/u0\/_0467_ ), .C(\u0\/u0\/_0069_ ), .Y(\u0\/u0\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u0/_1024_ ( .A_N(\u0\/u0\/_0211_ ), .B(\u0\/u0\/_0127_ ), .C(\u0\/u0\/_0212_ ), .D(\u0\/u0\/_0213_ ), .X(\u0\/u0\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1025_ ( .A(\u0\/u0\/_0137_ ), .Y(\u0\/u0\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1026_ ( .A(\u0\/u0\/_0128_ ), .B(\u0\/u0\/_0036_ ), .Y(\u0\/u0\/_0217_ ) );
sky130_fd_sc_hd__buf_2 \u0/u0/_1027_ ( .A(\u0\/u0\/_0478_ ), .X(\u0\/u0\/_0218_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1028_ ( .A1(\u0\/u0\/_0159_ ), .A2(\u0\/u0\/_0747_ ), .B1(\u0\/u0\/_0434_ ), .B2(\u0\/u0\/_0218_ ), .Y(\u0\/u0\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u0/_1029_ ( .A1(\u0\/u0\/_0116_ ), .A2(\u0\/u0\/_0215_ ), .B1(\u0\/u0\/_0217_ ), .C1(\u0\/u0\/_0219_ ), .X(\u0\/u0\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1030_ ( .A(\u0\/u0\/_0113_ ), .B(\u0\/u0\/_0746_ ), .X(\u0\/u0\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u0/_1031_ ( .A1(\u0\/u0\/_0098_ ), .A2(\u0\/u0\/_0746_ ), .B1(\u0\/u0\/_0434_ ), .B2(\u0\/u0\/_0750_ ), .X(\u0\/u0\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1032_ ( .A1(\u0\/u0\/_0047_ ), .A2(\u0\/u0\/_0113_ ), .B1(\u0\/u0\/_0221_ ), .C1(\u0\/u0\/_0222_ ), .Y(\u0\/u0\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u0/_1033_ ( .A1(\u0\/u0\/_0129_ ), .A2(\u0\/u0\/_0162_ ), .B1(\u0\/u0\/_0271_ ), .B2(\u0\/u0\/_0705_ ), .X(\u0\/u0\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1034_ ( .A1(\u0\/u0\/_0093_ ), .A2(\u0\/u0\/_0738_ ), .B1(\u0\/u0\/_0081_ ), .C1(\u0\/u0\/_0224_ ), .Y(\u0\/u0\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1035_ ( .A(\u0\/u0\/_0214_ ), .B(\u0\/u0\/_0220_ ), .C(\u0\/u0\/_0223_ ), .D(\u0\/u0\/_0225_ ), .X(\u0\/u0\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1036_ ( .A(\u0\/u0\/_0196_ ), .B(\u0\/u0\/_0204_ ), .C(\u0\/u0\/_0210_ ), .D(\u0\/u0\/_0226_ ), .X(\u0\/u0\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1037_ ( .A(\u0\/u0\/_0111_ ), .B(\u0\/u0\/_0554_ ), .X(\u0\/u0\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1038_ ( .A(\u0\/u0\/_0229_ ), .Y(\u0\/u0\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1039_ ( .A(\u0\/u0\/_0111_ ), .B(\u0\/u0\/_0129_ ), .Y(\u0\/u0\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1040_ ( .A(\u0\/u0\/_0018_ ), .B(\u0\/u0\/_0738_ ), .Y(\u0\/u0\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1041_ ( .A(\u0\/u0\/_0030_ ), .B(\u0\/u0\/_0304_ ), .Y(\u0\/u0\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1042_ ( .A(\u0\/u0\/_0230_ ), .B(\u0\/u0\/_0231_ ), .C(\u0\/u0\/_0232_ ), .D(\u0\/u0\/_0233_ ), .X(\u0\/u0\/_0234_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1043_ ( .A(\u0\/u0\/_0047_ ), .B(\u0\/u0\/_0478_ ), .X(\u0\/u0\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1044_ ( .A1(\u0\/u0\/_0129_ ), .A2(\u0\/u0\/_0554_ ), .B1(\u0\/u0\/_0137_ ), .Y(\u0\/u0\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u0/_1045_ ( .A(\u0\/u0\/_0235_ ), .B(\u0\/u0\/_0049_ ), .C_N(\u0\/u0\/_0236_ ), .Y(\u0\/u0\/_0237_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1046_ ( .A(\u0\/u0\/_0047_ ), .B(\u0\/u0\/_0077_ ), .X(\u0\/u0\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1047_ ( .A(\u0\/u0\/_0070_ ), .B(\u0\/u0\/_0036_ ), .X(\u0\/u0\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u0/_1048_ ( .A1(\u0\/u0\/_0047_ ), .A2(\u0\/u0\/_0736_ ), .B1(\u0\/u0\/_0023_ ), .B2(\u0\/u0\/_0099_ ), .X(\u0\/u0\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u0/_1049_ ( .A(\u0\/u0\/_0239_ ), .B(\u0\/u0\/_0240_ ), .C(\u0\/u0\/_0241_ ), .Y(\u0\/u0\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1050_ ( .A(\u0\/u0\/_0554_ ), .B(\u0\/u0\/_0072_ ), .X(\u0\/u0\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u0/_1051_ ( .A1(\u0\/u0\/_0142_ ), .A2(\u0\/u0\/_0137_ ), .B1(\u0\/u0\/_0159_ ), .B2(\u0\/u0\/_0082_ ), .X(\u0\/u0\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1052_ ( .A1(\u0\/u0\/_0608_ ), .A2(\u0\/u0\/_0072_ ), .B1(\u0\/u0\/_0243_ ), .C1(\u0\/u0\/_0244_ ), .Y(\u0\/u0\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1053_ ( .A(\u0\/u0\/_0234_ ), .B(\u0\/u0\/_0237_ ), .C(\u0\/u0\/_0242_ ), .D(\u0\/u0\/_0245_ ), .X(\u0\/u0\/_0246_ ) );
sky130_fd_sc_hd__buf_2 \u0/u0/_1054_ ( .A(\u0\/u0\/_0027_ ), .X(\u0\/u0\/_0247_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u0/_1055_ ( .A1(\u0\/u0\/_0554_ ), .A2(\u0\/u0\/_0586_ ), .B1(\u0\/u0\/_0247_ ), .X(\u0\/u0\/_0248_ ) );
sky130_fd_sc_hd__and2_1 \u0/u0/_1056_ ( .A(\u0\/u0\/_0082_ ), .B(\u0\/u0\/_0478_ ), .X(\u0\/u0\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_1057_ ( .A(\u0\/u0\/_0079_ ), .X(\u0\/u0\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1058_ ( .A(\u0\/u0\/_0251_ ), .B(\u0\/u0\/_0478_ ), .X(\u0\/u0\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_1059_ ( .A(\u0\/u0\/_0250_ ), .B(\u0\/u0\/_0252_ ), .Y(\u0\/u0\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1060_ ( .A(\u0\/u0\/_0016_ ), .B(\u0\/u0\/_0064_ ), .Y(\u0\/u0\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_1061_ ( .A(\u0\/u0\/_0304_ ), .X(\u0\/u0\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1062_ ( .A(\u0\/u0\/_0255_ ), .B(\u0\/u0\/_0651_ ), .Y(\u0\/u0\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u0/_1063_ ( .A_N(\u0\/u0\/_0248_ ), .B(\u0\/u0\/_0253_ ), .C(\u0\/u0\/_0254_ ), .D(\u0\/u0\/_0256_ ), .X(\u0\/u0\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1064_ ( .A(\u0\/u0\/_0099_ ), .B(\u0\/u0\/_0110_ ), .X(\u0\/u0\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \u0/u0/_1065_ ( .A1(\u0\/u0\/_0161_ ), .A2(\u0\/u0\/_0130_ ), .B1(\u0\/u0\/_0258_ ), .Y(\u0\/u0\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1066_ ( .A(\u0\/u0\/_0194_ ), .B(\u0\/u0\/_0001_ ), .X(\u0\/u0\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1068_ ( .A(\u0\/u0\/_0261_ ), .B(\u0\/u0\/_0153_ ), .Y(\u0\/u0\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u0/_1069_ ( .A_N(\u0\/u0\/_0154_ ), .B(\u0\/u0\/_0259_ ), .C(\u0\/u0\/_0263_ ), .X(\u0\/u0\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1070_ ( .A(\u0\/u0\/_0246_ ), .B(\u0\/u0\/_0174_ ), .C(\u0\/u0\/_0257_ ), .D(\u0\/u0\/_0264_ ), .X(\u0\/u0\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u0/_1071_ ( .A1(\u0\/u0\/_0261_ ), .A2(\u0\/u0\/_0554_ ), .B1(\u0\/u0\/_0159_ ), .X(\u0\/u0\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1072_ ( .A(\u0\/u0\/_0747_ ), .B(\u0\/u0\/_0150_ ), .Y(\u0\/u0\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1073_ ( .A(\u0\/u0\/_0175_ ), .Y(\u0\/u0\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \u0/u0/_1074_ ( .A(\u0\/u0\/_0423_ ), .B(\u0\/u0\/_0123_ ), .C(\u0\/u0\/_0151_ ), .X(\u0\/u0\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1075_ ( .A(\u0\/u0\/_0268_ ), .B(\u0\/u0\/_0269_ ), .Y(\u0\/u0\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u0/_1076_ ( .A_N(\u0\/u0\/_0266_ ), .B(\u0\/u0\/_0267_ ), .C(\u0\/u0\/_0270_ ), .X(\u0\/u0\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1077_ ( .A(\u0\/u0\/_0554_ ), .B(\u0\/u0\/_0150_ ), .X(\u0\/u0\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1078_ ( .A(\u0\/u0\/_0273_ ), .Y(\u0\/u0\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1079_ ( .A1(\u0\/u0\/_0734_ ), .A2(\u0\/u0\/_0325_ ), .B1(\u0\/u0\/_0380_ ), .Y(\u0\/u0\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1080_ ( .A(\u0\/u0\/_0275_ ), .Y(\u0\/u0\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1081_ ( .A(\u0\/u0\/_0276_ ), .B(\u0\/u0\/_0153_ ), .Y(\u0\/u0\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \u0/u0/_1082_ ( .A(\u0\/u0\/_0272_ ), .B(\u0\/u0\/_0274_ ), .C(\u0\/u0\/_0277_ ), .X(\u0\/u0\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_1083_ ( .A(\u0\/u0\/_0036_ ), .X(\u0\/u0\/_0279_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1085_ ( .A1(\u0\/u0\/_0218_ ), .A2(\u0\/u0\/_0279_ ), .B1(\u0\/u0\/_0084_ ), .B2(\u0\/u0\/_0060_ ), .Y(\u0\/u0\/_0281_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u0/_1086_ ( .A1(\u0\/u0\/_0251_ ), .A2(\u0\/u0\/_0434_ ), .B1(\u0\/u0\/_0304_ ), .Y(\u0\/u0\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1087_ ( .A(\u0\/u0\/_0091_ ), .B(\u0\/u0\/_0056_ ), .Y(\u0\/u0\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1088_ ( .A1(\u0\/u0\/_0743_ ), .A2(\u0\/u0\/_0050_ ), .B1(\u0\/u0\/_0038_ ), .C1(\u0\/u0\/_0255_ ), .Y(\u0\/u0\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1089_ ( .A(\u0\/u0\/_0281_ ), .B(\u0\/u0\/_0283_ ), .C(\u0\/u0\/_0284_ ), .D(\u0\/u0\/_0285_ ), .X(\u0\/u0\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1090_ ( .A(\u0\/u0\/_0082_ ), .B(\u0\/u0\/_0027_ ), .X(\u0\/u0\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1091_ ( .A(\u0\/u0\/_0129_ ), .B(\u0\/u0\/_0027_ ), .X(\u0\/u0\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_1092_ ( .A(\u0\/u0\/_0287_ ), .B(\u0\/u0\/_0288_ ), .Y(\u0\/u0\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1093_ ( .A1(\u0\/u0\/_0752_ ), .A2(\u0\/u0\/_0683_ ), .B1(\u0\/u0\/_0093_ ), .B2(\u0\/u0\/_0247_ ), .Y(\u0\/u0\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1094_ ( .A1(\u0\/u0\/_0092_ ), .A2(\u0\/u0\/_0575_ ), .B1(\u0\/u0\/_0056_ ), .Y(\u0\/u0\/_0291_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1096_ ( .A1(\u0\/u0\/_0218_ ), .A2(\u0\/u0\/_0672_ ), .B1(\u0\/u0\/_0084_ ), .B2(\u0\/u0\/_0056_ ), .Y(\u0\/u0\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1097_ ( .A(\u0\/u0\/_0289_ ), .B(\u0\/u0\/_0290_ ), .C(\u0\/u0\/_0291_ ), .D(\u0\/u0\/_0294_ ), .X(\u0\/u0\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1098_ ( .A(\u0\/u0\/_0750_ ), .B(\u0\/u0\/_0193_ ), .X(\u0\/u0\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1099_ ( .A(\u0\/u0\/_0705_ ), .B(\u0\/u0\/_0380_ ), .X(\u0\/u0\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1100_ ( .A(\u0\/u0\/_0752_ ), .B(\u0\/u0\/_0129_ ), .Y(\u0\/u0\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u0/_1101_ ( .A(\u0\/u0\/_0296_ ), .B(\u0\/u0\/_0297_ ), .C_N(\u0\/u0\/_0298_ ), .Y(\u0\/u0\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1102_ ( .A(\u0\/u0\/_0089_ ), .B(\u0\/u0\/_0532_ ), .Y(\u0\/u0\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1103_ ( .A(\w3\[18\] ), .Y(\u0\/u0\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u0/_1104_ ( .A(\u0\/u0\/_0301_ ), .B(\w3\[19\] ), .C(\u0\/u0\/_0743_ ), .Y(\u0\/u0\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1105_ ( .A(\u0\/u0\/_0072_ ), .B(\u0\/u0\/_0302_ ), .X(\u0\/u0\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1106_ ( .A(\u0\/u0\/_0303_ ), .Y(\u0\/u0\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1107_ ( .A(\u0\/u0\/_0147_ ), .B(\u0\/u0\/_0302_ ), .Y(\u0\/u0\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1108_ ( .A(\u0\/u0\/_0299_ ), .B(\u0\/u0\/_0300_ ), .C(\u0\/u0\/_0305_ ), .D(\u0\/u0\/_0306_ ), .X(\u0\/u0\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1109_ ( .A(\u0\/u0\/_0278_ ), .B(\u0\/u0\/_0286_ ), .C(\u0\/u0\/_0295_ ), .D(\u0\/u0\/_0307_ ), .X(\u0\/u0\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u0/_1110_ ( .A(\u0\/u0\/_0228_ ), .B(\u0\/u0\/_0265_ ), .C(\u0\/u0\/_0308_ ), .Y(\u0\/u0\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1111_ ( .A(\u0\/u0\/_0235_ ), .Y(\u0\/u0\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1112_ ( .A(\u0\/u0\/_0478_ ), .B(\u0\/u0\/_0640_ ), .X(\u0\/u0\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1113_ ( .A(\u0\/u0\/_0310_ ), .Y(\u0\/u0\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1114_ ( .A(\u0\/u0\/_0023_ ), .B(\u0\/u0\/_0218_ ), .Y(\u0\/u0\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1115_ ( .A(\u0\/u0\/_0218_ ), .B(\u0\/u0\/_0032_ ), .Y(\u0\/u0\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1116_ ( .A(\u0\/u0\/_0309_ ), .B(\u0\/u0\/_0311_ ), .C(\u0\/u0\/_0312_ ), .D(\u0\/u0\/_0313_ ), .X(\u0\/u0\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1117_ ( .A(\u0\/u0\/_0218_ ), .B(\u0\/u0\/_0064_ ), .Y(\u0\/u0\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1118_ ( .A(\u0\/u0\/_0218_ ), .B(\u0\/u0\/_0683_ ), .Y(\u0\/u0\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1119_ ( .A(\u0\/u0\/_0315_ ), .B(\u0\/u0\/_0316_ ), .C(\u0\/u0\/_0317_ ), .D(\u0\/u0\/_0253_ ), .X(\u0\/u0\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1120_ ( .A(\u0\/u0\/_0047_ ), .B(\u0\/u0\/_0304_ ), .Y(\u0\/u0\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1121_ ( .A(\u0\/u0\/_0586_ ), .B(\u0\/u0\/_0162_ ), .Y(\u0\/u0\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1122_ ( .A(\u0\/u0\/_0319_ ), .B(\u0\/u0\/_0320_ ), .Y(\u0\/u0\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_1123_ ( .A(\u0\/u0\/_0321_ ), .B(\u0\/u0\/_0238_ ), .Y(\u0\/u0\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1124_ ( .A(\u0\/u0\/_0304_ ), .B(\u0\/u0\/_0062_ ), .Y(\u0\/u0\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_1125_ ( .A(\u0\/u0\/_0251_ ), .X(\u0\/u0\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1126_ ( .A1(\u0\/u0\/_0324_ ), .A2(\u0\/u0\/_0084_ ), .B1(\u0\/u0\/_0255_ ), .Y(\u0\/u0\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1127_ ( .A1(\u0\/u0\/_0050_ ), .A2(\u0\/u0\/_0216_ ), .B1(\u0\/u0\/_0109_ ), .C1(\u0\/u0\/_0255_ ), .Y(\u0\/u0\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1128_ ( .A(\u0\/u0\/_0322_ ), .B(\u0\/u0\/_0323_ ), .C(\u0\/u0\/_0326_ ), .D(\u0\/u0\/_0327_ ), .X(\u0\/u0\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1129_ ( .A1(\u0\/u0\/_0733_ ), .A2(\u0\/u0\/_0279_ ), .A3(\u0\/u0\/_0058_ ), .B1(\u0\/u0\/_0056_ ), .Y(\u0\/u0\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_1130_ ( .A(\u0\/u0\/_0047_ ), .X(\u0\/u0\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1131_ ( .A(\u0\/u0\/_0330_ ), .B(\u0\/u0\/_0056_ ), .Y(\u0\/u0\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1132_ ( .A(\u0\/u0\/_0054_ ), .B(\u0\/u0\/_0045_ ), .Y(\u0\/u0\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1133_ ( .A(\u0\/u0\/_0329_ ), .B(\u0\/u0\/_0331_ ), .C(\u0\/u0\/_0284_ ), .D(\u0\/u0\/_0332_ ), .X(\u0\/u0\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u0/_1134_ ( .A1(\u0\/u0\/_0543_ ), .A2(\u0\/u0\/_0216_ ), .B1(\u0\/u0\/_0532_ ), .C1(\u0\/u0\/_0060_ ), .X(\u0\/u0\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1135_ ( .A(\u0\/u0\/_0084_ ), .B(\u0\/u0\/_0060_ ), .Y(\u0\/u0\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1136_ ( .A(\u0\/u0\/_0324_ ), .B(\u0\/u0\/_0060_ ), .Y(\u0\/u0\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1137_ ( .A(\u0\/u0\/_0335_ ), .B(\u0\/u0\/_0337_ ), .Y(\u0\/u0\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1138_ ( .A1(\u0\/u0\/_0276_ ), .A2(\u0\/u0\/_0060_ ), .B1(\u0\/u0\/_0334_ ), .C1(\u0\/u0\/_0338_ ), .Y(\u0\/u0\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1139_ ( .A(\u0\/u0\/_0318_ ), .B(\u0\/u0\/_0328_ ), .C(\u0\/u0\/_0333_ ), .D(\u0\/u0\/_0339_ ), .X(\u0\/u0\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u0/_1140_ ( .A1(\u0\/u0\/_0747_ ), .A2(\u0\/u0\/_0134_ ), .B1(\u0\/u0\/_0128_ ), .X(\u0\/u0\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u0/_1141_ ( .A_N(\u0\/u0\/_0086_ ), .B(\u0\/u0\/_0128_ ), .X(\u0\/u0\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1142_ ( .A(\u0\/u0\/_0079_ ), .B(\u0\/u0\/_0124_ ), .X(\u0\/u0\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_1143_ ( .A(\u0\/u0\/_0126_ ), .B(\u0\/u0\/_0343_ ), .Y(\u0\/u0\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u0/_1144_ ( .A(\u0\/u0\/_0341_ ), .B(\u0\/u0\/_0342_ ), .C_N(\u0\/u0\/_0344_ ), .Y(\u0\/u0\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1146_ ( .A1(\u0\/u0\/_0193_ ), .A2(\u0\/u0\/_0092_ ), .A3(\u0\/u0\/_0330_ ), .B1(\u0\/u0\/_0147_ ), .Y(\u0\/u0\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1147_ ( .A1(\u0\/u0\/_0130_ ), .A2(\u0\/u0\/_0084_ ), .A3(\u0\/u0\/_0134_ ), .B1(\u0\/u0\/_0139_ ), .Y(\u0\/u0\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1148_ ( .A1(\u0\/u0\/_0144_ ), .A2(\u0\/u0\/_0608_ ), .A3(\u0\/u0\/_0092_ ), .B1(\u0\/u0\/_0139_ ), .Y(\u0\/u0\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1149_ ( .A(\u0\/u0\/_0345_ ), .B(\u0\/u0\/_0348_ ), .C(\u0\/u0\/_0349_ ), .D(\u0\/u0\/_0350_ ), .X(\u0\/u0\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \u0/u0/_1150_ ( .A(\u0\/u0\/_0150_ ), .B(\u0\/u0\/_0194_ ), .C(\u0\/u0\/_0543_ ), .X(\u0\/u0\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u0/_1151_ ( .A(\u0\/u0\/_0277_ ), .SLEEP(\u0\/u0\/_0352_ ), .X(\u0\/u0\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \u0/u0/_1152_ ( .A1(\u0\/u0\/_0268_ ), .A2(\u0\/u0\/_0171_ ), .B1(\u0\/u0\/_0157_ ), .Y(\u0\/u0\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u0/_1153_ ( .A(\u0\/u0\/_0161_ ), .X(\u0\/u0\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1154_ ( .A1(\u0\/u0\/_0279_ ), .A2(\u0\/u0\/_0084_ ), .B1(\u0\/u0\/_0355_ ), .Y(\u0\/u0\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1155_ ( .A1(\u0\/u0\/_0020_ ), .A2(\u0\/u0\/_0193_ ), .A3(\u0\/u0\/_0091_ ), .B1(\u0\/u0\/_0355_ ), .Y(\u0\/u0\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1156_ ( .A(\u0\/u0\/_0353_ ), .B(\u0\/u0\/_0354_ ), .C(\u0\/u0\/_0356_ ), .D(\u0\/u0\/_0357_ ), .X(\u0\/u0\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1157_ ( .A(\u0\/u0\/_0111_ ), .B(\u0\/u0\/_0586_ ), .X(\u0\/u0\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1158_ ( .A(\u0\/u0\/_0360_ ), .Y(\u0\/u0\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u0/_1159_ ( .A1(\u0\/u0\/_0119_ ), .A2(\u0\/u0\/_0120_ ), .B1(\u0\/u0\/_0230_ ), .C1(\u0\/u0\/_0361_ ), .X(\u0\/u0\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1160_ ( .A1(\u0\/u0\/_0672_ ), .A2(\u0\/u0\/_0251_ ), .A3(\u0\/u0\/_0134_ ), .B1(\u0\/u0\/_0114_ ), .Y(\u0\/u0\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1162_ ( .A1(\u0\/u0\/_0036_ ), .A2(\u0\/u0\/_0251_ ), .A3(\u0\/u0\/_0134_ ), .B1(\u0\/u0\/_0099_ ), .Y(\u0\/u0\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1163_ ( .A1(\u0\/u0\/_0193_ ), .A2(\u0\/u0\/_0608_ ), .B1(\u0\/u0\/_0099_ ), .Y(\u0\/u0\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1164_ ( .A(\u0\/u0\/_0362_ ), .B(\u0\/u0\/_0363_ ), .C(\u0\/u0\/_0365_ ), .D(\u0\/u0\/_0366_ ), .X(\u0\/u0\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1165_ ( .A1(\u0\/u0\/_0575_ ), .A2(\u0\/u0\/_0092_ ), .A3(\u0\/u0\/_0330_ ), .B1(\u0\/u0\/_0089_ ), .Y(\u0\/u0\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1166_ ( .A1(\u0\/u0\/_0586_ ), .A2(\u0\/u0\/_0018_ ), .A3(\u0\/u0\/_0330_ ), .B1(\u0\/u0\/_0094_ ), .Y(\u0\/u0\/_0370_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1167_ ( .A1(\u0\/u0\/_0293_ ), .A2(\u0\/u0\/_0134_ ), .B1(\u0\/u0\/_0089_ ), .Y(\u0\/u0\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1168_ ( .A1(\u0\/u0\/_0279_ ), .A2(\u0\/u0\/_0134_ ), .B1(\u0\/u0\/_0094_ ), .Y(\u0\/u0\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1169_ ( .A(\u0\/u0\/_0368_ ), .B(\u0\/u0\/_0370_ ), .C(\u0\/u0\/_0371_ ), .D(\u0\/u0\/_0372_ ), .X(\u0\/u0\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1170_ ( .A(\u0\/u0\/_0351_ ), .B(\u0\/u0\/_0359_ ), .C(\u0\/u0\/_0367_ ), .D(\u0\/u0\/_0373_ ), .X(\u0\/u0\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1171_ ( .A1(\u0\/u0\/_0102_ ), .A2(\u0\/u0\/_0347_ ), .B1(\u0\/u0\/_0109_ ), .C1(\u0\/u0\/_0247_ ), .Y(\u0\/u0\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1172_ ( .A1(\u0\/u0\/_0102_ ), .A2(\u0\/u0\/_0347_ ), .B1(\u0\/u0\/_0532_ ), .C1(\u0\/u0\/_0247_ ), .Y(\u0\/u0\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1173_ ( .A1(\u0\/u0\/_0050_ ), .A2(\u0\/u0\/_0543_ ), .B1(\u0\/u0\/_0380_ ), .C1(\u0\/u0\/_0247_ ), .Y(\u0\/u0\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1174_ ( .A(\u0\/u0\/_0041_ ), .B(\u0\/u0\/_0375_ ), .C(\u0\/u0\/_0376_ ), .D(\u0\/u0\/_0377_ ), .X(\u0\/u0\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1175_ ( .A(\u0\/u0\/_0047_ ), .B(\u0\/u0\/_0750_ ), .X(\u0\/u0\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1176_ ( .A(\u0\/u0\/_0379_ ), .Y(\u0\/u0\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1177_ ( .A(\u0\/u0\/_0016_ ), .B(\u0\/u0\/_0608_ ), .Y(\u0\/u0\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1178_ ( .A(\u0\/u0\/_0752_ ), .B(\u0\/u0\/_0554_ ), .Y(\u0\/u0\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1179_ ( .A1(\u0\/u0\/_0001_ ), .A2(\u0\/u0\/_0734_ ), .B1(\u0\/u0\/_0109_ ), .C1(\u0\/u0\/_0016_ ), .Y(\u0\/u0\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1180_ ( .A(\u0\/u0\/_0381_ ), .B(\u0\/u0\/_0382_ ), .C(\u0\/u0\/_0383_ ), .D(\u0\/u0\/_0384_ ), .X(\u0\/u0\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \u0/u0/_1181_ ( .A(\u0\/u0\/_0086_ ), .B_N(\u0\/u0\/_0736_ ), .X(\u0\/u0\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1182_ ( .A1(\u0\/u0\/_0748_ ), .A2(\u0\/u0\/_0134_ ), .B1(\u0\/u0\/_0739_ ), .Y(\u0\/u0\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1183_ ( .A1(\u0\/u0\/_0743_ ), .A2(\u0\/u0\/_0543_ ), .B1(\u0\/u0\/_0109_ ), .C1(\u0\/u0\/_0739_ ), .Y(\u0\/u0\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1184_ ( .A1(\u0\/u0\/_0102_ ), .A2(\u0\/u0\/_0301_ ), .B1(\w3\[19\] ), .C1(\u0\/u0\/_0739_ ), .Y(\u0\/u0\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1185_ ( .A(\u0\/u0\/_0386_ ), .B(\u0\/u0\/_0387_ ), .C(\u0\/u0\/_0388_ ), .D(\u0\/u0\/_0389_ ), .X(\u0\/u0\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1186_ ( .A(\u0\/u0\/_0020_ ), .Y(\u0\/u0\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1187_ ( .A(\u0\/u0\/_0727_ ), .Y(\u0\/u0\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1188_ ( .A(\u0\/u0\/_0727_ ), .B(\u0\/u0\/_0064_ ), .Y(\u0\/u0\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1189_ ( .A1(\u0\/u0\/_0102_ ), .A2(\u0\/u0\/_0734_ ), .B1(\u0\/u0\/_0532_ ), .C1(\u0\/u0\/_0727_ ), .Y(\u0\/u0\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u0/_1190_ ( .A1(\u0\/u0\/_0392_ ), .A2(\u0\/u0\/_0393_ ), .B1(\u0\/u0\/_0394_ ), .C1(\u0\/u0\/_0395_ ), .X(\u0\/u0\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1191_ ( .A(\u0\/u0\/_0378_ ), .B(\u0\/u0\/_0385_ ), .C(\u0\/u0\/_0390_ ), .D(\u0\/u0\/_0396_ ), .X(\u0\/u0\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u0/_1192_ ( .A(\u0\/u0\/_0340_ ), .B(\u0\/u0\/_0374_ ), .C(\u0\/u0\/_0397_ ), .Y(\u0\/u0\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1193_ ( .A(\u0\/u0\/_0077_ ), .B(\u0\/u0\/_0129_ ), .X(\u0\/u0\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_1194_ ( .A(\u0\/u0\/_0398_ ), .B(\u0\/u0\/_0239_ ), .Y(\u0\/u0\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1195_ ( .A(\u0\/u0\/_0023_ ), .B(\u0\/u0\/_0111_ ), .X(\u0\/u0\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u0/_1196_ ( .A_N(\u0\/u0\/_0400_ ), .B(\u0\/u0\/_0231_ ), .Y(\u0\/u0\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u0/_1197_ ( .A(\u0\/u0\/_0399_ ), .SLEEP(\u0\/u0\/_0402_ ), .X(\u0\/u0\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_1198_ ( .A(\u0\/u0\/_0747_ ), .B(\u0\/u0\/_0251_ ), .Y(\u0\/u0\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u0/_1199_ ( .A_N(\u0\/u0\/_0404_ ), .B(\u0\/u0\/_0752_ ), .Y(\u0\/u0\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \u0/u0/_1200_ ( .A(\u0\/u0\/_0467_ ), .B(\u0\/u0\/_0194_ ), .C(\u0\/u0\/_0694_ ), .X(\u0\/u0\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u0/_1201_ ( .A_N(\u0\/u0\/_0175_ ), .B(\u0\/u0\/_0406_ ), .X(\u0\/u0\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1202_ ( .A(\u0\/u0\/_0407_ ), .Y(\u0\/u0\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1203_ ( .A1(\u0\/u0\/_0094_ ), .A2(\u0\/u0\/_0197_ ), .B1(\u0\/u0\/_0114_ ), .B2(\u0\/u0\/_0651_ ), .Y(\u0\/u0\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1204_ ( .A(\u0\/u0\/_0403_ ), .B(\u0\/u0\/_0405_ ), .C(\u0\/u0\/_0408_ ), .D(\u0\/u0\/_0409_ ), .X(\u0\/u0\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1205_ ( .A(\u0\/u0\/_0030_ ), .B(\u0\/u0\/_0150_ ), .Y(\u0\/u0\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u0/_1206_ ( .A_N(\u0\/u0\/_0169_ ), .B(\u0\/u0\/_0289_ ), .C(\u0\/u0\/_0411_ ), .X(\u0\/u0\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u0/_1207_ ( .A1(\u0\/u0\/_0467_ ), .A2(\u0\/u0\/_0151_ ), .B1(\u0\/u0\/_0140_ ), .C1(\u0\/u0\/_0129_ ), .X(\u0\/u0\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1208_ ( .A1(\u0\/u0\/_0608_ ), .A2(\u0\/u0\/_0099_ ), .B1(\u0\/u0\/_0037_ ), .C1(\u0\/u0\/_0414_ ), .Y(\u0\/u0\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1209_ ( .A(\u0\/u0\/_0738_ ), .Y(\u0\/u0\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1210_ ( .A(\u0\/u0\/_0586_ ), .B(\u0\/u0\/_0736_ ), .Y(\u0\/u0\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1211_ ( .A1(\u0\/u0\/_0194_ ), .A2(\u0\/u0\/_0038_ ), .B1(\u0\/u0\/_0743_ ), .C1(\u0\/u0\/_0153_ ), .Y(\u0\/u0\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u0/_1212_ ( .A1(\u0\/u0\/_0416_ ), .A2(\u0\/u0\/_0117_ ), .B1(\u0\/u0\/_0417_ ), .C1(\u0\/u0\/_0418_ ), .X(\u0\/u0\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1213_ ( .A(\u0\/u0\/_0077_ ), .B(\u0\/u0\/_0035_ ), .X(\u0\/u0\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1214_ ( .A(\u0\/u0\/_0672_ ), .B(\u0\/u0\/_0124_ ), .Y(\u0\/u0\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1215_ ( .A(\u0\/u0\/_0030_ ), .B(\u0\/u0\/_0137_ ), .Y(\u0\/u0\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1216_ ( .A(\u0\/u0\/_0072_ ), .B(\u0\/u0\/_0732_ ), .Y(\u0\/u0\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u0/_1217_ ( .A_N(\u0\/u0\/_0420_ ), .B(\u0\/u0\/_0421_ ), .C(\u0\/u0\/_0422_ ), .D(\u0\/u0\/_0424_ ), .X(\u0\/u0\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1218_ ( .A(\u0\/u0\/_0413_ ), .B(\u0\/u0\/_0415_ ), .C(\u0\/u0\/_0419_ ), .D(\u0\/u0\/_0425_ ), .X(\u0\/u0\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u0/_1219_ ( .A(\u0\/u0\/_0355_ ), .B(\u0\/u0\/_0102_ ), .C(\u0\/u0\/_0109_ ), .Y(\u0\/u0\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1220_ ( .A(\u0\/u0\/_0077_ ), .B(\u0\/u0\/_0018_ ), .X(\u0\/u0\/_0428_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1221_ ( .A(\u0\/u0\/_0077_ ), .B(\u0\/u0\/_0554_ ), .X(\u0\/u0\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u0/_1222_ ( .A1(\u0\/u0\/_0050_ ), .A2(\u0\/u0\/_0216_ ), .B1(\u0\/u0\/_0380_ ), .C1(\u0\/u0\/_0078_ ), .X(\u0\/u0\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u0/_1223_ ( .A(\u0\/u0\/_0428_ ), .B(\u0\/u0\/_0429_ ), .C(\u0\/u0\/_0430_ ), .Y(\u0\/u0\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u0/_1224_ ( .A_N(\u0\/u0\/_0209_ ), .B(\u0\/u0\/_0431_ ), .X(\u0\/u0\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u0/_1225_ ( .A1(\u0\/u0\/_0215_ ), .A2(\u0\/u0\/_0404_ ), .B1(\u0\/u0\/_0427_ ), .C1(\u0\/u0\/_0432_ ), .X(\u0\/u0\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1226_ ( .A(\u0\/u0\/_0043_ ), .B(\u0\/u0\/_0058_ ), .Y(\u0\/u0\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1227_ ( .A(\u0\/u0\/_0195_ ), .B(\u0\/u0\/_0233_ ), .C(\u0\/u0\/_0320_ ), .D(\u0\/u0\/_0435_ ), .X(\u0\/u0\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1228_ ( .A(\u0\/u0\/_0261_ ), .B(\u0\/u0\/_0738_ ), .Y(\u0\/u0\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1229_ ( .A1(\u0\/u0\/_0218_ ), .A2(\u0\/u0\/_0651_ ), .B1(\u0\/u0\/_0261_ ), .B2(\u0\/u0\/_0056_ ), .Y(\u0\/u0\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1230_ ( .A(\u0\/u0\/_0436_ ), .B(\u0\/u0\/_0394_ ), .C(\u0\/u0\/_0437_ ), .D(\u0\/u0\/_0438_ ), .X(\u0\/u0\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1231_ ( .A(\u0\/u0\/_0410_ ), .B(\u0\/u0\/_0426_ ), .C(\u0\/u0\/_0433_ ), .D(\u0\/u0\/_0439_ ), .X(\u0\/u0\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u0/_1232_ ( .A(\u0\/u0\/_0135_ ), .SLEEP(\u0\/u0\/_0273_ ), .X(\u0\/u0\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1233_ ( .A1(\u0\/u0\/_0279_ ), .A2(\u0\/u0\/_0134_ ), .B1(\u0\/u0\/_0099_ ), .Y(\u0\/u0\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1234_ ( .A(\u0\/u0\/_0441_ ), .B(\u0\/u0\/_0164_ ), .C(\u0\/u0\/_0270_ ), .D(\u0\/u0\/_0442_ ), .X(\u0\/u0\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1235_ ( .A(\u0\/u0\/_0051_ ), .B(\u0\/u0\/_0672_ ), .Y(\u0\/u0\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1236_ ( .A(\u0\/u0\/_0051_ ), .B(\u0\/u0\/_0271_ ), .Y(\u0\/u0\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1237_ ( .A(\u0\/u0\/_0444_ ), .B(\u0\/u0\/_0446_ ), .X(\u0\/u0\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1238_ ( .A(\u0\/u0\/_0193_ ), .B(\u0\/u0\/_0304_ ), .X(\u0\/u0\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1239_ ( .A(\u0\/u0\/_0448_ ), .Y(\u0\/u0\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1240_ ( .A(\u0\/u0\/_0162_ ), .B(\u0\/u0\/_0130_ ), .X(\u0\/u0\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1241_ ( .A(\u0\/u0\/_0450_ ), .Y(\u0\/u0\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1242_ ( .A1(\u0\/u0\/_0129_ ), .A2(\u0\/u0\/_0554_ ), .B1(\u0\/u0\/_0043_ ), .Y(\u0\/u0\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1243_ ( .A(\u0\/u0\/_0447_ ), .B(\u0\/u0\/_0449_ ), .C(\u0\/u0\/_0451_ ), .D(\u0\/u0\/_0452_ ), .X(\u0\/u0\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1244_ ( .A(\u0\/u0\/_0056_ ), .B(\u0\/u0\/_0064_ ), .Y(\u0\/u0\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u0/_1245_ ( .A_N(\u0\/u0\/_0248_ ), .B(\u0\/u0\/_0454_ ), .C(\u0\/u0\/_0254_ ), .D(\u0\/u0\/_0256_ ), .X(\u0\/u0\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1246_ ( .A1(\u0\/u0\/_0330_ ), .A2(\u0\/u0\/_0099_ ), .B1(\u0\/u0\/_0134_ ), .B2(\u0\/u0\/_0705_ ), .Y(\u0\/u0\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1247_ ( .A1(\u0\/u0\/_0748_ ), .A2(\u0\/u0\/_0738_ ), .B1(\u0\/u0\/_0092_ ), .B2(\u0\/u0\/_0752_ ), .Y(\u0\/u0\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1248_ ( .A1(\u0\/u0\/_0072_ ), .A2(\u0\/u0\/_0036_ ), .B1(\u0\/u0\/_0748_ ), .B2(\u0\/u0\/_0056_ ), .Y(\u0\/u0\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1249_ ( .A1(\u0\/u0\/_0748_ ), .A2(\u0\/u0\/_0251_ ), .B1(\u0\/u0\/_0247_ ), .Y(\u0\/u0\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1250_ ( .A(\u0\/u0\/_0457_ ), .B(\u0\/u0\/_0458_ ), .C(\u0\/u0\/_0459_ ), .D(\u0\/u0\/_0460_ ), .X(\u0\/u0\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1251_ ( .A(\u0\/u0\/_0443_ ), .B(\u0\/u0\/_0453_ ), .C(\u0\/u0\/_0455_ ), .D(\u0\/u0\/_0461_ ), .X(\u0\/u0\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1252_ ( .A(\u0\/u0\/_0705_ ), .B(\u0\/u0\/_0079_ ), .X(\u0\/u0\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1253_ ( .A(\u0\/u0\/_0586_ ), .B(\u0\/u0\/_0124_ ), .Y(\u0\/u0\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1254_ ( .A(\u0\/u0\/_0218_ ), .B(\u0\/u0\/_0747_ ), .Y(\u0\/u0\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u0/_1255_ ( .A_N(\u0\/u0\/_0463_ ), .B(\u0\/u0\/_0464_ ), .C(\u0\/u0\/_0465_ ), .X(\u0\/u0\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u0/_1256_ ( .A1(\u0\/u0\/_0271_ ), .A2(\u0\/u0\/_0072_ ), .B1(\u0\/u0\/_0142_ ), .B2(\u0\/u0\/_0027_ ), .X(\u0\/u0\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1257_ ( .A1(\u0\/u0\/_0144_ ), .A2(\u0\/u0\/_0099_ ), .B1(\u0\/u0\/_0360_ ), .C1(\u0\/u0\/_0468_ ), .Y(\u0\/u0\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u0/_1258_ ( .A1(\u0\/u0\/_0672_ ), .A2(\u0\/u0\/_0251_ ), .B1(\u0\/u0\/_0218_ ), .X(\u0\/u0\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1259_ ( .A1(\u0\/u0\/_0575_ ), .A2(\u0\/u0\/_0056_ ), .B1(\u0\/u0\/_0379_ ), .C1(\u0\/u0\/_0470_ ), .Y(\u0\/u0\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1260_ ( .A(\u0\/u0\/_0466_ ), .B(\u0\/u0\/_0469_ ), .C(\u0\/u0\/_0471_ ), .D(\u0\/u0\/_0305_ ), .X(\u0\/u0\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u0/_1261_ ( .A1(\u0\/u0\/_0247_ ), .A2(\u0\/u0\/_0683_ ), .B1(\u0\/u0\/_0324_ ), .B2(\u0\/u0\/_0056_ ), .X(\u0\/u0\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1262_ ( .A(\u0\/u0\/_0084_ ), .B(\u0\/u0\/_0099_ ), .X(\u0\/u0\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \u0/u0/_1263_ ( .A1(\u0\/u0\/_0092_ ), .A2(\u0\/u0\/_0247_ ), .B1(\u0\/u0\/_0474_ ), .X(\u0\/u0\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u0/_1264_ ( .A(\u0\/u0\/_0075_ ), .B(\u0\/u0\/_0473_ ), .C(\u0\/u0\/_0475_ ), .Y(\u0\/u0\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1265_ ( .A1(\u0\/u0\/_0279_ ), .A2(\u0\/u0\/_0255_ ), .B1(\u0\/u0\/_0084_ ), .B2(\u0\/u0\/_0060_ ), .Y(\u0\/u0\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1266_ ( .A1(\u0\/u0\/_0093_ ), .A2(\u0\/u0\/_0056_ ), .B1(\u0\/u0\/_0134_ ), .B2(\u0\/u0\/_0114_ ), .Y(\u0\/u0\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1267_ ( .A1(\u0\/u0\/_0161_ ), .A2(\u0\/u0\/_0032_ ), .B1(\u0\/u0\/_0324_ ), .B2(\u0\/u0\/_0147_ ), .Y(\u0\/u0\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1268_ ( .A1(\u0\/u0\/_0054_ ), .A2(\u0\/u0\/_0732_ ), .B1(\u0\/u0\/_0748_ ), .B2(\u0\/u0\/_0304_ ), .Y(\u0\/u0\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1269_ ( .A(\u0\/u0\/_0477_ ), .B(\u0\/u0\/_0479_ ), .C(\u0\/u0\/_0480_ ), .D(\u0\/u0\/_0481_ ), .X(\u0\/u0\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1270_ ( .A(\u0\/u0\/_0161_ ), .B(\u0\/u0\/_0064_ ), .Y(\u0\/u0\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u0/_1271_ ( .A(\u0\/u0\/_0732_ ), .B(\u0\/u0\/_0123_ ), .C(\u0\/u0\/_0467_ ), .Y(\u0\/u0\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1272_ ( .A(\u0\/u0\/_0483_ ), .B(\u0\/u0\/_0484_ ), .Y(\u0\/u0\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1273_ ( .A(\u0\/u0\/_0297_ ), .Y(\u0\/u0\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u0/_1274_ ( .A_N(\u0\/u0\/_0485_ ), .B(\u0\/u0\/_0181_ ), .C(\u0\/u0\/_0486_ ), .D(\u0\/u0\/_0386_ ), .X(\u0\/u0\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1275_ ( .A(\u0\/u0\/_0472_ ), .B(\u0\/u0\/_0476_ ), .C(\u0\/u0\/_0482_ ), .D(\u0\/u0\/_0487_ ), .X(\u0\/u0\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u0/_1276_ ( .A(\u0\/u0\/_0440_ ), .B(\u0\/u0\/_0462_ ), .C(\u0\/u0\/_0488_ ), .Y(\u0\/u0\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1277_ ( .A(\u0\/u0\/_0403_ ), .B(\u0\/u0\/_0230_ ), .C(\u0\/u0\/_0451_ ), .D(\u0\/u0\/_0361_ ), .X(\u0\/u0\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1278_ ( .A1(\u0\/u0\/_0743_ ), .A2(\u0\/u0\/_0050_ ), .B1(\u0\/u0\/_0109_ ), .C1(\u0\/u0\/_0139_ ), .Y(\u0\/u0\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1279_ ( .A(\u0\/u0\/_0447_ ), .B(\u0\/u0\/_0437_ ), .C(\u0\/u0\/_0491_ ), .D(\u0\/u0\/_0427_ ), .X(\u0\/u0\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1280_ ( .A1(\u0\/u0\/_0084_ ), .A2(\u0\/u0\/_0255_ ), .B1(\u0\/u0\/_0608_ ), .B2(\u0\/u0\/_0247_ ), .Y(\u0\/u0\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1281_ ( .A1(\u0\/u0\/_0144_ ), .A2(\u0\/u0\/_0147_ ), .B1(\u0\/u0\/_0355_ ), .B2(\u0\/u0\/_0093_ ), .Y(\u0\/u0\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1282_ ( .A1(\u0\/u0\/_0705_ ), .A2(\u0\/u0\/_0279_ ), .B1(\u0\/u0\/_0330_ ), .B2(\u0\/u0\/_0247_ ), .Y(\u0\/u0\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1283_ ( .A1(\u0\/u0\/_0279_ ), .A2(\u0\/u0\/_0084_ ), .B1(\u0\/u0\/_0114_ ), .Y(\u0\/u0\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1284_ ( .A(\u0\/u0\/_0493_ ), .B(\u0\/u0\/_0494_ ), .C(\u0\/u0\/_0495_ ), .D(\u0\/u0\/_0496_ ), .X(\u0\/u0\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1285_ ( .A1(\u0\/u0\/_0134_ ), .A2(\u0\/u0\/_0137_ ), .B1(\u0\/u0\/_0355_ ), .B2(\u0\/u0\/_0575_ ), .Y(\u0\/u0\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1286_ ( .A1(\u0\/u0\/_0099_ ), .A2(\u0\/u0\/_0733_ ), .B1(\u0\/u0\/_0093_ ), .B2(\u0\/u0\/_0218_ ), .Y(\u0\/u0\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1287_ ( .A(\u0\/u0\/_0147_ ), .B(\u0\/u0\/_0651_ ), .Y(\u0\/u0\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1288_ ( .A1(\u0\/u0\/_0153_ ), .A2(\u0\/u0\/_0056_ ), .B1(\u0\/u0\/_0748_ ), .Y(\u0\/u0\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1289_ ( .A(\u0\/u0\/_0498_ ), .B(\u0\/u0\/_0500_ ), .C(\u0\/u0\/_0501_ ), .D(\u0\/u0\/_0502_ ), .X(\u0\/u0\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1290_ ( .A(\u0\/u0\/_0490_ ), .B(\u0\/u0\/_0492_ ), .C(\u0\/u0\/_0497_ ), .D(\u0\/u0\/_0503_ ), .X(\u0\/u0\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u0/_1291_ ( .A_N(\u0\/u0\/_0275_ ), .B(\u0\/u0\/_0705_ ), .X(\u0\/u0\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1292_ ( .A(\u0\/u0\/_0505_ ), .Y(\u0\/u0\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1293_ ( .A(\u0\/u0\/_0380_ ), .B(\u0\/u0\/_0347_ ), .X(\u0\/u0\/_0507_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u0/_1294_ ( .A1(\u0\/u0\/_0507_ ), .A2(\u0\/u0\/_0093_ ), .B1(\u0\/u0\/_0056_ ), .Y(\u0\/u0\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1295_ ( .A(\u0\/u0\/_0322_ ), .B(\u0\/u0\/_0277_ ), .C(\u0\/u0\/_0506_ ), .D(\u0\/u0\/_0508_ ), .X(\u0\/u0\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1296_ ( .A(\u0\/u0\/_0084_ ), .B(\u0\/u0\/_0705_ ), .X(\u0\/u0\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1297_ ( .A1(\u0\/u0\/_0733_ ), .A2(\u0\/u0\/_0114_ ), .B1(\u0\/u0\/_0429_ ), .C1(\u0\/u0\/_0511_ ), .Y(\u0\/u0\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_1298_ ( .A(\u0\/u0\/_0019_ ), .B(\u0\/u0\/_0024_ ), .Y(\u0\/u0\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1299_ ( .A(\u0\/u0\/_0512_ ), .B(\u0\/u0\/_0513_ ), .C(\u0\/u0\/_0742_ ), .D(\u0\/u0\/_0306_ ), .X(\u0\/u0\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1300_ ( .A1(\u0\/u0\/_0532_ ), .A2(\u0\/u0\/_0089_ ), .B1(\u0\/u0\/_0154_ ), .C1(\u0\/u0\/_0169_ ), .Y(\u0\/u0\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u0/_1301_ ( .A1(\u0\/u0\/_0749_ ), .A2(\u0\/u0\/_0026_ ), .B1(\u0\/u0\/_0069_ ), .C1(\u0\/u0\/_0032_ ), .X(\u0\/u0\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u0/_1302_ ( .A1(\u0\/u0\/_0324_ ), .A2(\u0\/u0\/_0355_ ), .B1(\u0\/u0\/_0330_ ), .B2(\u0\/u0\/_0727_ ), .X(\u0\/u0\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u0/_1303_ ( .A(\u0\/u0\/_0133_ ), .B(\u0\/u0\/_0516_ ), .C(\u0\/u0\/_0517_ ), .Y(\u0\/u0\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1304_ ( .A(\u0\/u0\/_0509_ ), .B(\u0\/u0\/_0514_ ), .C(\u0\/u0\/_0515_ ), .D(\u0\/u0\/_0518_ ), .X(\u0\/u0\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1305_ ( .A(\u0\/u0\/_0747_ ), .B(\u0\/u0\/_0072_ ), .Y(\u0\/u0\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1306_ ( .A1(\u0\/u0\/_0082_ ), .A2(\u0\/u0\/_0070_ ), .B1(\u0\/u0\/_0043_ ), .B2(\u0\/u0\/_0193_ ), .Y(\u0\/u0\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1307_ ( .A(\u0\/u0\/_0311_ ), .B(\u0\/u0\/_0520_ ), .C(\u0\/u0\/_0332_ ), .D(\u0\/u0\/_0522_ ), .X(\u0\/u0\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1308_ ( .A(\u0\/u0\/_0129_ ), .B(\u0\/u0\/_0218_ ), .X(\u0\/u0\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_1309_ ( .A(\u0\/u0\/_0235_ ), .B(\u0\/u0\/_0524_ ), .Y(\u0\/u0\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u0/_1310_ ( .A(\u0\/u0\/_0081_ ), .B(\u0\/u0\/_0085_ ), .Y(\u0\/u0\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1311_ ( .A1(\u0\/u0\/_0051_ ), .A2(\u0\/u0\/_0045_ ), .B1(\u0\/u0\/_0130_ ), .B2(\u0\/u0\/_0094_ ), .Y(\u0\/u0\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1312_ ( .A(\u0\/u0\/_0523_ ), .B(\u0\/u0\/_0525_ ), .C(\u0\/u0\/_0526_ ), .D(\u0\/u0\/_0527_ ), .X(\u0\/u0\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u0/_1313_ ( .A_N(\u0\/u0\/_0250_ ), .B(\u0\/u0\/_0521_ ), .Y(\u0\/u0\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1314_ ( .A(\u0\/u0\/_0128_ ), .B(\u0\/u0\/_0020_ ), .X(\u0\/u0\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1315_ ( .A(\u0\/u0\/_0530_ ), .Y(\u0\/u0\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1316_ ( .A(\u0\/u0\/_0099_ ), .B(\u0\/u0\/_0058_ ), .X(\u0\/u0\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1317_ ( .A(\u0\/u0\/_0533_ ), .Y(\u0\/u0\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u0/_1318_ ( .A_N(\u0\/u0\/_0529_ ), .B(\u0\/u0\/_0531_ ), .C(\u0\/u0\/_0534_ ), .D(\u0\/u0\/_0192_ ), .X(\u0\/u0\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1319_ ( .A(\u0\/u0\/_0434_ ), .B(\u0\/u0\/_0078_ ), .X(\u0\/u0\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u0/_1320_ ( .A1(\u0\/u0\/_0750_ ), .A2(\u0\/u0\/_0079_ ), .B1(\u0\/u0\/_0129_ ), .B2(\u0\/u0\/_0705_ ), .X(\u0\/u0\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1321_ ( .A1(\u0\/u0\/_0161_ ), .A2(\u0\/u0\/_0032_ ), .B1(\u0\/u0\/_0536_ ), .C1(\u0\/u0\/_0537_ ), .Y(\u0\/u0\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u0/_1322_ ( .A1(\u0\/u0\/_0747_ ), .A2(\u0\/u0\/_0162_ ), .B1(\u0\/u0\/_0079_ ), .B2(\u0\/u0\/_0043_ ), .X(\u0\/u0\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1323_ ( .A1(\u0\/u0\/_0093_ ), .A2(\u0\/u0\/_0247_ ), .B1(\u0\/u0\/_0240_ ), .C1(\u0\/u0\/_0539_ ), .Y(\u0\/u0\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1324_ ( .A(\u0\/u0\/_0434_ ), .B(\u0\/u0\/_0043_ ), .X(\u0\/u0\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u0/_1325_ ( .A1(\u0\/u0\/_0142_ ), .A2(\u0\/u0\/_0150_ ), .B1(\u0\/u0\/_0023_ ), .B2(\u0\/u0\/_0137_ ), .X(\u0\/u0\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1326_ ( .A1(\u0\/u0\/_0279_ ), .A2(\u0\/u0\/_0051_ ), .B1(\u0\/u0\/_0541_ ), .C1(\u0\/u0\/_0542_ ), .Y(\u0\/u0\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1327_ ( .A(\u0\/u0\/_0159_ ), .B(\u0\/u0\/_0036_ ), .X(\u0\/u0\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u0/_1328_ ( .A1(\u0\/u0\/_0271_ ), .A2(\u0\/u0\/_0434_ ), .B1(\u0\/u0\/_0027_ ), .X(\u0\/u0\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1329_ ( .A1(\u0\/u0\/_0091_ ), .A2(\u0\/u0\/_0128_ ), .B1(\u0\/u0\/_0545_ ), .C1(\u0\/u0\/_0546_ ), .Y(\u0\/u0\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1330_ ( .A(\u0\/u0\/_0538_ ), .B(\u0\/u0\/_0540_ ), .C(\u0\/u0\/_0544_ ), .D(\u0\/u0\/_0547_ ), .X(\u0\/u0\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1331_ ( .A(\u0\/u0\/_0099_ ), .B(\u0\/u0\/_0193_ ), .X(\u0\/u0\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u0/_1332_ ( .A(\u0\/u0\/_0549_ ), .B(\u0\/u0\/_0186_ ), .C(\u0\/u0\/_0187_ ), .Y(\u0\/u0\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1333_ ( .A(\u0\/u0\/_0062_ ), .B(\u0\/u0\/_0347_ ), .C(\u0\/u0\/_0749_ ), .D(\u0\/u0\/_0694_ ), .X(\u0\/u0\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1334_ ( .A1(\u0\/u0\/_0130_ ), .A2(\u0\/u0\/_0218_ ), .B1(\u0\/u0\/_0551_ ), .C1(\u0\/u0\/_0101_ ), .Y(\u0\/u0\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1335_ ( .A(\u0\/u0\/_0139_ ), .B(\u0\/u0\/_0651_ ), .Y(\u0\/u0\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1336_ ( .A1(\u0\/u0\/_0752_ ), .A2(\u0\/u0\/_0672_ ), .B1(\u0\/u0\/_0084_ ), .B2(\u0\/u0\/_0099_ ), .Y(\u0\/u0\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1337_ ( .A(\u0\/u0\/_0550_ ), .B(\u0\/u0\/_0552_ ), .C(\u0\/u0\/_0553_ ), .D(\u0\/u0\/_0555_ ), .X(\u0\/u0\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1338_ ( .A(\u0\/u0\/_0528_ ), .B(\u0\/u0\/_0535_ ), .C(\u0\/u0\/_0548_ ), .D(\u0\/u0\/_0556_ ), .X(\u0\/u0\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u0/_1339_ ( .A(\u0\/u0\/_0504_ ), .B(\u0\/u0\/_0519_ ), .C(\u0\/u0\/_0557_ ), .Y(\u0\/u0\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1340_ ( .A(\u0\/u0\/_0054_ ), .B(\u0\/u0\/_0507_ ), .X(\u0\/u0\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u0/_1341_ ( .A_N(\u0\/u0\/_0558_ ), .B(\u0\/u0\/_0408_ ), .C(\u0\/u0\/_0451_ ), .D(\u0\/u0\/_0452_ ), .X(\u0\/u0\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1342_ ( .A(\u0\/u0\/_0549_ ), .Y(\u0\/u0\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1343_ ( .A(\u0\/u0\/_0559_ ), .B(\u0\/u0\/_0403_ ), .C(\u0\/u0\/_0560_ ), .D(\u0\/u0\/_0371_ ), .X(\u0\/u0\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1344_ ( .A(\u0\/u0\/_0181_ ), .B(\u0\/u0\/_0178_ ), .X(\u0\/u0\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1345_ ( .A(\u0\/u0\/_0562_ ), .B(\u0\/u0\/_0552_ ), .C(\u0\/u0\/_0553_ ), .D(\u0\/u0\/_0555_ ), .X(\u0\/u0\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1346_ ( .A(\u0\/u0\/_0247_ ), .B(\u0\/u0\/_0020_ ), .Y(\u0\/u0\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1347_ ( .A(\u0\/u0\/_0051_ ), .B(\u0\/u0\/_0130_ ), .X(\u0\/u0\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1348_ ( .A(\u0\/u0\/_0566_ ), .Y(\u0\/u0\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1349_ ( .A(\u0\/u0\/_0159_ ), .B(\u0\/u0\/_0423_ ), .X(\u0\/u0\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1350_ ( .A1(\u0\/u0\/_0752_ ), .A2(\u0\/u0\/_0651_ ), .B1(\u0\/u0\/_0568_ ), .B2(\u0\/u0\/_0175_ ), .Y(\u0\/u0\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1351_ ( .A(\u0\/u0\/_0076_ ), .B(\u0\/u0\/_0565_ ), .C(\u0\/u0\/_0567_ ), .D(\u0\/u0\/_0569_ ), .X(\u0\/u0\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u0/_1352_ ( .A1(\u0\/u0\/_0036_ ), .A2(\u0\/u0\/_0142_ ), .B1(\u0\/u0\/_0161_ ), .X(\u0\/u0\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1353_ ( .A(\u0\/u0\/_0099_ ), .B(\u0\/u0\/_0672_ ), .Y(\u0\/u0\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u0/_1354_ ( .A(\u0\/u0\/_0420_ ), .B(\u0\/u0\/_0571_ ), .C_N(\u0\/u0\/_0572_ ), .Y(\u0\/u0\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1355_ ( .A(\u0\/u0\/_0051_ ), .B(\u0\/u0\/_0747_ ), .Y(\u0\/u0\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1356_ ( .A(\u0\/u0\/_0574_ ), .B(\u0\/u0\/_0319_ ), .C(\u0\/u0\/_0320_ ), .D(\u0\/u0\/_0411_ ), .X(\u0\/u0\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1357_ ( .A(\u0\/u0\/_0736_ ), .B(\u0\/u0\/_0035_ ), .Y(\u0\/u0\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1358_ ( .A(\u0\/u0\/_0736_ ), .B(\u0\/u0\/_0030_ ), .Y(\u0\/u0\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1359_ ( .A(\u0\/u0\/_0298_ ), .B(\u0\/u0\/_0208_ ), .C(\u0\/u0\/_0577_ ), .D(\u0\/u0\/_0578_ ), .X(\u0\/u0\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1360_ ( .A1(\u0\/u0\/_0020_ ), .A2(\u0\/u0\/_0137_ ), .B1(\u0\/u0\/_0261_ ), .B2(\u0\/u0\/_0128_ ), .Y(\u0\/u0\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1361_ ( .A(\u0\/u0\/_0573_ ), .B(\u0\/u0\/_0576_ ), .C(\u0\/u0\/_0579_ ), .D(\u0\/u0\/_0580_ ), .X(\u0\/u0\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1362_ ( .A(\u0\/u0\/_0561_ ), .B(\u0\/u0\/_0563_ ), .C(\u0\/u0\/_0570_ ), .D(\u0\/u0\/_0581_ ), .X(\u0\/u0\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1363_ ( .A(\u0\/u0\/_0128_ ), .B(\u0\/u0\/_0193_ ), .X(\u0\/u0\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1364_ ( .A(\u0\/u0\/_0082_ ), .B(\u0\/u0\/_0162_ ), .X(\u0\/u0\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u0/_1365_ ( .A(\u0\/u0\/_0583_ ), .B(\u0\/u0\/_0584_ ), .C_N(\u0\/u0\/_0437_ ), .Y(\u0\/u0\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u0/_1366_ ( .A(\u0\/u0\/_0150_ ), .B(\u0\/u0\/_0743_ ), .C(\u0\/u0\/_0380_ ), .Y(\u0\/u0\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u0/_1367_ ( .A_N(\u0\/u0\/_0182_ ), .B(\u0\/u0\/_0587_ ), .C(\u0\/u0\/_0323_ ), .X(\u0\/u0\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1368_ ( .A1(\u0\/u0\/_0575_ ), .A2(\u0\/u0\/_0153_ ), .B1(\u0\/u0\/_0727_ ), .B2(\u0\/u0\/_0058_ ), .Y(\u0\/u0\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1369_ ( .A1(\u0\/u0\/_0218_ ), .A2(\u0\/u0\/_0064_ ), .B1(\u0\/u0\/_0134_ ), .B2(\u0\/u0\/_0255_ ), .Y(\u0\/u0\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1370_ ( .A(\u0\/u0\/_0585_ ), .B(\u0\/u0\/_0588_ ), .C(\u0\/u0\/_0589_ ), .D(\u0\/u0\/_0590_ ), .X(\u0\/u0\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \u0/u0/_1371_ ( .A1(\u0\/u0\/_0091_ ), .A2(\u0\/u0\/_0139_ ), .B1(\u0\/u0\/_0250_ ), .Y(\u0\/u0\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1372_ ( .A1(\u0\/u0\/_0092_ ), .A2(\u0\/u0\/_0739_ ), .B1(\u0\/u0\/_0324_ ), .B2(\u0\/u0\/_0247_ ), .Y(\u0\/u0\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1373_ ( .A1(\u0\/u0\/_0144_ ), .A2(\u0\/u0\/_0153_ ), .B1(\u0\/u0\/_0683_ ), .B2(\u0\/u0\/_0056_ ), .Y(\u0\/u0\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1374_ ( .A1(\u0\/u0\/_0091_ ), .A2(\u0\/u0\/_0218_ ), .B1(\u0\/u0\/_0330_ ), .B2(\u0\/u0\/_0056_ ), .Y(\u0\/u0\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1375_ ( .A(\u0\/u0\/_0592_ ), .B(\u0\/u0\/_0593_ ), .C(\u0\/u0\/_0594_ ), .D(\u0\/u0\/_0595_ ), .X(\u0\/u0\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1376_ ( .A(\u0\/u0\/_0218_ ), .B(\u0\/u0\/_0144_ ), .Y(\u0\/u0\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1377_ ( .A(\u0\/u0\/_0312_ ), .B(\u0\/u0\/_0598_ ), .Y(\u0\/u0\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1378_ ( .A(\u0\/u0\/_0575_ ), .B(\u0\/u0\/_0147_ ), .Y(\u0\/u0\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1379_ ( .A1(\u0\/u0\/_0293_ ), .A2(\u0\/u0\/_0137_ ), .B1(\u0\/u0\/_0093_ ), .B2(\u0\/u0\/_0739_ ), .Y(\u0\/u0\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1380_ ( .A1(\u0\/u0\/_0734_ ), .A2(\u0\/u0\/_0531_ ), .B1(\u0\/u0\/_0600_ ), .C1(\u0\/u0\/_0601_ ), .Y(\u0\/u0\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1381_ ( .A1(\u0\/u0\/_0153_ ), .A2(\u0\/u0\/_0261_ ), .B1(\u0\/u0\/_0599_ ), .C1(\u0\/u0\/_0602_ ), .Y(\u0\/u0\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1382_ ( .A(\u0\/u0\/_0591_ ), .B(\u0\/u0\/_0596_ ), .C(\u0\/u0\/_0174_ ), .D(\u0\/u0\/_0603_ ), .X(\u0\/u0\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1383_ ( .A(\u0\/u0\/_0247_ ), .B(\u0\/u0\/_0144_ ), .Y(\u0\/u0\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1384_ ( .A(\u0\/u0\/_0113_ ), .B(\u0\/u0\/_0018_ ), .Y(\u0\/u0\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1385_ ( .A(\u0\/u0\/_0381_ ), .B(\u0\/u0\/_0605_ ), .C(\u0\/u0\/_0361_ ), .D(\u0\/u0\/_0606_ ), .X(\u0\/u0\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1386_ ( .A1(\u0\/u0\/_0016_ ), .A2(\u0\/u0\/_0727_ ), .B1(\u0\/u0\/_0733_ ), .Y(\u0\/u0\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1387_ ( .A1(\u0\/u0\/_0586_ ), .A2(\u0\/u0\/_0159_ ), .B1(\u0\/u0\/_0082_ ), .B2(\u0\/u0\/_0750_ ), .Y(\u0\/u0\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1388_ ( .A1(\u0\/u0\/_0142_ ), .A2(\u0\/u0\/_0162_ ), .B1(\u0\/u0\/_0079_ ), .B2(\u0\/u0\/_0054_ ), .Y(\u0\/u0\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1389_ ( .A(\u0\/u0\/_0610_ ), .B(\u0\/u0\/_0611_ ), .C(\u0\/u0\/_0105_ ), .D(\u0\/u0\/_0106_ ), .X(\u0\/u0\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1390_ ( .A1(\u0\/u0\/_0094_ ), .A2(\u0\/u0\/_0302_ ), .B1(\u0\/u0\/_0324_ ), .B2(\u0\/u0\/_0089_ ), .Y(\u0\/u0\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1391_ ( .A(\u0\/u0\/_0607_ ), .B(\u0\/u0\/_0609_ ), .C(\u0\/u0\/_0612_ ), .D(\u0\/u0\/_0613_ ), .X(\u0\/u0\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1392_ ( .A(\u0\/u0\/_0041_ ), .B(\u0\/u0\/_0170_ ), .X(\u0\/u0\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1393_ ( .A(\u0\/u0\/_0554_ ), .B(\u0\/u0\/_0027_ ), .X(\u0\/u0\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1394_ ( .A(\u0\/u0\/_0027_ ), .B(\u0\/u0\/_0261_ ), .Y(\u0\/u0\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u0/_1395_ ( .A_N(\u0\/u0\/_0616_ ), .B(\u0\/u0\/_0617_ ), .Y(\u0\/u0\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1396_ ( .A1(\u0\/u0\/_0147_ ), .A2(\u0\/u0\/_0302_ ), .B1(\u0\/u0\/_0342_ ), .C1(\u0\/u0\/_0618_ ), .Y(\u0\/u0\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1397_ ( .A(\u0\/u0\/_0614_ ), .B(\u0\/u0\/_0272_ ), .C(\u0\/u0\/_0615_ ), .D(\u0\/u0\/_0620_ ), .X(\u0\/u0\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u0/_1398_ ( .A(\u0\/u0\/_0582_ ), .B(\u0\/u0\/_0604_ ), .C(\u0\/u0\/_0621_ ), .Y(\u0\/u0\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1399_ ( .A1(\u0\/u0\/_0084_ ), .A2(\u0\/u0\/_0134_ ), .B1(\u0\/u0\/_0089_ ), .Y(\u0\/u0\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1400_ ( .A1(\u0\/u0\/_0144_ ), .A2(\u0\/u0\/_0608_ ), .A3(\u0\/u0\/_0330_ ), .B1(\u0\/u0\/_0089_ ), .Y(\u0\/u0\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1401_ ( .A1(\u0\/u0\/_0197_ ), .A2(\u0\/u0\/_0130_ ), .A3(\u0\/u0\/_0110_ ), .B1(\u0\/u0\/_0094_ ), .Y(\u0\/u0\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1402_ ( .A(\u0\/u0\/_0432_ ), .B(\u0\/u0\/_0622_ ), .C(\u0\/u0\/_0623_ ), .D(\u0\/u0\/_0624_ ), .X(\u0\/u0\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \u0/u0/_1403_ ( .A1(\u0\/u0\/_0554_ ), .A2(\u0\/u0\/_0018_ ), .A3(\u0\/u0\/_0023_ ), .B1(\u0\/u0\/_0161_ ), .X(\u0\/u0\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u0/_1404_ ( .A_N(\u0\/u0\/_0269_ ), .B(\u0\/u0\/_0170_ ), .X(\u0\/u0\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1405_ ( .A1(\u0\/u0\/_0109_ ), .A2(\u0\/u0\/_0064_ ), .A3(\u0\/u0\/_0733_ ), .B1(\u0\/u0\/_0355_ ), .Y(\u0\/u0\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u0/_1406_ ( .A_N(\u0\/u0\/_0626_ ), .B(\u0\/u0\/_0627_ ), .C(\u0\/u0\/_0353_ ), .D(\u0\/u0\/_0628_ ), .X(\u0\/u0\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1407_ ( .A1(\u0\/u0\/_0091_ ), .A2(\u0\/u0\/_0110_ ), .A3(\u0\/u0\/_0176_ ), .B1(\u0\/u0\/_0139_ ), .Y(\u0\/u0\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1408_ ( .A1(\u0\/u0\/_0020_ ), .A2(\u0\/u0\/_0261_ ), .B1(\u0\/u0\/_0147_ ), .Y(\u0\/u0\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1409_ ( .A(\u0\/u0\/_0631_ ), .B(\u0\/u0\/_0344_ ), .C(\u0\/u0\/_0421_ ), .D(\u0\/u0\/_0632_ ), .X(\u0\/u0\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u0/_1410_ ( .A1(\u0\/u0\/_0325_ ), .A2(\u0\/u0\/_0734_ ), .B1(\u0\/u0\/_0038_ ), .C1(\u0\/u0\/_0113_ ), .X(\u0\/u0\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1411_ ( .A1(\u0\/u0\/_0134_ ), .A2(\u0\/u0\/_0114_ ), .B1(\u0\/u0\/_0221_ ), .C1(\u0\/u0\/_0634_ ), .Y(\u0\/u0\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u0/_1412_ ( .A(\u0\/u0\/_0119_ ), .B_N(\u0\/u0\/_0111_ ), .Y(\u0\/u0\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1413_ ( .A1(\u0\/u0\/_0032_ ), .A2(\u0\/u0\/_0113_ ), .B1(\u0\/u0\/_0636_ ), .C1(\u0\/u0\/_0400_ ), .Y(\u0\/u0\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1414_ ( .A1(\u0\/u0\/_0732_ ), .A2(\u0\/u0\/_0293_ ), .A3(\u0\/u0\/_0251_ ), .B1(\u0\/u0\/_0099_ ), .Y(\u0\/u0\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1415_ ( .A(\u0\/u0\/_0189_ ), .B(\u0\/u0\/_0635_ ), .C(\u0\/u0\/_0637_ ), .D(\u0\/u0\/_0638_ ), .X(\u0\/u0\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1416_ ( .A(\u0\/u0\/_0625_ ), .B(\u0\/u0\/_0630_ ), .C(\u0\/u0\/_0633_ ), .D(\u0\/u0\/_0639_ ), .X(\u0\/u0\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1417_ ( .A(\u0\/u0\/_0747_ ), .B(\u0\/u0\/_0738_ ), .X(\u0\/u0\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1418_ ( .A(\u0\/u0\/_0736_ ), .B(\u0\/u0\/_0731_ ), .X(\u0\/u0\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u0/_1419_ ( .A_N(\u0\/u0\/_0643_ ), .B(\u0\/u0\/_0577_ ), .Y(\u0\/u0\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1420_ ( .A1(\u0\/u0\/_0084_ ), .A2(\u0\/u0\/_0739_ ), .B1(\u0\/u0\/_0642_ ), .C1(\u0\/u0\/_0644_ ), .Y(\u0\/u0\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1421_ ( .A1(\u0\/u0\/_0050_ ), .A2(\u0\/u0\/_0543_ ), .B1(\u0\/u0\/_0194_ ), .C1(\u0\/u0\/_0738_ ), .Y(\u0\/u0\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1422_ ( .A(\u0\/u0\/_0646_ ), .B(\u0\/u0\/_0232_ ), .C(\u0\/u0\/_0417_ ), .D(\u0\/u0\/_0578_ ), .X(\u0\/u0\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1423_ ( .A1(\u0\/u0\/_0064_ ), .A2(\u0\/u0\/_0733_ ), .B1(\u0\/u0\/_0727_ ), .Y(\u0\/u0\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1424_ ( .A1(\u0\/u0\/_0193_ ), .A2(\u0\/u0\/_0276_ ), .B1(\u0\/u0\/_0727_ ), .Y(\u0\/u0\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1425_ ( .A(\u0\/u0\/_0645_ ), .B(\u0\/u0\/_0647_ ), .C(\u0\/u0\/_0648_ ), .D(\u0\/u0\/_0649_ ), .X(\u0\/u0\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1426_ ( .A1(\u0\/u0\/_0325_ ), .A2(\u0\/u0\/_0734_ ), .B1(\u0\/u0\/_0038_ ), .C1(\u0\/u0\/_0247_ ), .Y(\u0\/u0\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1427_ ( .A1(\u0\/u0\/_0543_ ), .A2(\u0\/u0\/_0216_ ), .B1(\u0\/u0\/_0423_ ), .C1(\u0\/u0\/_0247_ ), .Y(\u0\/u0\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1428_ ( .A(\u0\/u0\/_0652_ ), .B(\u0\/u0\/_0653_ ), .X(\u0\/u0\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1429_ ( .A1(\u0\/u0\/_0733_ ), .A2(\u0\/u0\/_0748_ ), .A3(\u0\/u0\/_0324_ ), .B1(\u0\/u0\/_0016_ ), .Y(\u0\/u0\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1430_ ( .A1(\u0\/u0\/_0651_ ), .A2(\u0\/u0\/_0193_ ), .A3(\u0\/u0\/_0091_ ), .B1(\u0\/u0\/_0016_ ), .Y(\u0\/u0\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1431_ ( .A1(\u0\/u0\/_0102_ ), .A2(\u0\/u0\/_0301_ ), .B1(\w3\[19\] ), .C1(\u0\/u0\/_0247_ ), .Y(\u0\/u0\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1432_ ( .A(\u0\/u0\/_0654_ ), .B(\u0\/u0\/_0655_ ), .C(\u0\/u0\/_0656_ ), .D(\u0\/u0\/_0657_ ), .X(\u0\/u0\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1433_ ( .A1(\u0\/u0\/_0743_ ), .A2(\u0\/u0\/_0050_ ), .B1(\u0\/u0\/_0038_ ), .C1(\u0\/u0\/_0478_ ), .Y(\u0\/u0\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u0/_1434_ ( .A_N(\u0\/u0\/_0250_ ), .B(\u0\/u0\/_0465_ ), .C(\u0\/u0\/_0659_ ), .X(\u0\/u0\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1435_ ( .A1(\u0\/u0\/_0683_ ), .A2(\u0\/u0\/_0324_ ), .B1(\u0\/u0\/_0255_ ), .Y(\u0\/u0\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1436_ ( .A1(\u0\/u0\/_0032_ ), .A2(\u0\/u0\/_0193_ ), .A3(\u0\/u0\/_0047_ ), .B1(\u0\/u0\/_0255_ ), .Y(\u0\/u0\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1437_ ( .A1(\u0\/u0\/_0144_ ), .A2(\u0\/u0\/_0586_ ), .A3(\u0\/u0\/_0047_ ), .B1(\u0\/u0\/_0218_ ), .Y(\u0\/u0\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1438_ ( .A(\u0\/u0\/_0660_ ), .B(\u0\/u0\/_0661_ ), .C(\u0\/u0\/_0663_ ), .D(\u0\/u0\/_0664_ ), .X(\u0\/u0\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1439_ ( .A1(\u0\/u0\/_0091_ ), .A2(\u0\/u0\/_0276_ ), .B1(\u0\/u0\/_0060_ ), .Y(\u0\/u0\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1440_ ( .A1(\u0\/u0\/_0144_ ), .A2(\u0\/u0\/_0608_ ), .B1(\u0\/u0\/_0056_ ), .Y(\u0\/u0\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1441_ ( .A1(\u0\/u0\/_0423_ ), .A2(\u0\/u0\/_0038_ ), .B1(\u0\/u0\/_0102_ ), .C1(\u0\/u0\/_0060_ ), .Y(\u0\/u0\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1442_ ( .A1(\u0\/u0\/_0001_ ), .A2(\u0\/u0\/_0734_ ), .B1(\u0\/u0\/_0109_ ), .C1(\u0\/u0\/_0056_ ), .Y(\u0\/u0\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1443_ ( .A(\u0\/u0\/_0666_ ), .B(\u0\/u0\/_0667_ ), .C(\u0\/u0\/_0668_ ), .D(\u0\/u0\/_0669_ ), .X(\u0\/u0\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1444_ ( .A(\u0\/u0\/_0650_ ), .B(\u0\/u0\/_0658_ ), .C(\u0\/u0\/_0665_ ), .D(\u0\/u0\/_0670_ ), .X(\u0\/u0\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u0/_1445_ ( .A(\u0\/u0\/_0641_ ), .B(\u0\/u0\/_0174_ ), .C(\u0\/u0\/_0671_ ), .Y(\u0\/u0\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u0/_1446_ ( .A(\u0\/u0\/_0049_ ), .B(\u0\/u0\/_0618_ ), .C_N(\u0\/u0\/_0052_ ), .Y(\u0\/u0\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \u0/u0/_1447_ ( .A(\u0\/u0\/_0239_ ), .Y(\u0\/u0\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1448_ ( .A(\u0\/u0\/_0705_ ), .B(\u0\/u0\/_0032_ ), .Y(\u0\/u0\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1449_ ( .A1(\u0\/u0\/_0054_ ), .A2(\u0\/u0\/_0732_ ), .B1(\u0\/u0\/_0036_ ), .B2(\u0\/u0\/_0705_ ), .Y(\u0\/u0\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1450_ ( .A1(\u0\/u0\/_0304_ ), .A2(\u0\/u0\/_0732_ ), .B1(\u0\/u0\/_0047_ ), .B2(\u0\/u0\/_0750_ ), .Y(\u0\/u0\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1451_ ( .A(\u0\/u0\/_0674_ ), .B(\u0\/u0\/_0675_ ), .C(\u0\/u0\/_0676_ ), .D(\u0\/u0\/_0677_ ), .X(\u0\/u0\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u0/_1452_ ( .A_N(\u0\/u0\/_0584_ ), .B(\u0\/u0\/_0283_ ), .X(\u0\/u0\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1453_ ( .A(\u0\/u0\/_0673_ ), .B(\u0\/u0\/_0678_ ), .C(\u0\/u0\/_0679_ ), .D(\u0\/u0\/_0508_ ), .X(\u0\/u0\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1454_ ( .A1(\u0\/u0\/_0016_ ), .A2(\u0\/u0\/_0733_ ), .B1(\u0\/u0\/_0355_ ), .B2(\u0\/u0\/_0092_ ), .Y(\u0\/u0\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1455_ ( .A(\u0\/u0\/_0681_ ), .B(\u0\/u0\/_0034_ ), .X(\u0\/u0\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u0/_1456_ ( .A1(\u0\/u0\/_0330_ ), .A2(\u0\/u0\/_0139_ ), .B1(\u0\/u0\/_0324_ ), .B2(\u0\/u0\/_0089_ ), .X(\u0\/u0\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1457_ ( .A1(\u0\/u0\/_0146_ ), .A2(\u0\/u0\/_0147_ ), .B1(\u0\/u0\/_0133_ ), .C1(\u0\/u0\/_0684_ ), .Y(\u0\/u0\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1458_ ( .A(\u0\/u0\/_0113_ ), .B(\u0\/u0\/_0251_ ), .Y(\u0\/u0\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u0/_1459_ ( .A_N(\u0\/u0\/_0463_ ), .B(\u0\/u0\/_0686_ ), .C(\u0\/u0\/_0383_ ), .D(\u0\/u0\/_0464_ ), .X(\u0\/u0\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1460_ ( .A1(\u0\/u0\/_0051_ ), .A2(\u0\/u0\/_0293_ ), .B1(\u0\/u0\/_0084_ ), .B2(\u0\/u0\/_0705_ ), .Y(\u0\/u0\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1461_ ( .A1(\u0\/u0\/_0018_ ), .A2(\u0\/u0\/_0072_ ), .B1(\u0\/u0\/_0134_ ), .B2(\u0\/u0\/_0078_ ), .Y(\u0\/u0\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1462_ ( .A(\u0\/u0\/_0687_ ), .B(\u0\/u0\/_0236_ ), .C(\u0\/u0\/_0688_ ), .D(\u0\/u0\/_0689_ ), .X(\u0\/u0\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1463_ ( .A(\u0\/u0\/_0680_ ), .B(\u0\/u0\/_0682_ ), .C(\u0\/u0\/_0685_ ), .D(\u0\/u0\/_0690_ ), .X(\u0\/u0\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u0/_1464_ ( .A1(\u0\/u0\/_0532_ ), .A2(\u0\/u0\/_0380_ ), .B1(\u0\/u0\/_0102_ ), .C1(\u0\/u0\/_0355_ ), .X(\u0\/u0\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u0/_1465_ ( .A(\u0\/u0\/_0692_ ), .B(\u0\/u0\/_0338_ ), .C(\u0\/u0\/_0644_ ), .Y(\u0\/u0\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1466_ ( .A(\u0\/u0\/_0016_ ), .B(\u0\/u0\/_0020_ ), .Y(\u0\/u0\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1467_ ( .A1(\u0\/u0\/_0032_ ), .A2(\u0\/u0\/_0137_ ), .B1(\u0\/u0\/_0279_ ), .B2(\u0\/u0\/_0094_ ), .Y(\u0\/u0\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1468_ ( .A1(\u0\/u0\/_0575_ ), .A2(\u0\/u0\/_0153_ ), .B1(\u0\/u0\/_0161_ ), .B2(\u0\/u0\/_0293_ ), .Y(\u0\/u0\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1469_ ( .A(\u0\/u0\/_0259_ ), .B(\u0\/u0\/_0695_ ), .C(\u0\/u0\/_0696_ ), .D(\u0\/u0\/_0697_ ), .X(\u0\/u0\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u0/_1470_ ( .A1(\u0\/u0\/_0255_ ), .A2(\u0\/u0\/_0651_ ), .B1(\u0\/u0\/_0016_ ), .B2(\u0\/u0\/_0193_ ), .X(\u0\/u0\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1471_ ( .A1(\u0\/u0\/_0060_ ), .A2(\u0\/u0\/_0176_ ), .B1(\u0\/u0\/_0699_ ), .C1(\u0\/u0\/_0177_ ), .Y(\u0\/u0\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1472_ ( .A1(\u0\/u0\/_0091_ ), .A2(\u0\/u0\/_0218_ ), .B1(\u0\/u0\/_0092_ ), .B2(\u0\/u0\/_0705_ ), .Y(\u0\/u0\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u0/_1473_ ( .A1(\u0\/u0\/_0705_ ), .A2(\u0\/u0\/_0683_ ), .B1(\u0\/u0\/_0093_ ), .B2(\u0\/u0\/_0114_ ), .Y(\u0\/u0\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u0/_1474_ ( .A1(\u0\/u0\/_0683_ ), .A2(\u0\/u0\/_0084_ ), .B1(\u0\/u0\/_0094_ ), .Y(\u0\/u0\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u0/_1475_ ( .A1(\u0\/u0\/_0543_ ), .A2(\u0\/u0\/_0216_ ), .B1(\u0\/u0\/_0038_ ), .C1(\u0\/u0\/_0056_ ), .Y(\u0\/u0\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1476_ ( .A(\u0\/u0\/_0701_ ), .B(\u0\/u0\/_0702_ ), .C(\u0\/u0\/_0703_ ), .D(\u0\/u0\/_0704_ ), .X(\u0\/u0\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1477_ ( .A(\u0\/u0\/_0693_ ), .B(\u0\/u0\/_0698_ ), .C(\u0\/u0\/_0700_ ), .D(\u0\/u0\/_0706_ ), .X(\u0\/u0\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u0/_1478_ ( .A1(\u0\/u0\/_0113_ ), .A2(\u0\/u0\/_0640_ ), .B1(\u0\/u0\/_0099_ ), .B2(\u0\/u0\/_0058_ ), .X(\u0\/u0\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u0/_1479_ ( .A(\u0\/u0\/_0407_ ), .B(\u0\/u0\/_0708_ ), .C(\u0\/u0\/_0529_ ), .Y(\u0\/u0\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1480_ ( .A(\u0\/u0\/_0568_ ), .B(\u0\/u0\/_0175_ ), .Y(\u0\/u0\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u0/_1481_ ( .A1(\u0\/u0\/_0247_ ), .A2(\u0\/u0\/_0114_ ), .A3(\u0\/u0\/_0051_ ), .B1(\u0\/u0\/_0130_ ), .Y(\u0\/u0\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1482_ ( .A(\u0\/u0\/_0709_ ), .B(\u0\/u0\/_0550_ ), .C(\u0\/u0\/_0710_ ), .D(\u0\/u0\/_0711_ ), .X(\u0\/u0\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u0/_1483_ ( .A1(\u0\/u0\/_0114_ ), .A2(\u0\/u0\/_0064_ ), .B1(\u0\/u0\/_0261_ ), .B2(\u0\/u0\/_0089_ ), .X(\u0\/u0\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1484_ ( .A1(\u0\/u0\/_0355_ ), .A2(\u0\/u0\/_0261_ ), .B1(\u0\/u0\/_0198_ ), .C1(\u0\/u0\/_0713_ ), .Y(\u0\/u0\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1485_ ( .A(\u0\/u0\/_0586_ ), .B(\u0\/u0\/_0478_ ), .Y(\u0\/u0\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u0/_1486_ ( .A_N(\u0\/u0\/_0541_ ), .B(\u0\/u0\/_0267_ ), .C(\u0\/u0\/_0715_ ), .D(\u0\/u0\/_0320_ ), .X(\u0\/u0\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1487_ ( .A(\u0\/u0\/_0586_ ), .B(\u0\/u0\/_0070_ ), .Y(\u0\/u0\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u0/_1488_ ( .A_N(\u0\/u0\/_0211_ ), .B(\u0\/u0\/_0155_ ), .C(\u0\/u0\/_0202_ ), .D(\u0\/u0\/_0718_ ), .X(\u0\/u0\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u0/_1489_ ( .A(\u0\/u0\/_0150_ ), .B(\u0\/u0\/_0216_ ), .C(\u0\/u0\/_0380_ ), .Y(\u0\/u0\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \u0/u0/_1490_ ( .A(\u0\/u0\/_0411_ ), .B(\u0\/u0\/_0720_ ), .X(\u0\/u0\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u0/_1491_ ( .A1(\u0\/u0\/_0018_ ), .A2(\u0\/u0\/_0023_ ), .B1(\u0\/u0\/_0078_ ), .X(\u0\/u0\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u0/_1492_ ( .A1(\u0\/u0\/_0134_ ), .A2(\u0\/u0\/_0738_ ), .B1(\u0\/u0\/_0101_ ), .C1(\u0\/u0\/_0722_ ), .Y(\u0\/u0\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1493_ ( .A(\u0\/u0\/_0717_ ), .B(\u0\/u0\/_0719_ ), .C(\u0\/u0\/_0721_ ), .D(\u0\/u0\/_0723_ ), .X(\u0\/u0\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u0/_1494_ ( .A(\u0\/u0\/_0739_ ), .B(\u0\/u0\/_0193_ ), .Y(\u0\/u0\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1495_ ( .A(\u0\/u0\/_0344_ ), .B(\u0\/u0\/_0184_ ), .C(\u0\/u0\/_0449_ ), .D(\u0\/u0\/_0725_ ), .X(\u0\/u0\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \u0/u0/_1496_ ( .A(\u0\/u0\/_0712_ ), .B(\u0\/u0\/_0714_ ), .C(\u0\/u0\/_0724_ ), .D(\u0\/u0\/_0726_ ), .X(\u0\/u0\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u0/_1497_ ( .A(\u0\/u0\/_0691_ ), .B(\u0\/u0\/_0707_ ), .C(\u0\/u0\/_0728_ ), .Y(\u0\/u0\/_0015_ ) );
sky130_fd_sc_hd__buf_2 \u0/u0/_1502_ ( .A(\w3\[17\] ), .X(\u0\/u0\/_0001_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u1/_0753_ ( .A(\w3\[10\] ), .B_N(\w3\[11\] ), .Y(\u0\/u1\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_0755_ ( .A(\w3\[9\] ), .B(\w3\[8\] ), .X(\u0\/u1\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_0756_ ( .A(\u0\/u1\/_0096_ ), .B(\u0\/u1\/_0118_ ), .X(\u0\/u1\/_0129_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_0757_ ( .A(\w3\[15\] ), .B(\w3\[14\] ), .X(\u0\/u1\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_0758_ ( .A(\w3\[12\] ), .B(\w3\[13\] ), .Y(\u0\/u1\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0759_ ( .A(\u0\/u1\/_0140_ ), .B(\u0\/u1\/_0151_ ), .X(\u0\/u1\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0761_ ( .A(\u0\/u1\/_0129_ ), .B(\u0\/u1\/_0162_ ), .X(\u0\/u1\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0762_ ( .A(\u0\/u1\/_0096_ ), .X(\u0\/u1\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u1/_0763_ ( .A(\w3\[9\] ), .B_N(\w3\[8\] ), .Y(\u0\/u1\/_0205_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0764_ ( .A(\u0\/u1\/_0205_ ), .X(\u0\/u1\/_0216_ ) );
sky130_fd_sc_hd__and3_1 \u0/u1/_0765_ ( .A(\u0\/u1\/_0162_ ), .B(\u0\/u1\/_0194_ ), .C(\u0\/u1\/_0216_ ), .X(\u0\/u1\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \u0/u1/_0766_ ( .A(\u0\/u1\/_0183_ ), .SLEEP(\u0\/u1\/_0227_ ), .X(\u0\/u1\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u1/_0767_ ( .A(\w3\[8\] ), .B_N(\w3\[9\] ), .Y(\u0\/u1\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_0768_ ( .A(\w3\[10\] ), .B(\w3\[11\] ), .Y(\u0\/u1\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0769_ ( .A(\u0\/u1\/_0249_ ), .B(\u0\/u1\/_0260_ ), .X(\u0\/u1\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0771_ ( .A(\u0\/u1\/_0271_ ), .X(\u0\/u1\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0772_ ( .A(\u0\/u1\/_0162_ ), .X(\u0\/u1\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_0773_ ( .A(\u0\/u1\/_0293_ ), .B(\u0\/u1\/_0304_ ), .Y(\u0\/u1\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \u0/u1/_0774_ ( .A(\w3\[9\] ), .Y(\u0\/u1\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \u0/u1/_0776_ ( .A(\w3\[8\] ), .Y(\u0\/u1\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0777_ ( .A(\w3\[10\] ), .B(\w3\[11\] ), .X(\u0\/u1\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0779_ ( .A(\u0\/u1\/_0358_ ), .X(\u0\/u1\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_0780_ ( .A1(\u0\/u1\/_0325_ ), .A2(\u0\/u1\/_0347_ ), .B1(\u0\/u1\/_0380_ ), .C1(\u0\/u1\/_0304_ ), .Y(\u0\/u1\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u1/_0781_ ( .A_N(\u0\/u1\/_0238_ ), .B(\u0\/u1\/_0314_ ), .C(\u0\/u1\/_0391_ ), .X(\u0\/u1\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u1/_0782_ ( .A(\w3\[11\] ), .B_N(\w3\[10\] ), .Y(\u0\/u1\/_0412_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0784_ ( .A(\u0\/u1\/_0412_ ), .B(\u0\/u1\/_0205_ ), .X(\u0\/u1\/_0434_ ) );
sky130_fd_sc_hd__buf_2 \u0/u1/_0786_ ( .A(\u0\/u1\/_0434_ ), .X(\u0\/u1\/_0456_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u1/_0787_ ( .A(\w3\[13\] ), .B_N(\w3\[12\] ), .Y(\u0\/u1\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0788_ ( .A(\u0\/u1\/_0467_ ), .B(\u0\/u1\/_0140_ ), .X(\u0\/u1\/_0478_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_0791_ ( .A(\u0\/u1\/_0456_ ), .B(\u0\/u1\/_0218_ ), .Y(\u0\/u1\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_0792_ ( .A(\u0\/u1\/_0478_ ), .B(\u0\/u1\/_0271_ ), .Y(\u0\/u1\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0793_ ( .A(\u0\/u1\/_0194_ ), .X(\u0\/u1\/_0532_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0794_ ( .A(\u0\/u1\/_0249_ ), .X(\u0\/u1\/_0543_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_0795_ ( .A(\u0\/u1\/_0543_ ), .B(\u0\/u1\/_0358_ ), .X(\u0\/u1\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0797_ ( .A(\u0\/u1\/_0554_ ), .X(\u0\/u1\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_0798_ ( .A(\u0\/u1\/_0216_ ), .B(\u0\/u1\/_0358_ ), .X(\u0\/u1\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0800_ ( .A(\u0\/u1\/_0586_ ), .X(\u0\/u1\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_0801_ ( .A1(\u0\/u1\/_0532_ ), .A2(\u0\/u1\/_0575_ ), .A3(\u0\/u1\/_0608_ ), .B1(\u0\/u1\/_0218_ ), .Y(\u0\/u1\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_0802_ ( .A(\u0\/u1\/_0401_ ), .B(\u0\/u1\/_0510_ ), .C(\u0\/u1\/_0521_ ), .D(\u0\/u1\/_0619_ ), .X(\u0\/u1\/_0629_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_0803_ ( .A(\u0\/u1\/_0358_ ), .B(\w3\[9\] ), .X(\u0\/u1\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0805_ ( .A(\u0\/u1\/_0205_ ), .B(\u0\/u1\/_0260_ ), .X(\u0\/u1\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0807_ ( .A(\u0\/u1\/_0662_ ), .X(\u0\/u1\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u1/_0808_ ( .A(\w3\[14\] ), .B_N(\w3\[15\] ), .Y(\u0\/u1\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_0809_ ( .A(\u0\/u1\/_0467_ ), .B(\u0\/u1\/_0694_ ), .X(\u0\/u1\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0811_ ( .A(\u0\/u1\/_0705_ ), .X(\u0\/u1\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_0812_ ( .A1(\u0\/u1\/_0640_ ), .A2(\u0\/u1\/_0293_ ), .A3(\u0\/u1\/_0683_ ), .B1(\u0\/u1\/_0727_ ), .Y(\u0\/u1\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_0813_ ( .A(\w3\[9\] ), .B(\w3\[8\] ), .Y(\u0\/u1\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0814_ ( .A(\u0\/u1\/_0730_ ), .B(\u0\/u1\/_0260_ ), .X(\u0\/u1\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0816_ ( .A(\u0\/u1\/_0731_ ), .X(\u0\/u1\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0817_ ( .A(\w3\[8\] ), .X(\u0\/u1\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u1/_0818_ ( .A1(\u0\/u1\/_0325_ ), .A2(\u0\/u1\/_0734_ ), .B1(\u0\/u1\/_0412_ ), .X(\u0\/u1\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0819_ ( .A(\u0\/u1\/_0694_ ), .B(\u0\/u1\/_0151_ ), .X(\u0\/u1\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0821_ ( .A(\u0\/u1\/_0736_ ), .X(\u0\/u1\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0822_ ( .A(\u0\/u1\/_0738_ ), .X(\u0\/u1\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_0823_ ( .A1(\u0\/u1\/_0733_ ), .A2(\u0\/u1\/_0735_ ), .A3(\u0\/u1\/_0293_ ), .B1(\u0\/u1\/_0739_ ), .Y(\u0\/u1\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u1/_0824_ ( .A(\u0\/u1\/_0730_ ), .B_N(\u0\/u1\/_0358_ ), .Y(\u0\/u1\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_0825_ ( .A(\u0\/u1\/_0741_ ), .B(\u0\/u1\/_0739_ ), .Y(\u0\/u1\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_0827_ ( .A1(\u0\/u1\/_0118_ ), .A2(\u0\/u1\/_0216_ ), .B1(\u0\/u1\/_0532_ ), .C1(\u0\/u1\/_0739_ ), .Y(\u0\/u1\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_0828_ ( .A(\u0\/u1\/_0729_ ), .B(\u0\/u1\/_0740_ ), .C(\u0\/u1\/_0742_ ), .D(\u0\/u1\/_0744_ ), .X(\u0\/u1\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0829_ ( .A(\u0\/u1\/_0412_ ), .B(\u0\/u1\/_0730_ ), .X(\u0\/u1\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0831_ ( .A(\u0\/u1\/_0746_ ), .X(\u0\/u1\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u1/_0832_ ( .A(\w3\[12\] ), .B_N(\w3\[13\] ), .Y(\u0\/u1\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0833_ ( .A(\u0\/u1\/_0749_ ), .B(\u0\/u1\/_0694_ ), .X(\u0\/u1\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0835_ ( .A(\u0\/u1\/_0750_ ), .X(\u0\/u1\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0836_ ( .A(\u0\/u1\/_0752_ ), .X(\u0\/u1\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0837_ ( .A(\u0\/u1\/_0118_ ), .B(\u0\/u1\/_0358_ ), .X(\u0\/u1\/_0017_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0839_ ( .A(\u0\/u1\/_0752_ ), .B(\u0\/u1\/_0017_ ), .X(\u0\/u1\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0840_ ( .A(\u0\/u1\/_0358_ ), .B(\u0\/u1\/_0325_ ), .X(\u0\/u1\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0842_ ( .A(\u0\/u1\/_0096_ ), .B(\u0\/u1\/_0205_ ), .X(\u0\/u1\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u1/_0844_ ( .A1(\u0\/u1\/_0020_ ), .A2(\u0\/u1\/_0022_ ), .B1(\u0\/u1\/_0752_ ), .X(\u0\/u1\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_0845_ ( .A1(\u0\/u1\/_0748_ ), .A2(\u0\/u1\/_0016_ ), .B1(\u0\/u1\/_0019_ ), .C1(\u0\/u1\/_0024_ ), .Y(\u0\/u1\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_0846_ ( .A(\w3\[12\] ), .B(\w3\[13\] ), .X(\u0\/u1\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0847_ ( .A(\u0\/u1\/_0694_ ), .B(\u0\/u1\/_0026_ ), .X(\u0\/u1\/_0027_ ) );
sky130_fd_sc_hd__buf_2 \u0/u1/_0849_ ( .A(\u0\/u1\/_0027_ ), .X(\u0\/u1\/_0029_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0850_ ( .A(\u0\/u1\/_0358_ ), .B(\u0\/u1\/_0730_ ), .X(\u0\/u1\/_0030_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0852_ ( .A(\u0\/u1\/_0030_ ), .X(\u0\/u1\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_0853_ ( .A(\u0\/u1\/_0029_ ), .B(\u0\/u1\/_0032_ ), .Y(\u0\/u1\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_0854_ ( .A(\u0\/u1\/_0029_ ), .B(\u0\/u1\/_0735_ ), .Y(\u0\/u1\/_0034_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0855_ ( .A(\u0\/u1\/_0118_ ), .B(\u0\/u1\/_0260_ ), .X(\u0\/u1\/_0035_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0857_ ( .A(\u0\/u1\/_0027_ ), .B(\u0\/u1\/_0035_ ), .X(\u0\/u1\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0858_ ( .A(\u0\/u1\/_0260_ ), .X(\u0\/u1\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_0859_ ( .A(\u0\/u1\/_0038_ ), .B(\u0\/u1\/_0347_ ), .Y(\u0\/u1\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u1/_0860_ ( .A_N(\u0\/u1\/_0039_ ), .B(\u0\/u1\/_0027_ ), .X(\u0\/u1\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_0861_ ( .A(\u0\/u1\/_0037_ ), .B(\u0\/u1\/_0040_ ), .Y(\u0\/u1\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_0862_ ( .A(\u0\/u1\/_0025_ ), .B(\u0\/u1\/_0033_ ), .C(\u0\/u1\/_0034_ ), .D(\u0\/u1\/_0041_ ), .X(\u0\/u1\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0863_ ( .A(\u0\/u1\/_0749_ ), .B(\u0\/u1\/_0140_ ), .X(\u0\/u1\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \u0/u1/_0865_ ( .A(\w3\[8\] ), .B(\w3\[10\] ), .C(\w3\[11\] ), .X(\u0\/u1\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0866_ ( .A(\u0\/u1\/_0043_ ), .B(\u0\/u1\/_0045_ ), .X(\u0\/u1\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0867_ ( .A(\u0\/u1\/_0096_ ), .B(\u0\/u1\/_0543_ ), .X(\u0\/u1\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0869_ ( .A(\u0\/u1\/_0047_ ), .B(\u0\/u1\/_0043_ ), .X(\u0\/u1\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0870_ ( .A(\u0\/u1\/_0730_ ), .X(\u0\/u1\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0871_ ( .A(\u0\/u1\/_0043_ ), .X(\u0\/u1\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_0872_ ( .A1(\u0\/u1\/_0118_ ), .A2(\u0\/u1\/_0050_ ), .B1(\u0\/u1\/_0194_ ), .C1(\u0\/u1\/_0051_ ), .Y(\u0\/u1\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u1/_0873_ ( .A(\u0\/u1\/_0046_ ), .B(\u0\/u1\/_0049_ ), .C_N(\u0\/u1\/_0052_ ), .Y(\u0\/u1\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0874_ ( .A(\u0\/u1\/_0026_ ), .B(\u0\/u1\/_0140_ ), .X(\u0\/u1\/_0054_ ) );
sky130_fd_sc_hd__buf_2 \u0/u1/_0876_ ( .A(\u0\/u1\/_0054_ ), .X(\u0\/u1\/_0056_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_0877_ ( .A1(\u0\/u1\/_0532_ ), .A2(\u0\/u1\/_0575_ ), .B1(\u0\/u1\/_0056_ ), .Y(\u0\/u1\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0878_ ( .A(\u0\/u1\/_0412_ ), .B(\u0\/u1\/_0325_ ), .X(\u0\/u1\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0880_ ( .A(\u0\/u1\/_0051_ ), .X(\u0\/u1\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_0881_ ( .A1(\u0\/u1\/_0731_ ), .A2(\u0\/u1\/_0035_ ), .A3(\u0\/u1\/_0058_ ), .B1(\u0\/u1\/_0060_ ), .Y(\u0\/u1\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0882_ ( .A(\u0\/u1\/_0260_ ), .B(\w3\[9\] ), .X(\u0\/u1\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0884_ ( .A(\u0\/u1\/_0062_ ), .X(\u0\/u1\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_0885_ ( .A1(\u0\/u1\/_0064_ ), .A2(\u0\/u1\/_0748_ ), .A3(\u0\/u1\/_0683_ ), .B1(\u0\/u1\/_0056_ ), .Y(\u0\/u1\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_0886_ ( .A(\u0\/u1\/_0053_ ), .B(\u0\/u1\/_0057_ ), .C(\u0\/u1\/_0061_ ), .D(\u0\/u1\/_0065_ ), .X(\u0\/u1\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_0887_ ( .A(\u0\/u1\/_0629_ ), .B(\u0\/u1\/_0745_ ), .C(\u0\/u1\/_0042_ ), .D(\u0\/u1\/_0066_ ), .X(\u0\/u1\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u1/_0889_ ( .A(\w3\[15\] ), .B_N(\w3\[14\] ), .Y(\u0\/u1\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0890_ ( .A(\u0\/u1\/_0069_ ), .B(\u0\/u1\/_0151_ ), .X(\u0\/u1\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0892_ ( .A(\u0\/u1\/_0070_ ), .X(\u0\/u1\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_0893_ ( .A1(\u0\/u1\/_0129_ ), .A2(\u0\/u1\/_0586_ ), .B1(\u0\/u1\/_0072_ ), .Y(\u0\/u1\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_0894_ ( .A1(\u0\/u1\/_0380_ ), .A2(\u0\/u1\/_0347_ ), .B1(\u0\/u1\/_0194_ ), .B2(\u0\/u1\/_0216_ ), .Y(\u0\/u1\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u1/_0895_ ( .A(\u0\/u1\/_0074_ ), .B_N(\u0\/u1\/_0070_ ), .Y(\u0\/u1\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u1/_0896_ ( .A(\u0\/u1\/_0073_ ), .SLEEP(\u0\/u1\/_0075_ ), .X(\u0\/u1\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_0897_ ( .A(\u0\/u1\/_0467_ ), .B(\u0\/u1\/_0069_ ), .X(\u0\/u1\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0898_ ( .A(\u0\/u1\/_0077_ ), .X(\u0\/u1\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0899_ ( .A(\u0\/u1\/_0412_ ), .B(\u0\/u1\/_0118_ ), .X(\u0\/u1\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0901_ ( .A(\u0\/u1\/_0078_ ), .B(\u0\/u1\/_0079_ ), .X(\u0\/u1\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0902_ ( .A(\u0\/u1\/_0412_ ), .B(\u0\/u1\/_0249_ ), .X(\u0\/u1\/_0082_ ) );
sky130_fd_sc_hd__buf_2 \u0/u1/_0904_ ( .A(\u0\/u1\/_0082_ ), .X(\u0\/u1\/_0084_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0905_ ( .A(\u0\/u1\/_0084_ ), .B(\u0\/u1\/_0078_ ), .X(\u0\/u1\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u1/_0906_ ( .A1(\w3\[8\] ), .A2(\u0\/u1\/_0325_ ), .B1(\u0\/u1\/_0260_ ), .Y(\u0\/u1\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u1/_0907_ ( .A_N(\u0\/u1\/_0086_ ), .B(\u0\/u1\/_0078_ ), .X(\u0\/u1\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u1/_0908_ ( .A(\u0\/u1\/_0081_ ), .B(\u0\/u1\/_0085_ ), .C(\u0\/u1\/_0087_ ), .Y(\u0\/u1\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0909_ ( .A(\u0\/u1\/_0072_ ), .X(\u0\/u1\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_0910_ ( .A1(\u0\/u1\/_0733_ ), .A2(\u0\/u1\/_0748_ ), .A3(\u0\/u1\/_0683_ ), .B1(\u0\/u1\/_0089_ ), .Y(\u0\/u1\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0911_ ( .A(\u0\/u1\/_0129_ ), .X(\u0\/u1\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0912_ ( .A(\u0\/u1\/_0017_ ), .X(\u0\/u1\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0913_ ( .A(\u0\/u1\/_0022_ ), .X(\u0\/u1\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0914_ ( .A(\u0\/u1\/_0078_ ), .X(\u0\/u1\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_0915_ ( .A1(\u0\/u1\/_0091_ ), .A2(\u0\/u1\/_0092_ ), .A3(\u0\/u1\/_0093_ ), .B1(\u0\/u1\/_0094_ ), .Y(\u0\/u1\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_0916_ ( .A(\u0\/u1\/_0076_ ), .B(\u0\/u1\/_0088_ ), .C(\u0\/u1\/_0090_ ), .D(\u0\/u1\/_0095_ ), .X(\u0\/u1\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_0917_ ( .A(\u0\/u1\/_0069_ ), .B(\u0\/u1\/_0026_ ), .X(\u0\/u1\/_0098_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0918_ ( .A(\u0\/u1\/_0098_ ), .X(\u0\/u1\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0919_ ( .A(\u0\/u1\/_0434_ ), .B(\u0\/u1\/_0099_ ), .X(\u0\/u1\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0920_ ( .A(\u0\/u1\/_0079_ ), .B(\u0\/u1\/_0098_ ), .X(\u0\/u1\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0921_ ( .A(\u0\/u1\/_0325_ ), .X(\u0\/u1\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_0922_ ( .A1(\u0\/u1\/_0102_ ), .A2(\u0\/u1\/_0734_ ), .B1(\u0\/u1\/_0038_ ), .C1(\u0\/u1\/_0099_ ), .Y(\u0\/u1\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u1/_0923_ ( .A(\u0\/u1\/_0100_ ), .B(\u0\/u1\/_0101_ ), .C_N(\u0\/u1\/_0103_ ), .Y(\u0\/u1\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_0924_ ( .A1(\u0\/u1\/_0554_ ), .A2(\u0\/u1\/_0586_ ), .B1(\u0\/u1\/_0099_ ), .Y(\u0\/u1\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_0925_ ( .A(\u0\/u1\/_0129_ ), .B(\u0\/u1\/_0099_ ), .Y(\u0\/u1\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0926_ ( .A(\u0\/u1\/_0105_ ), .B(\u0\/u1\/_0106_ ), .X(\u0\/u1\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0927_ ( .A(\u0\/u1\/_0412_ ), .X(\u0\/u1\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_0928_ ( .A(\u0\/u1\/_0260_ ), .B(\w3\[8\] ), .X(\u0\/u1\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0929_ ( .A(\u0\/u1\/_0069_ ), .B(\u0\/u1\/_0749_ ), .X(\u0\/u1\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0931_ ( .A(\u0\/u1\/_0111_ ), .X(\u0\/u1\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0932_ ( .A(\u0\/u1\/_0113_ ), .X(\u0\/u1\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_0933_ ( .A1(\u0\/u1\/_0109_ ), .A2(\u0\/u1\/_0110_ ), .B1(\u0\/u1\/_0114_ ), .Y(\u0\/u1\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_0934_ ( .A(\u0\/u1\/_0022_ ), .Y(\u0\/u1\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_0935_ ( .A(\u0\/u1\/_0554_ ), .Y(\u0\/u1\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u1/_0936_ ( .A1(\u0\/u1\/_0050_ ), .A2(\u0\/u1\/_0118_ ), .B1(\u0\/u1\/_0194_ ), .Y(\u0\/u1\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_0937_ ( .A(\u0\/u1\/_0113_ ), .Y(\u0\/u1\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \u0/u1/_0938_ ( .A1(\u0\/u1\/_0116_ ), .A2(\u0\/u1\/_0117_ ), .A3(\u0\/u1\/_0119_ ), .B1(\u0\/u1\/_0120_ ), .X(\u0\/u1\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_0939_ ( .A(\u0\/u1\/_0104_ ), .B(\u0\/u1\/_0108_ ), .C(\u0\/u1\/_0115_ ), .D(\u0\/u1\/_0121_ ), .X(\u0\/u1\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_0940_ ( .A(\w3\[15\] ), .B(\w3\[14\] ), .Y(\u0\/u1\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0941_ ( .A(\u0\/u1\/_0749_ ), .B(\u0\/u1\/_0123_ ), .X(\u0\/u1\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0943_ ( .A(\u0\/u1\/_0082_ ), .B(\u0\/u1\/_0124_ ), .X(\u0\/u1\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_0944_ ( .A(\u0\/u1\/_0271_ ), .B(\u0\/u1\/_0124_ ), .Y(\u0\/u1\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0945_ ( .A(\u0\/u1\/_0124_ ), .X(\u0\/u1\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0946_ ( .A(\u0\/u1\/_0260_ ), .B(\u0\/u1\/_0325_ ), .X(\u0\/u1\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_0948_ ( .A(\u0\/u1\/_0128_ ), .B(\u0\/u1\/_0130_ ), .Y(\u0\/u1\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_0949_ ( .A(\u0\/u1\/_0127_ ), .B(\u0\/u1\/_0132_ ), .Y(\u0\/u1\/_0133_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_0951_ ( .A(\u0\/u1\/_0456_ ), .B(\u0\/u1\/_0128_ ), .Y(\u0\/u1\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u1/_0952_ ( .A(\u0\/u1\/_0126_ ), .B(\u0\/u1\/_0133_ ), .C_N(\u0\/u1\/_0135_ ), .Y(\u0\/u1\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_0953_ ( .A(\u0\/u1\/_0026_ ), .B(\u0\/u1\/_0123_ ), .X(\u0\/u1\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0955_ ( .A(\u0\/u1\/_0137_ ), .X(\u0\/u1\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_0956_ ( .A1(\u0\/u1\/_0110_ ), .A2(\u0\/u1\/_0293_ ), .A3(\u0\/u1\/_0084_ ), .B1(\u0\/u1\/_0139_ ), .Y(\u0\/u1\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0957_ ( .A(\u0\/u1\/_0096_ ), .B(\u0\/u1\/_0730_ ), .X(\u0\/u1\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0959_ ( .A(\u0\/u1\/_0142_ ), .X(\u0\/u1\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_0960_ ( .A1(\u0\/u1\/_0020_ ), .A2(\u0\/u1\/_0144_ ), .A3(\u0\/u1\/_0017_ ), .B1(\u0\/u1\/_0139_ ), .Y(\u0\/u1\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u1/_0961_ ( .A(\w3\[10\] ), .B(\u0\/u1\/_0050_ ), .C_N(\w3\[11\] ), .Y(\u0\/u1\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0962_ ( .A(\u0\/u1\/_0128_ ), .X(\u0\/u1\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_0963_ ( .A1(\u0\/u1\/_0146_ ), .A2(\u0\/u1\/_0032_ ), .A3(\u0\/u1\/_0640_ ), .B1(\u0\/u1\/_0147_ ), .Y(\u0\/u1\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_0964_ ( .A(\u0\/u1\/_0136_ ), .B(\u0\/u1\/_0141_ ), .C(\u0\/u1\/_0145_ ), .D(\u0\/u1\/_0148_ ), .X(\u0\/u1\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0965_ ( .A(\u0\/u1\/_0123_ ), .B(\u0\/u1\/_0151_ ), .X(\u0\/u1\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0967_ ( .A(\u0\/u1\/_0150_ ), .X(\u0\/u1\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_0968_ ( .A(\u0\/u1\/_0150_ ), .B(\u0\/u1\/_0062_ ), .X(\u0\/u1\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_0969_ ( .A(\u0\/u1\/_0079_ ), .B(\u0\/u1\/_0150_ ), .Y(\u0\/u1\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u1/_0970_ ( .A(\u0\/u1\/_0150_ ), .B(\u0\/u1\/_0412_ ), .C(\u0\/u1\/_0543_ ), .Y(\u0\/u1\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_0971_ ( .A(\u0\/u1\/_0155_ ), .B(\u0\/u1\/_0156_ ), .Y(\u0\/u1\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_0972_ ( .A1(\u0\/u1\/_0153_ ), .A2(\u0\/u1\/_0456_ ), .B1(\u0\/u1\/_0154_ ), .C1(\u0\/u1\/_0157_ ), .Y(\u0\/u1\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0973_ ( .A(\u0\/u1\/_0467_ ), .B(\u0\/u1\/_0123_ ), .X(\u0\/u1\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_0975_ ( .A(\u0\/u1\/_0159_ ), .X(\u0\/u1\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u1/_0976_ ( .A_N(\u0\/u1\/_0119_ ), .B(\u0\/u1\/_0161_ ), .X(\u0\/u1\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_0977_ ( .A(\u0\/u1\/_0163_ ), .Y(\u0\/u1\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_0978_ ( .A1(\u0\/u1\/_0146_ ), .A2(\u0\/u1\/_0575_ ), .A3(\u0\/u1\/_0608_ ), .B1(\u0\/u1\/_0153_ ), .Y(\u0\/u1\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_0979_ ( .A1(\u0\/u1\/_0062_ ), .A2(\u0\/u1\/_0084_ ), .A3(\u0\/u1\/_0456_ ), .B1(\u0\/u1\/_0161_ ), .Y(\u0\/u1\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_0980_ ( .A(\u0\/u1\/_0158_ ), .B(\u0\/u1\/_0164_ ), .C(\u0\/u1\/_0165_ ), .D(\u0\/u1\/_0166_ ), .X(\u0\/u1\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_0981_ ( .A(\u0\/u1\/_0097_ ), .B(\u0\/u1\/_0122_ ), .C(\u0\/u1\/_0149_ ), .D(\u0\/u1\/_0167_ ), .X(\u0\/u1\/_0168_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0982_ ( .A(\u0\/u1\/_0662_ ), .B(\u0\/u1\/_0150_ ), .X(\u0\/u1\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_0983_ ( .A(\u0\/u1\/_0154_ ), .B(\u0\/u1\/_0169_ ), .Y(\u0\/u1\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \u0/u1/_0984_ ( .A(\u0\/u1\/_0123_ ), .B(\u0\/u1\/_0151_ ), .C(\u0\/u1\/_0038_ ), .X(\u0\/u1\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0985_ ( .A(\u0\/u1\/_0170_ ), .B(\u0\/u1\/_0171_ ), .X(\u0\/u1\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_0986_ ( .A(\u0\/u1\/_0172_ ), .Y(\u0\/u1\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u1/_0987_ ( .A(\u0\/u1\/_0067_ ), .B(\u0\/u1\/_0168_ ), .C(\u0\/u1\/_0174_ ), .Y(\u0\/u1\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/u1/_0988_ ( .A(\w3\[9\] ), .B(\w3\[8\] ), .Y(\u0\/u1\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_0989_ ( .A(\u0\/u1\/_0175_ ), .B(\u0\/u1\/_0358_ ), .X(\u0\/u1\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0990_ ( .A(\u0\/u1\/_0176_ ), .B(\u0\/u1\/_0478_ ), .X(\u0\/u1\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_0991_ ( .A(\u0\/u1\/_0084_ ), .B(\u0\/u1\/_0113_ ), .Y(\u0\/u1\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0992_ ( .A(\u0\/u1\/_0111_ ), .B(\u0\/u1\/_0062_ ), .X(\u0\/u1\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0993_ ( .A(\u0\/u1\/_0111_ ), .B(\u0\/u1\/_0662_ ), .X(\u0\/u1\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_0994_ ( .A(\u0\/u1\/_0179_ ), .B(\u0\/u1\/_0180_ ), .Y(\u0\/u1\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0995_ ( .A(\u0\/u1\/_0054_ ), .B(\u0\/u1\/_0058_ ), .X(\u0\/u1\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_0996_ ( .A(\u0\/u1\/_0182_ ), .Y(\u0\/u1\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u1/_0997_ ( .A_N(\u0\/u1\/_0177_ ), .B(\u0\/u1\/_0178_ ), .C(\u0\/u1\/_0181_ ), .D(\u0\/u1\/_0184_ ), .X(\u0\/u1\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0998_ ( .A(\u0\/u1\/_0098_ ), .B(\u0\/u1\/_0741_ ), .X(\u0\/u1\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_0999_ ( .A(\u0\/u1\/_0047_ ), .B(\u0\/u1\/_0098_ ), .X(\u0\/u1\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \u0/u1/_1000_ ( .A(\u0\/u1\/_0186_ ), .B(\u0\/u1\/_0187_ ), .X(\u0\/u1\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1001_ ( .A(\u0\/u1\/_0188_ ), .Y(\u0\/u1\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1002_ ( .A(\u0\/u1\/_0738_ ), .B(\u0\/u1\/_0735_ ), .X(\u0\/u1\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1003_ ( .A(\u0\/u1\/_0271_ ), .B(\u0\/u1\/_0736_ ), .X(\u0\/u1\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_1004_ ( .A(\u0\/u1\/_0190_ ), .B(\u0\/u1\/_0191_ ), .Y(\u0\/u1\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_1005_ ( .A(\u0\/u1\/_0096_ ), .B(\u0\/u1\/_0325_ ), .X(\u0\/u1\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1006_ ( .A1(\u0\/u1\/_0193_ ), .A2(\u0\/u1\/_0176_ ), .B1(\u0\/u1\/_0043_ ), .Y(\u0\/u1\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1007_ ( .A(\u0\/u1\/_0185_ ), .B(\u0\/u1\/_0189_ ), .C(\u0\/u1\/_0192_ ), .D(\u0\/u1\/_0195_ ), .X(\u0\/u1\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u1/_1008_ ( .A_N(\w3\[11\] ), .B(\u0\/u1\/_0734_ ), .C(\w3\[10\] ), .X(\u0\/u1\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1009_ ( .A(\u0\/u1\/_0137_ ), .B(\u0\/u1\/_0197_ ), .X(\u0\/u1\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_1010_ ( .A(\u0\/u1\/_0198_ ), .B(\u0\/u1\/_0040_ ), .Y(\u0\/u1\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1011_ ( .A(\u0\/u1\/_0293_ ), .B(\u0\/u1\/_0137_ ), .X(\u0\/u1\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1012_ ( .A(\u0\/u1\/_0200_ ), .Y(\u0\/u1\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1013_ ( .A(\u0\/u1\/_0137_ ), .B(\u0\/u1\/_0110_ ), .Y(\u0\/u1\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1014_ ( .A(\u0\/u1\/_0139_ ), .B(\u0\/u1\/_0020_ ), .Y(\u0\/u1\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1015_ ( .A(\u0\/u1\/_0199_ ), .B(\u0\/u1\/_0201_ ), .C(\u0\/u1\/_0202_ ), .D(\u0\/u1\/_0203_ ), .X(\u0\/u1\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u1/_1016_ ( .A1(\u0\/u1\/_0532_ ), .A2(\u0\/u1\/_0109_ ), .B1(\u0\/u1\/_0102_ ), .C1(\u0\/u1\/_0727_ ), .X(\u0\/u1\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1017_ ( .A(\u0\/u1\/_0022_ ), .B(\u0\/u1\/_0078_ ), .Y(\u0\/u1\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1018_ ( .A(\u0\/u1\/_0078_ ), .B(\u0\/u1\/_0142_ ), .Y(\u0\/u1\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1019_ ( .A(\u0\/u1\/_0207_ ), .B(\u0\/u1\/_0208_ ), .Y(\u0\/u1\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1020_ ( .A1(\u0\/u1\/_0094_ ), .A2(\u0\/u1\/_0176_ ), .B1(\u0\/u1\/_0206_ ), .C1(\u0\/u1\/_0209_ ), .Y(\u0\/u1\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1021_ ( .A(\u0\/u1\/_0662_ ), .B(\u0\/u1\/_0070_ ), .X(\u0\/u1\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u1/_1022_ ( .A(\u0\/u1\/_0731_ ), .B(\u0\/u1\/_0123_ ), .C(\u0\/u1\/_0749_ ), .Y(\u0\/u1\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u1/_1023_ ( .A(\u0\/u1\/_0731_ ), .B(\u0\/u1\/_0467_ ), .C(\u0\/u1\/_0069_ ), .Y(\u0\/u1\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u1/_1024_ ( .A_N(\u0\/u1\/_0211_ ), .B(\u0\/u1\/_0127_ ), .C(\u0\/u1\/_0212_ ), .D(\u0\/u1\/_0213_ ), .X(\u0\/u1\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1025_ ( .A(\u0\/u1\/_0137_ ), .Y(\u0\/u1\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1026_ ( .A(\u0\/u1\/_0128_ ), .B(\u0\/u1\/_0035_ ), .Y(\u0\/u1\/_0217_ ) );
sky130_fd_sc_hd__buf_2 \u0/u1/_1027_ ( .A(\u0\/u1\/_0478_ ), .X(\u0\/u1\/_0218_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1028_ ( .A1(\u0\/u1\/_0159_ ), .A2(\u0\/u1\/_0746_ ), .B1(\u0\/u1\/_0434_ ), .B2(\u0\/u1\/_0218_ ), .Y(\u0\/u1\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u1/_1029_ ( .A1(\u0\/u1\/_0116_ ), .A2(\u0\/u1\/_0215_ ), .B1(\u0\/u1\/_0217_ ), .C1(\u0\/u1\/_0219_ ), .X(\u0\/u1\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1030_ ( .A(\u0\/u1\/_0113_ ), .B(\u0\/u1\/_0746_ ), .X(\u0\/u1\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u1/_1031_ ( .A1(\u0\/u1\/_0098_ ), .A2(\u0\/u1\/_0746_ ), .B1(\u0\/u1\/_0434_ ), .B2(\u0\/u1\/_0750_ ), .X(\u0\/u1\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1032_ ( .A1(\u0\/u1\/_0047_ ), .A2(\u0\/u1\/_0113_ ), .B1(\u0\/u1\/_0221_ ), .C1(\u0\/u1\/_0222_ ), .Y(\u0\/u1\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u1/_1033_ ( .A1(\u0\/u1\/_0129_ ), .A2(\u0\/u1\/_0162_ ), .B1(\u0\/u1\/_0271_ ), .B2(\u0\/u1\/_0705_ ), .X(\u0\/u1\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1034_ ( .A1(\u0\/u1\/_0093_ ), .A2(\u0\/u1\/_0738_ ), .B1(\u0\/u1\/_0081_ ), .C1(\u0\/u1\/_0224_ ), .Y(\u0\/u1\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1035_ ( .A(\u0\/u1\/_0214_ ), .B(\u0\/u1\/_0220_ ), .C(\u0\/u1\/_0223_ ), .D(\u0\/u1\/_0225_ ), .X(\u0\/u1\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1036_ ( .A(\u0\/u1\/_0196_ ), .B(\u0\/u1\/_0204_ ), .C(\u0\/u1\/_0210_ ), .D(\u0\/u1\/_0226_ ), .X(\u0\/u1\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1037_ ( .A(\u0\/u1\/_0111_ ), .B(\u0\/u1\/_0554_ ), .X(\u0\/u1\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1038_ ( .A(\u0\/u1\/_0229_ ), .Y(\u0\/u1\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1039_ ( .A(\u0\/u1\/_0111_ ), .B(\u0\/u1\/_0129_ ), .Y(\u0\/u1\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1040_ ( .A(\u0\/u1\/_0017_ ), .B(\u0\/u1\/_0738_ ), .Y(\u0\/u1\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1041_ ( .A(\u0\/u1\/_0030_ ), .B(\u0\/u1\/_0304_ ), .Y(\u0\/u1\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1042_ ( .A(\u0\/u1\/_0230_ ), .B(\u0\/u1\/_0231_ ), .C(\u0\/u1\/_0232_ ), .D(\u0\/u1\/_0233_ ), .X(\u0\/u1\/_0234_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1043_ ( .A(\u0\/u1\/_0047_ ), .B(\u0\/u1\/_0478_ ), .X(\u0\/u1\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1044_ ( .A1(\u0\/u1\/_0129_ ), .A2(\u0\/u1\/_0554_ ), .B1(\u0\/u1\/_0137_ ), .Y(\u0\/u1\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u1/_1045_ ( .A(\u0\/u1\/_0235_ ), .B(\u0\/u1\/_0049_ ), .C_N(\u0\/u1\/_0236_ ), .Y(\u0\/u1\/_0237_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_1046_ ( .A(\u0\/u1\/_0047_ ), .B(\u0\/u1\/_0077_ ), .X(\u0\/u1\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1047_ ( .A(\u0\/u1\/_0070_ ), .B(\u0\/u1\/_0035_ ), .X(\u0\/u1\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u1/_1048_ ( .A1(\u0\/u1\/_0047_ ), .A2(\u0\/u1\/_0736_ ), .B1(\u0\/u1\/_0022_ ), .B2(\u0\/u1\/_0099_ ), .X(\u0\/u1\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u1/_1049_ ( .A(\u0\/u1\/_0239_ ), .B(\u0\/u1\/_0240_ ), .C(\u0\/u1\/_0241_ ), .Y(\u0\/u1\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1050_ ( .A(\u0\/u1\/_0554_ ), .B(\u0\/u1\/_0072_ ), .X(\u0\/u1\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u1/_1051_ ( .A1(\u0\/u1\/_0142_ ), .A2(\u0\/u1\/_0137_ ), .B1(\u0\/u1\/_0159_ ), .B2(\u0\/u1\/_0082_ ), .X(\u0\/u1\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1052_ ( .A1(\u0\/u1\/_0608_ ), .A2(\u0\/u1\/_0072_ ), .B1(\u0\/u1\/_0243_ ), .C1(\u0\/u1\/_0244_ ), .Y(\u0\/u1\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1053_ ( .A(\u0\/u1\/_0234_ ), .B(\u0\/u1\/_0237_ ), .C(\u0\/u1\/_0242_ ), .D(\u0\/u1\/_0245_ ), .X(\u0\/u1\/_0246_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u1/_1055_ ( .A1(\u0\/u1\/_0554_ ), .A2(\u0\/u1\/_0586_ ), .B1(\u0\/u1\/_0029_ ), .X(\u0\/u1\/_0248_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1056_ ( .A(\u0\/u1\/_0082_ ), .B(\u0\/u1\/_0478_ ), .X(\u0\/u1\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_1057_ ( .A(\u0\/u1\/_0079_ ), .X(\u0\/u1\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1058_ ( .A(\u0\/u1\/_0251_ ), .B(\u0\/u1\/_0478_ ), .X(\u0\/u1\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_1059_ ( .A(\u0\/u1\/_0250_ ), .B(\u0\/u1\/_0252_ ), .Y(\u0\/u1\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1060_ ( .A(\u0\/u1\/_0016_ ), .B(\u0\/u1\/_0064_ ), .Y(\u0\/u1\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_1061_ ( .A(\u0\/u1\/_0304_ ), .X(\u0\/u1\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1062_ ( .A(\u0\/u1\/_0255_ ), .B(\u0\/u1\/_0640_ ), .Y(\u0\/u1\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u1/_1063_ ( .A_N(\u0\/u1\/_0248_ ), .B(\u0\/u1\/_0253_ ), .C(\u0\/u1\/_0254_ ), .D(\u0\/u1\/_0256_ ), .X(\u0\/u1\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1064_ ( .A(\u0\/u1\/_0099_ ), .B(\u0\/u1\/_0110_ ), .X(\u0\/u1\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \u0/u1/_1065_ ( .A1(\u0\/u1\/_0161_ ), .A2(\u0\/u1\/_0130_ ), .B1(\u0\/u1\/_0258_ ), .Y(\u0\/u1\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1066_ ( .A(\u0\/u1\/_0194_ ), .B(\w3\[9\] ), .X(\u0\/u1\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1068_ ( .A(\u0\/u1\/_0261_ ), .B(\u0\/u1\/_0153_ ), .Y(\u0\/u1\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u1/_1069_ ( .A_N(\u0\/u1\/_0154_ ), .B(\u0\/u1\/_0259_ ), .C(\u0\/u1\/_0263_ ), .X(\u0\/u1\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1070_ ( .A(\u0\/u1\/_0246_ ), .B(\u0\/u1\/_0174_ ), .C(\u0\/u1\/_0257_ ), .D(\u0\/u1\/_0264_ ), .X(\u0\/u1\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u1/_1071_ ( .A1(\u0\/u1\/_0261_ ), .A2(\u0\/u1\/_0554_ ), .B1(\u0\/u1\/_0159_ ), .X(\u0\/u1\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1072_ ( .A(\u0\/u1\/_0746_ ), .B(\u0\/u1\/_0150_ ), .Y(\u0\/u1\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1073_ ( .A(\u0\/u1\/_0175_ ), .Y(\u0\/u1\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \u0/u1/_1074_ ( .A(\u0\/u1\/_0412_ ), .B(\u0\/u1\/_0123_ ), .C(\u0\/u1\/_0151_ ), .X(\u0\/u1\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1075_ ( .A(\u0\/u1\/_0268_ ), .B(\u0\/u1\/_0269_ ), .Y(\u0\/u1\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u1/_1076_ ( .A_N(\u0\/u1\/_0266_ ), .B(\u0\/u1\/_0267_ ), .C(\u0\/u1\/_0270_ ), .X(\u0\/u1\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1077_ ( .A(\u0\/u1\/_0554_ ), .B(\u0\/u1\/_0150_ ), .X(\u0\/u1\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1078_ ( .A(\u0\/u1\/_0273_ ), .Y(\u0\/u1\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1079_ ( .A1(\u0\/u1\/_0734_ ), .A2(\u0\/u1\/_0325_ ), .B1(\u0\/u1\/_0380_ ), .Y(\u0\/u1\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1080_ ( .A(\u0\/u1\/_0275_ ), .Y(\u0\/u1\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1081_ ( .A(\u0\/u1\/_0276_ ), .B(\u0\/u1\/_0153_ ), .Y(\u0\/u1\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \u0/u1/_1082_ ( .A(\u0\/u1\/_0272_ ), .B(\u0\/u1\/_0274_ ), .C(\u0\/u1\/_0277_ ), .X(\u0\/u1\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_1083_ ( .A(\u0\/u1\/_0035_ ), .X(\u0\/u1\/_0279_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1085_ ( .A1(\u0\/u1\/_0218_ ), .A2(\u0\/u1\/_0279_ ), .B1(\u0\/u1\/_0084_ ), .B2(\u0\/u1\/_0060_ ), .Y(\u0\/u1\/_0281_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u1/_1086_ ( .A1(\u0\/u1\/_0251_ ), .A2(\u0\/u1\/_0434_ ), .B1(\u0\/u1\/_0304_ ), .Y(\u0\/u1\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1087_ ( .A(\u0\/u1\/_0091_ ), .B(\u0\/u1\/_0056_ ), .Y(\u0\/u1\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1088_ ( .A1(\u0\/u1\/_0118_ ), .A2(\u0\/u1\/_0050_ ), .B1(\u0\/u1\/_0038_ ), .C1(\u0\/u1\/_0255_ ), .Y(\u0\/u1\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1089_ ( .A(\u0\/u1\/_0281_ ), .B(\u0\/u1\/_0283_ ), .C(\u0\/u1\/_0284_ ), .D(\u0\/u1\/_0285_ ), .X(\u0\/u1\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1090_ ( .A(\u0\/u1\/_0082_ ), .B(\u0\/u1\/_0027_ ), .X(\u0\/u1\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1091_ ( .A(\u0\/u1\/_0129_ ), .B(\u0\/u1\/_0027_ ), .X(\u0\/u1\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_1092_ ( .A(\u0\/u1\/_0287_ ), .B(\u0\/u1\/_0288_ ), .Y(\u0\/u1\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1093_ ( .A1(\u0\/u1\/_0752_ ), .A2(\u0\/u1\/_0683_ ), .B1(\u0\/u1\/_0093_ ), .B2(\u0\/u1\/_0029_ ), .Y(\u0\/u1\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1094_ ( .A1(\u0\/u1\/_0092_ ), .A2(\u0\/u1\/_0575_ ), .B1(\u0\/u1\/_0056_ ), .Y(\u0\/u1\/_0291_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1096_ ( .A1(\u0\/u1\/_0218_ ), .A2(\u0\/u1\/_0662_ ), .B1(\u0\/u1\/_0084_ ), .B2(\u0\/u1\/_0056_ ), .Y(\u0\/u1\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1097_ ( .A(\u0\/u1\/_0289_ ), .B(\u0\/u1\/_0290_ ), .C(\u0\/u1\/_0291_ ), .D(\u0\/u1\/_0294_ ), .X(\u0\/u1\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1098_ ( .A(\u0\/u1\/_0750_ ), .B(\u0\/u1\/_0193_ ), .X(\u0\/u1\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1099_ ( .A(\u0\/u1\/_0705_ ), .B(\u0\/u1\/_0380_ ), .X(\u0\/u1\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1100_ ( .A(\u0\/u1\/_0752_ ), .B(\u0\/u1\/_0129_ ), .Y(\u0\/u1\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u1/_1101_ ( .A(\u0\/u1\/_0296_ ), .B(\u0\/u1\/_0297_ ), .C_N(\u0\/u1\/_0298_ ), .Y(\u0\/u1\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1102_ ( .A(\u0\/u1\/_0089_ ), .B(\u0\/u1\/_0532_ ), .Y(\u0\/u1\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1103_ ( .A(\w3\[10\] ), .Y(\u0\/u1\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u1/_1104_ ( .A(\u0\/u1\/_0301_ ), .B(\w3\[11\] ), .C(\u0\/u1\/_0118_ ), .Y(\u0\/u1\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1105_ ( .A(\u0\/u1\/_0072_ ), .B(\u0\/u1\/_0302_ ), .X(\u0\/u1\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1106_ ( .A(\u0\/u1\/_0303_ ), .Y(\u0\/u1\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1107_ ( .A(\u0\/u1\/_0147_ ), .B(\u0\/u1\/_0302_ ), .Y(\u0\/u1\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1108_ ( .A(\u0\/u1\/_0299_ ), .B(\u0\/u1\/_0300_ ), .C(\u0\/u1\/_0305_ ), .D(\u0\/u1\/_0306_ ), .X(\u0\/u1\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1109_ ( .A(\u0\/u1\/_0278_ ), .B(\u0\/u1\/_0286_ ), .C(\u0\/u1\/_0295_ ), .D(\u0\/u1\/_0307_ ), .X(\u0\/u1\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u1/_1110_ ( .A(\u0\/u1\/_0228_ ), .B(\u0\/u1\/_0265_ ), .C(\u0\/u1\/_0308_ ), .Y(\u0\/u1\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1111_ ( .A(\u0\/u1\/_0235_ ), .Y(\u0\/u1\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1112_ ( .A(\u0\/u1\/_0478_ ), .B(\u0\/u1\/_0640_ ), .X(\u0\/u1\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1113_ ( .A(\u0\/u1\/_0310_ ), .Y(\u0\/u1\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1114_ ( .A(\u0\/u1\/_0022_ ), .B(\u0\/u1\/_0218_ ), .Y(\u0\/u1\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1115_ ( .A(\u0\/u1\/_0218_ ), .B(\u0\/u1\/_0032_ ), .Y(\u0\/u1\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1116_ ( .A(\u0\/u1\/_0309_ ), .B(\u0\/u1\/_0311_ ), .C(\u0\/u1\/_0312_ ), .D(\u0\/u1\/_0313_ ), .X(\u0\/u1\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1117_ ( .A(\u0\/u1\/_0218_ ), .B(\u0\/u1\/_0064_ ), .Y(\u0\/u1\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1118_ ( .A(\u0\/u1\/_0218_ ), .B(\u0\/u1\/_0683_ ), .Y(\u0\/u1\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1119_ ( .A(\u0\/u1\/_0315_ ), .B(\u0\/u1\/_0316_ ), .C(\u0\/u1\/_0317_ ), .D(\u0\/u1\/_0253_ ), .X(\u0\/u1\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1120_ ( .A(\u0\/u1\/_0047_ ), .B(\u0\/u1\/_0304_ ), .Y(\u0\/u1\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1121_ ( .A(\u0\/u1\/_0586_ ), .B(\u0\/u1\/_0162_ ), .Y(\u0\/u1\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1122_ ( .A(\u0\/u1\/_0319_ ), .B(\u0\/u1\/_0320_ ), .Y(\u0\/u1\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_1123_ ( .A(\u0\/u1\/_0321_ ), .B(\u0\/u1\/_0238_ ), .Y(\u0\/u1\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1124_ ( .A(\u0\/u1\/_0304_ ), .B(\u0\/u1\/_0062_ ), .Y(\u0\/u1\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_1125_ ( .A(\u0\/u1\/_0251_ ), .X(\u0\/u1\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1126_ ( .A1(\u0\/u1\/_0324_ ), .A2(\u0\/u1\/_0084_ ), .B1(\u0\/u1\/_0255_ ), .Y(\u0\/u1\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1127_ ( .A1(\u0\/u1\/_0050_ ), .A2(\u0\/u1\/_0216_ ), .B1(\u0\/u1\/_0109_ ), .C1(\u0\/u1\/_0255_ ), .Y(\u0\/u1\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1128_ ( .A(\u0\/u1\/_0322_ ), .B(\u0\/u1\/_0323_ ), .C(\u0\/u1\/_0326_ ), .D(\u0\/u1\/_0327_ ), .X(\u0\/u1\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1129_ ( .A1(\u0\/u1\/_0733_ ), .A2(\u0\/u1\/_0279_ ), .A3(\u0\/u1\/_0058_ ), .B1(\u0\/u1\/_0056_ ), .Y(\u0\/u1\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_1130_ ( .A(\u0\/u1\/_0047_ ), .X(\u0\/u1\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1131_ ( .A(\u0\/u1\/_0330_ ), .B(\u0\/u1\/_0056_ ), .Y(\u0\/u1\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1132_ ( .A(\u0\/u1\/_0054_ ), .B(\u0\/u1\/_0045_ ), .Y(\u0\/u1\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1133_ ( .A(\u0\/u1\/_0329_ ), .B(\u0\/u1\/_0331_ ), .C(\u0\/u1\/_0284_ ), .D(\u0\/u1\/_0332_ ), .X(\u0\/u1\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u1/_1134_ ( .A1(\u0\/u1\/_0543_ ), .A2(\u0\/u1\/_0216_ ), .B1(\u0\/u1\/_0532_ ), .C1(\u0\/u1\/_0060_ ), .X(\u0\/u1\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1135_ ( .A(\u0\/u1\/_0084_ ), .B(\u0\/u1\/_0060_ ), .Y(\u0\/u1\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1136_ ( .A(\u0\/u1\/_0324_ ), .B(\u0\/u1\/_0060_ ), .Y(\u0\/u1\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1137_ ( .A(\u0\/u1\/_0335_ ), .B(\u0\/u1\/_0337_ ), .Y(\u0\/u1\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1138_ ( .A1(\u0\/u1\/_0276_ ), .A2(\u0\/u1\/_0060_ ), .B1(\u0\/u1\/_0334_ ), .C1(\u0\/u1\/_0338_ ), .Y(\u0\/u1\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1139_ ( .A(\u0\/u1\/_0318_ ), .B(\u0\/u1\/_0328_ ), .C(\u0\/u1\/_0333_ ), .D(\u0\/u1\/_0339_ ), .X(\u0\/u1\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u1/_1140_ ( .A1(\u0\/u1\/_0746_ ), .A2(\u0\/u1\/_0456_ ), .B1(\u0\/u1\/_0128_ ), .X(\u0\/u1\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u1/_1141_ ( .A_N(\u0\/u1\/_0086_ ), .B(\u0\/u1\/_0128_ ), .X(\u0\/u1\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1142_ ( .A(\u0\/u1\/_0079_ ), .B(\u0\/u1\/_0124_ ), .X(\u0\/u1\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_1143_ ( .A(\u0\/u1\/_0126_ ), .B(\u0\/u1\/_0343_ ), .Y(\u0\/u1\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u1/_1144_ ( .A(\u0\/u1\/_0341_ ), .B(\u0\/u1\/_0342_ ), .C_N(\u0\/u1\/_0344_ ), .Y(\u0\/u1\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1146_ ( .A1(\u0\/u1\/_0193_ ), .A2(\u0\/u1\/_0092_ ), .A3(\u0\/u1\/_0330_ ), .B1(\u0\/u1\/_0147_ ), .Y(\u0\/u1\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1147_ ( .A1(\u0\/u1\/_0130_ ), .A2(\u0\/u1\/_0084_ ), .A3(\u0\/u1\/_0456_ ), .B1(\u0\/u1\/_0139_ ), .Y(\u0\/u1\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1148_ ( .A1(\u0\/u1\/_0144_ ), .A2(\u0\/u1\/_0608_ ), .A3(\u0\/u1\/_0092_ ), .B1(\u0\/u1\/_0139_ ), .Y(\u0\/u1\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1149_ ( .A(\u0\/u1\/_0345_ ), .B(\u0\/u1\/_0348_ ), .C(\u0\/u1\/_0349_ ), .D(\u0\/u1\/_0350_ ), .X(\u0\/u1\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \u0/u1/_1150_ ( .A(\u0\/u1\/_0150_ ), .B(\u0\/u1\/_0194_ ), .C(\u0\/u1\/_0543_ ), .X(\u0\/u1\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u1/_1151_ ( .A(\u0\/u1\/_0277_ ), .SLEEP(\u0\/u1\/_0352_ ), .X(\u0\/u1\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \u0/u1/_1152_ ( .A1(\u0\/u1\/_0268_ ), .A2(\u0\/u1\/_0171_ ), .B1(\u0\/u1\/_0157_ ), .Y(\u0\/u1\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u1/_1153_ ( .A(\u0\/u1\/_0161_ ), .X(\u0\/u1\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1154_ ( .A1(\u0\/u1\/_0279_ ), .A2(\u0\/u1\/_0084_ ), .B1(\u0\/u1\/_0355_ ), .Y(\u0\/u1\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1155_ ( .A1(\u0\/u1\/_0020_ ), .A2(\u0\/u1\/_0193_ ), .A3(\u0\/u1\/_0091_ ), .B1(\u0\/u1\/_0355_ ), .Y(\u0\/u1\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1156_ ( .A(\u0\/u1\/_0353_ ), .B(\u0\/u1\/_0354_ ), .C(\u0\/u1\/_0356_ ), .D(\u0\/u1\/_0357_ ), .X(\u0\/u1\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1157_ ( .A(\u0\/u1\/_0111_ ), .B(\u0\/u1\/_0586_ ), .X(\u0\/u1\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1158_ ( .A(\u0\/u1\/_0360_ ), .Y(\u0\/u1\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u1/_1159_ ( .A1(\u0\/u1\/_0119_ ), .A2(\u0\/u1\/_0120_ ), .B1(\u0\/u1\/_0230_ ), .C1(\u0\/u1\/_0361_ ), .X(\u0\/u1\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1160_ ( .A1(\u0\/u1\/_0662_ ), .A2(\u0\/u1\/_0251_ ), .A3(\u0\/u1\/_0456_ ), .B1(\u0\/u1\/_0114_ ), .Y(\u0\/u1\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1162_ ( .A1(\u0\/u1\/_0035_ ), .A2(\u0\/u1\/_0251_ ), .A3(\u0\/u1\/_0456_ ), .B1(\u0\/u1\/_0099_ ), .Y(\u0\/u1\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1163_ ( .A1(\u0\/u1\/_0193_ ), .A2(\u0\/u1\/_0608_ ), .B1(\u0\/u1\/_0099_ ), .Y(\u0\/u1\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1164_ ( .A(\u0\/u1\/_0362_ ), .B(\u0\/u1\/_0363_ ), .C(\u0\/u1\/_0365_ ), .D(\u0\/u1\/_0366_ ), .X(\u0\/u1\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1165_ ( .A1(\u0\/u1\/_0575_ ), .A2(\u0\/u1\/_0092_ ), .A3(\u0\/u1\/_0330_ ), .B1(\u0\/u1\/_0089_ ), .Y(\u0\/u1\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1166_ ( .A1(\u0\/u1\/_0586_ ), .A2(\u0\/u1\/_0017_ ), .A3(\u0\/u1\/_0330_ ), .B1(\u0\/u1\/_0094_ ), .Y(\u0\/u1\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u1/_1167_ ( .A1(\u0\/u1\/_0293_ ), .A2(\u0\/u1\/_0456_ ), .B1(\u0\/u1\/_0089_ ), .Y(\u0\/u1\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1168_ ( .A1(\u0\/u1\/_0279_ ), .A2(\u0\/u1\/_0456_ ), .B1(\u0\/u1\/_0094_ ), .Y(\u0\/u1\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1169_ ( .A(\u0\/u1\/_0368_ ), .B(\u0\/u1\/_0370_ ), .C(\u0\/u1\/_0371_ ), .D(\u0\/u1\/_0372_ ), .X(\u0\/u1\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1170_ ( .A(\u0\/u1\/_0351_ ), .B(\u0\/u1\/_0359_ ), .C(\u0\/u1\/_0367_ ), .D(\u0\/u1\/_0373_ ), .X(\u0\/u1\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1171_ ( .A1(\u0\/u1\/_0102_ ), .A2(\u0\/u1\/_0347_ ), .B1(\u0\/u1\/_0109_ ), .C1(\u0\/u1\/_0029_ ), .Y(\u0\/u1\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1172_ ( .A1(\u0\/u1\/_0102_ ), .A2(\u0\/u1\/_0347_ ), .B1(\u0\/u1\/_0532_ ), .C1(\u0\/u1\/_0029_ ), .Y(\u0\/u1\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1173_ ( .A1(\u0\/u1\/_0050_ ), .A2(\u0\/u1\/_0543_ ), .B1(\u0\/u1\/_0380_ ), .C1(\u0\/u1\/_0029_ ), .Y(\u0\/u1\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1174_ ( .A(\u0\/u1\/_0041_ ), .B(\u0\/u1\/_0375_ ), .C(\u0\/u1\/_0376_ ), .D(\u0\/u1\/_0377_ ), .X(\u0\/u1\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1175_ ( .A(\u0\/u1\/_0047_ ), .B(\u0\/u1\/_0750_ ), .X(\u0\/u1\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1176_ ( .A(\u0\/u1\/_0379_ ), .Y(\u0\/u1\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1177_ ( .A(\u0\/u1\/_0016_ ), .B(\u0\/u1\/_0608_ ), .Y(\u0\/u1\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1178_ ( .A(\u0\/u1\/_0752_ ), .B(\u0\/u1\/_0554_ ), .Y(\u0\/u1\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1179_ ( .A1(\w3\[9\] ), .A2(\u0\/u1\/_0734_ ), .B1(\u0\/u1\/_0109_ ), .C1(\u0\/u1\/_0016_ ), .Y(\u0\/u1\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1180_ ( .A(\u0\/u1\/_0381_ ), .B(\u0\/u1\/_0382_ ), .C(\u0\/u1\/_0383_ ), .D(\u0\/u1\/_0384_ ), .X(\u0\/u1\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \u0/u1/_1181_ ( .A(\u0\/u1\/_0086_ ), .B_N(\u0\/u1\/_0736_ ), .X(\u0\/u1\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1182_ ( .A1(\u0\/u1\/_0748_ ), .A2(\u0\/u1\/_0456_ ), .B1(\u0\/u1\/_0739_ ), .Y(\u0\/u1\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1183_ ( .A1(\u0\/u1\/_0118_ ), .A2(\u0\/u1\/_0543_ ), .B1(\u0\/u1\/_0109_ ), .C1(\u0\/u1\/_0739_ ), .Y(\u0\/u1\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1184_ ( .A1(\u0\/u1\/_0102_ ), .A2(\u0\/u1\/_0301_ ), .B1(\w3\[11\] ), .C1(\u0\/u1\/_0739_ ), .Y(\u0\/u1\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1185_ ( .A(\u0\/u1\/_0386_ ), .B(\u0\/u1\/_0387_ ), .C(\u0\/u1\/_0388_ ), .D(\u0\/u1\/_0389_ ), .X(\u0\/u1\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1186_ ( .A(\u0\/u1\/_0020_ ), .Y(\u0\/u1\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1187_ ( .A(\u0\/u1\/_0727_ ), .Y(\u0\/u1\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1188_ ( .A(\u0\/u1\/_0727_ ), .B(\u0\/u1\/_0064_ ), .Y(\u0\/u1\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1189_ ( .A1(\u0\/u1\/_0102_ ), .A2(\u0\/u1\/_0734_ ), .B1(\u0\/u1\/_0532_ ), .C1(\u0\/u1\/_0727_ ), .Y(\u0\/u1\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u1/_1190_ ( .A1(\u0\/u1\/_0392_ ), .A2(\u0\/u1\/_0393_ ), .B1(\u0\/u1\/_0394_ ), .C1(\u0\/u1\/_0395_ ), .X(\u0\/u1\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1191_ ( .A(\u0\/u1\/_0378_ ), .B(\u0\/u1\/_0385_ ), .C(\u0\/u1\/_0390_ ), .D(\u0\/u1\/_0396_ ), .X(\u0\/u1\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u1/_1192_ ( .A(\u0\/u1\/_0340_ ), .B(\u0\/u1\/_0374_ ), .C(\u0\/u1\/_0397_ ), .Y(\u0\/u1\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1193_ ( .A(\u0\/u1\/_0077_ ), .B(\u0\/u1\/_0129_ ), .X(\u0\/u1\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_1194_ ( .A(\u0\/u1\/_0398_ ), .B(\u0\/u1\/_0239_ ), .Y(\u0\/u1\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1195_ ( .A(\u0\/u1\/_0022_ ), .B(\u0\/u1\/_0111_ ), .X(\u0\/u1\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u1/_1196_ ( .A_N(\u0\/u1\/_0400_ ), .B(\u0\/u1\/_0231_ ), .Y(\u0\/u1\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u1/_1197_ ( .A(\u0\/u1\/_0399_ ), .SLEEP(\u0\/u1\/_0402_ ), .X(\u0\/u1\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_1198_ ( .A(\u0\/u1\/_0746_ ), .B(\u0\/u1\/_0251_ ), .Y(\u0\/u1\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u1/_1199_ ( .A_N(\u0\/u1\/_0404_ ), .B(\u0\/u1\/_0752_ ), .Y(\u0\/u1\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \u0/u1/_1200_ ( .A(\u0\/u1\/_0467_ ), .B(\u0\/u1\/_0194_ ), .C(\u0\/u1\/_0694_ ), .X(\u0\/u1\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u1/_1201_ ( .A_N(\u0\/u1\/_0175_ ), .B(\u0\/u1\/_0406_ ), .X(\u0\/u1\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1202_ ( .A(\u0\/u1\/_0407_ ), .Y(\u0\/u1\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1203_ ( .A1(\u0\/u1\/_0094_ ), .A2(\u0\/u1\/_0197_ ), .B1(\u0\/u1\/_0114_ ), .B2(\u0\/u1\/_0640_ ), .Y(\u0\/u1\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1204_ ( .A(\u0\/u1\/_0403_ ), .B(\u0\/u1\/_0405_ ), .C(\u0\/u1\/_0408_ ), .D(\u0\/u1\/_0409_ ), .X(\u0\/u1\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1205_ ( .A(\u0\/u1\/_0030_ ), .B(\u0\/u1\/_0150_ ), .Y(\u0\/u1\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u1/_1206_ ( .A_N(\u0\/u1\/_0169_ ), .B(\u0\/u1\/_0289_ ), .C(\u0\/u1\/_0411_ ), .X(\u0\/u1\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u1/_1207_ ( .A1(\u0\/u1\/_0467_ ), .A2(\u0\/u1\/_0151_ ), .B1(\u0\/u1\/_0140_ ), .C1(\u0\/u1\/_0129_ ), .X(\u0\/u1\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1208_ ( .A1(\u0\/u1\/_0608_ ), .A2(\u0\/u1\/_0099_ ), .B1(\u0\/u1\/_0037_ ), .C1(\u0\/u1\/_0414_ ), .Y(\u0\/u1\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1209_ ( .A(\u0\/u1\/_0738_ ), .Y(\u0\/u1\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1210_ ( .A(\u0\/u1\/_0586_ ), .B(\u0\/u1\/_0736_ ), .Y(\u0\/u1\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1211_ ( .A1(\u0\/u1\/_0194_ ), .A2(\u0\/u1\/_0038_ ), .B1(\u0\/u1\/_0118_ ), .C1(\u0\/u1\/_0153_ ), .Y(\u0\/u1\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u1/_1212_ ( .A1(\u0\/u1\/_0416_ ), .A2(\u0\/u1\/_0117_ ), .B1(\u0\/u1\/_0417_ ), .C1(\u0\/u1\/_0418_ ), .X(\u0\/u1\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1213_ ( .A(\u0\/u1\/_0077_ ), .B(\u0\/u1\/_0035_ ), .X(\u0\/u1\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1214_ ( .A(\u0\/u1\/_0662_ ), .B(\u0\/u1\/_0124_ ), .Y(\u0\/u1\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1215_ ( .A(\u0\/u1\/_0030_ ), .B(\u0\/u1\/_0137_ ), .Y(\u0\/u1\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1216_ ( .A(\u0\/u1\/_0072_ ), .B(\u0\/u1\/_0731_ ), .Y(\u0\/u1\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u1/_1217_ ( .A_N(\u0\/u1\/_0420_ ), .B(\u0\/u1\/_0421_ ), .C(\u0\/u1\/_0422_ ), .D(\u0\/u1\/_0424_ ), .X(\u0\/u1\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1218_ ( .A(\u0\/u1\/_0413_ ), .B(\u0\/u1\/_0415_ ), .C(\u0\/u1\/_0419_ ), .D(\u0\/u1\/_0425_ ), .X(\u0\/u1\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u1/_1219_ ( .A(\u0\/u1\/_0355_ ), .B(\u0\/u1\/_0102_ ), .C(\u0\/u1\/_0109_ ), .Y(\u0\/u1\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1220_ ( .A(\u0\/u1\/_0077_ ), .B(\u0\/u1\/_0017_ ), .X(\u0\/u1\/_0428_ ) );
sky130_fd_sc_hd__and2_1 \u0/u1/_1221_ ( .A(\u0\/u1\/_0077_ ), .B(\u0\/u1\/_0554_ ), .X(\u0\/u1\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u1/_1222_ ( .A1(\u0\/u1\/_0050_ ), .A2(\u0\/u1\/_0216_ ), .B1(\u0\/u1\/_0380_ ), .C1(\u0\/u1\/_0078_ ), .X(\u0\/u1\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u1/_1223_ ( .A(\u0\/u1\/_0428_ ), .B(\u0\/u1\/_0429_ ), .C(\u0\/u1\/_0430_ ), .Y(\u0\/u1\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u1/_1224_ ( .A_N(\u0\/u1\/_0209_ ), .B(\u0\/u1\/_0431_ ), .X(\u0\/u1\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u1/_1225_ ( .A1(\u0\/u1\/_0215_ ), .A2(\u0\/u1\/_0404_ ), .B1(\u0\/u1\/_0427_ ), .C1(\u0\/u1\/_0432_ ), .X(\u0\/u1\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1226_ ( .A(\u0\/u1\/_0043_ ), .B(\u0\/u1\/_0058_ ), .Y(\u0\/u1\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1227_ ( .A(\u0\/u1\/_0195_ ), .B(\u0\/u1\/_0233_ ), .C(\u0\/u1\/_0320_ ), .D(\u0\/u1\/_0435_ ), .X(\u0\/u1\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1228_ ( .A(\u0\/u1\/_0261_ ), .B(\u0\/u1\/_0738_ ), .Y(\u0\/u1\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1229_ ( .A1(\u0\/u1\/_0218_ ), .A2(\u0\/u1\/_0640_ ), .B1(\u0\/u1\/_0261_ ), .B2(\u0\/u1\/_0056_ ), .Y(\u0\/u1\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1230_ ( .A(\u0\/u1\/_0436_ ), .B(\u0\/u1\/_0394_ ), .C(\u0\/u1\/_0437_ ), .D(\u0\/u1\/_0438_ ), .X(\u0\/u1\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1231_ ( .A(\u0\/u1\/_0410_ ), .B(\u0\/u1\/_0426_ ), .C(\u0\/u1\/_0433_ ), .D(\u0\/u1\/_0439_ ), .X(\u0\/u1\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u1/_1232_ ( .A(\u0\/u1\/_0135_ ), .SLEEP(\u0\/u1\/_0273_ ), .X(\u0\/u1\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1233_ ( .A1(\u0\/u1\/_0279_ ), .A2(\u0\/u1\/_0456_ ), .B1(\u0\/u1\/_0099_ ), .Y(\u0\/u1\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1234_ ( .A(\u0\/u1\/_0441_ ), .B(\u0\/u1\/_0164_ ), .C(\u0\/u1\/_0270_ ), .D(\u0\/u1\/_0442_ ), .X(\u0\/u1\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1235_ ( .A(\u0\/u1\/_0051_ ), .B(\u0\/u1\/_0662_ ), .Y(\u0\/u1\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1236_ ( .A(\u0\/u1\/_0051_ ), .B(\u0\/u1\/_0271_ ), .Y(\u0\/u1\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1237_ ( .A(\u0\/u1\/_0444_ ), .B(\u0\/u1\/_0446_ ), .X(\u0\/u1\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1238_ ( .A(\u0\/u1\/_0193_ ), .B(\u0\/u1\/_0304_ ), .X(\u0\/u1\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1239_ ( .A(\u0\/u1\/_0448_ ), .Y(\u0\/u1\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1240_ ( .A(\u0\/u1\/_0162_ ), .B(\u0\/u1\/_0130_ ), .X(\u0\/u1\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1241_ ( .A(\u0\/u1\/_0450_ ), .Y(\u0\/u1\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1242_ ( .A1(\u0\/u1\/_0129_ ), .A2(\u0\/u1\/_0554_ ), .B1(\u0\/u1\/_0043_ ), .Y(\u0\/u1\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1243_ ( .A(\u0\/u1\/_0447_ ), .B(\u0\/u1\/_0449_ ), .C(\u0\/u1\/_0451_ ), .D(\u0\/u1\/_0452_ ), .X(\u0\/u1\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1244_ ( .A(\u0\/u1\/_0056_ ), .B(\u0\/u1\/_0064_ ), .Y(\u0\/u1\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u1/_1245_ ( .A_N(\u0\/u1\/_0248_ ), .B(\u0\/u1\/_0454_ ), .C(\u0\/u1\/_0254_ ), .D(\u0\/u1\/_0256_ ), .X(\u0\/u1\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1246_ ( .A1(\u0\/u1\/_0330_ ), .A2(\u0\/u1\/_0099_ ), .B1(\u0\/u1\/_0456_ ), .B2(\u0\/u1\/_0705_ ), .Y(\u0\/u1\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1247_ ( .A1(\u0\/u1\/_0748_ ), .A2(\u0\/u1\/_0738_ ), .B1(\u0\/u1\/_0092_ ), .B2(\u0\/u1\/_0752_ ), .Y(\u0\/u1\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1248_ ( .A1(\u0\/u1\/_0072_ ), .A2(\u0\/u1\/_0035_ ), .B1(\u0\/u1\/_0748_ ), .B2(\u0\/u1\/_0056_ ), .Y(\u0\/u1\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1249_ ( .A1(\u0\/u1\/_0748_ ), .A2(\u0\/u1\/_0251_ ), .B1(\u0\/u1\/_0029_ ), .Y(\u0\/u1\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1250_ ( .A(\u0\/u1\/_0457_ ), .B(\u0\/u1\/_0458_ ), .C(\u0\/u1\/_0459_ ), .D(\u0\/u1\/_0460_ ), .X(\u0\/u1\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1251_ ( .A(\u0\/u1\/_0443_ ), .B(\u0\/u1\/_0453_ ), .C(\u0\/u1\/_0455_ ), .D(\u0\/u1\/_0461_ ), .X(\u0\/u1\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1252_ ( .A(\u0\/u1\/_0705_ ), .B(\u0\/u1\/_0079_ ), .X(\u0\/u1\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1253_ ( .A(\u0\/u1\/_0586_ ), .B(\u0\/u1\/_0124_ ), .Y(\u0\/u1\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1254_ ( .A(\u0\/u1\/_0218_ ), .B(\u0\/u1\/_0746_ ), .Y(\u0\/u1\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u1/_1255_ ( .A_N(\u0\/u1\/_0463_ ), .B(\u0\/u1\/_0464_ ), .C(\u0\/u1\/_0465_ ), .X(\u0\/u1\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u1/_1256_ ( .A1(\u0\/u1\/_0271_ ), .A2(\u0\/u1\/_0072_ ), .B1(\u0\/u1\/_0142_ ), .B2(\u0\/u1\/_0027_ ), .X(\u0\/u1\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1257_ ( .A1(\u0\/u1\/_0144_ ), .A2(\u0\/u1\/_0099_ ), .B1(\u0\/u1\/_0360_ ), .C1(\u0\/u1\/_0468_ ), .Y(\u0\/u1\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u1/_1258_ ( .A1(\u0\/u1\/_0662_ ), .A2(\u0\/u1\/_0251_ ), .B1(\u0\/u1\/_0218_ ), .X(\u0\/u1\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1259_ ( .A1(\u0\/u1\/_0575_ ), .A2(\u0\/u1\/_0056_ ), .B1(\u0\/u1\/_0379_ ), .C1(\u0\/u1\/_0470_ ), .Y(\u0\/u1\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1260_ ( .A(\u0\/u1\/_0466_ ), .B(\u0\/u1\/_0469_ ), .C(\u0\/u1\/_0471_ ), .D(\u0\/u1\/_0305_ ), .X(\u0\/u1\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u1/_1261_ ( .A1(\u0\/u1\/_0029_ ), .A2(\u0\/u1\/_0683_ ), .B1(\u0\/u1\/_0324_ ), .B2(\u0\/u1\/_0056_ ), .X(\u0\/u1\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1262_ ( .A(\u0\/u1\/_0084_ ), .B(\u0\/u1\/_0099_ ), .X(\u0\/u1\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \u0/u1/_1263_ ( .A1(\u0\/u1\/_0092_ ), .A2(\u0\/u1\/_0029_ ), .B1(\u0\/u1\/_0474_ ), .X(\u0\/u1\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u1/_1264_ ( .A(\u0\/u1\/_0075_ ), .B(\u0\/u1\/_0473_ ), .C(\u0\/u1\/_0475_ ), .Y(\u0\/u1\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1265_ ( .A1(\u0\/u1\/_0279_ ), .A2(\u0\/u1\/_0255_ ), .B1(\u0\/u1\/_0084_ ), .B2(\u0\/u1\/_0060_ ), .Y(\u0\/u1\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1266_ ( .A1(\u0\/u1\/_0093_ ), .A2(\u0\/u1\/_0056_ ), .B1(\u0\/u1\/_0456_ ), .B2(\u0\/u1\/_0114_ ), .Y(\u0\/u1\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1267_ ( .A1(\u0\/u1\/_0161_ ), .A2(\u0\/u1\/_0032_ ), .B1(\u0\/u1\/_0324_ ), .B2(\u0\/u1\/_0147_ ), .Y(\u0\/u1\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1268_ ( .A1(\u0\/u1\/_0054_ ), .A2(\u0\/u1\/_0731_ ), .B1(\u0\/u1\/_0748_ ), .B2(\u0\/u1\/_0304_ ), .Y(\u0\/u1\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1269_ ( .A(\u0\/u1\/_0477_ ), .B(\u0\/u1\/_0479_ ), .C(\u0\/u1\/_0480_ ), .D(\u0\/u1\/_0481_ ), .X(\u0\/u1\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1270_ ( .A(\u0\/u1\/_0161_ ), .B(\u0\/u1\/_0064_ ), .Y(\u0\/u1\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u1/_1271_ ( .A(\u0\/u1\/_0731_ ), .B(\u0\/u1\/_0123_ ), .C(\u0\/u1\/_0467_ ), .Y(\u0\/u1\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1272_ ( .A(\u0\/u1\/_0483_ ), .B(\u0\/u1\/_0484_ ), .Y(\u0\/u1\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1273_ ( .A(\u0\/u1\/_0297_ ), .Y(\u0\/u1\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u1/_1274_ ( .A_N(\u0\/u1\/_0485_ ), .B(\u0\/u1\/_0181_ ), .C(\u0\/u1\/_0486_ ), .D(\u0\/u1\/_0386_ ), .X(\u0\/u1\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1275_ ( .A(\u0\/u1\/_0472_ ), .B(\u0\/u1\/_0476_ ), .C(\u0\/u1\/_0482_ ), .D(\u0\/u1\/_0487_ ), .X(\u0\/u1\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u1/_1276_ ( .A(\u0\/u1\/_0440_ ), .B(\u0\/u1\/_0462_ ), .C(\u0\/u1\/_0488_ ), .Y(\u0\/u1\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1277_ ( .A(\u0\/u1\/_0403_ ), .B(\u0\/u1\/_0230_ ), .C(\u0\/u1\/_0451_ ), .D(\u0\/u1\/_0361_ ), .X(\u0\/u1\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1278_ ( .A1(\u0\/u1\/_0118_ ), .A2(\u0\/u1\/_0050_ ), .B1(\u0\/u1\/_0109_ ), .C1(\u0\/u1\/_0139_ ), .Y(\u0\/u1\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1279_ ( .A(\u0\/u1\/_0447_ ), .B(\u0\/u1\/_0437_ ), .C(\u0\/u1\/_0491_ ), .D(\u0\/u1\/_0427_ ), .X(\u0\/u1\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1280_ ( .A1(\u0\/u1\/_0084_ ), .A2(\u0\/u1\/_0255_ ), .B1(\u0\/u1\/_0608_ ), .B2(\u0\/u1\/_0029_ ), .Y(\u0\/u1\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1281_ ( .A1(\u0\/u1\/_0144_ ), .A2(\u0\/u1\/_0147_ ), .B1(\u0\/u1\/_0355_ ), .B2(\u0\/u1\/_0093_ ), .Y(\u0\/u1\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1282_ ( .A1(\u0\/u1\/_0705_ ), .A2(\u0\/u1\/_0279_ ), .B1(\u0\/u1\/_0330_ ), .B2(\u0\/u1\/_0029_ ), .Y(\u0\/u1\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1283_ ( .A1(\u0\/u1\/_0279_ ), .A2(\u0\/u1\/_0084_ ), .B1(\u0\/u1\/_0114_ ), .Y(\u0\/u1\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1284_ ( .A(\u0\/u1\/_0493_ ), .B(\u0\/u1\/_0494_ ), .C(\u0\/u1\/_0495_ ), .D(\u0\/u1\/_0496_ ), .X(\u0\/u1\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1285_ ( .A1(\u0\/u1\/_0456_ ), .A2(\u0\/u1\/_0137_ ), .B1(\u0\/u1\/_0355_ ), .B2(\u0\/u1\/_0575_ ), .Y(\u0\/u1\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1286_ ( .A1(\u0\/u1\/_0099_ ), .A2(\u0\/u1\/_0733_ ), .B1(\u0\/u1\/_0093_ ), .B2(\u0\/u1\/_0218_ ), .Y(\u0\/u1\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1287_ ( .A(\u0\/u1\/_0147_ ), .B(\u0\/u1\/_0640_ ), .Y(\u0\/u1\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1288_ ( .A1(\u0\/u1\/_0153_ ), .A2(\u0\/u1\/_0056_ ), .B1(\u0\/u1\/_0748_ ), .Y(\u0\/u1\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1289_ ( .A(\u0\/u1\/_0498_ ), .B(\u0\/u1\/_0500_ ), .C(\u0\/u1\/_0501_ ), .D(\u0\/u1\/_0502_ ), .X(\u0\/u1\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1290_ ( .A(\u0\/u1\/_0490_ ), .B(\u0\/u1\/_0492_ ), .C(\u0\/u1\/_0497_ ), .D(\u0\/u1\/_0503_ ), .X(\u0\/u1\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u1/_1291_ ( .A_N(\u0\/u1\/_0275_ ), .B(\u0\/u1\/_0705_ ), .X(\u0\/u1\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1292_ ( .A(\u0\/u1\/_0505_ ), .Y(\u0\/u1\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1293_ ( .A(\u0\/u1\/_0380_ ), .B(\u0\/u1\/_0347_ ), .X(\u0\/u1\/_0507_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u1/_1294_ ( .A1(\u0\/u1\/_0507_ ), .A2(\u0\/u1\/_0093_ ), .B1(\u0\/u1\/_0056_ ), .Y(\u0\/u1\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1295_ ( .A(\u0\/u1\/_0322_ ), .B(\u0\/u1\/_0277_ ), .C(\u0\/u1\/_0506_ ), .D(\u0\/u1\/_0508_ ), .X(\u0\/u1\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1296_ ( .A(\u0\/u1\/_0084_ ), .B(\u0\/u1\/_0705_ ), .X(\u0\/u1\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1297_ ( .A1(\u0\/u1\/_0733_ ), .A2(\u0\/u1\/_0114_ ), .B1(\u0\/u1\/_0429_ ), .C1(\u0\/u1\/_0511_ ), .Y(\u0\/u1\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_1298_ ( .A(\u0\/u1\/_0019_ ), .B(\u0\/u1\/_0024_ ), .Y(\u0\/u1\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1299_ ( .A(\u0\/u1\/_0512_ ), .B(\u0\/u1\/_0513_ ), .C(\u0\/u1\/_0742_ ), .D(\u0\/u1\/_0306_ ), .X(\u0\/u1\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1300_ ( .A1(\u0\/u1\/_0532_ ), .A2(\u0\/u1\/_0089_ ), .B1(\u0\/u1\/_0154_ ), .C1(\u0\/u1\/_0169_ ), .Y(\u0\/u1\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u1/_1301_ ( .A1(\u0\/u1\/_0749_ ), .A2(\u0\/u1\/_0026_ ), .B1(\u0\/u1\/_0069_ ), .C1(\u0\/u1\/_0032_ ), .X(\u0\/u1\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u1/_1302_ ( .A1(\u0\/u1\/_0324_ ), .A2(\u0\/u1\/_0355_ ), .B1(\u0\/u1\/_0330_ ), .B2(\u0\/u1\/_0727_ ), .X(\u0\/u1\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u1/_1303_ ( .A(\u0\/u1\/_0133_ ), .B(\u0\/u1\/_0516_ ), .C(\u0\/u1\/_0517_ ), .Y(\u0\/u1\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1304_ ( .A(\u0\/u1\/_0509_ ), .B(\u0\/u1\/_0514_ ), .C(\u0\/u1\/_0515_ ), .D(\u0\/u1\/_0518_ ), .X(\u0\/u1\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1305_ ( .A(\u0\/u1\/_0746_ ), .B(\u0\/u1\/_0072_ ), .Y(\u0\/u1\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1306_ ( .A1(\u0\/u1\/_0082_ ), .A2(\u0\/u1\/_0070_ ), .B1(\u0\/u1\/_0043_ ), .B2(\u0\/u1\/_0193_ ), .Y(\u0\/u1\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1307_ ( .A(\u0\/u1\/_0311_ ), .B(\u0\/u1\/_0520_ ), .C(\u0\/u1\/_0332_ ), .D(\u0\/u1\/_0522_ ), .X(\u0\/u1\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1308_ ( .A(\u0\/u1\/_0129_ ), .B(\u0\/u1\/_0218_ ), .X(\u0\/u1\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_1309_ ( .A(\u0\/u1\/_0235_ ), .B(\u0\/u1\/_0524_ ), .Y(\u0\/u1\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u1/_1310_ ( .A(\u0\/u1\/_0081_ ), .B(\u0\/u1\/_0085_ ), .Y(\u0\/u1\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1311_ ( .A1(\u0\/u1\/_0051_ ), .A2(\u0\/u1\/_0045_ ), .B1(\u0\/u1\/_0130_ ), .B2(\u0\/u1\/_0094_ ), .Y(\u0\/u1\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1312_ ( .A(\u0\/u1\/_0523_ ), .B(\u0\/u1\/_0525_ ), .C(\u0\/u1\/_0526_ ), .D(\u0\/u1\/_0527_ ), .X(\u0\/u1\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u1/_1313_ ( .A_N(\u0\/u1\/_0250_ ), .B(\u0\/u1\/_0521_ ), .Y(\u0\/u1\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1314_ ( .A(\u0\/u1\/_0128_ ), .B(\u0\/u1\/_0020_ ), .X(\u0\/u1\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1315_ ( .A(\u0\/u1\/_0530_ ), .Y(\u0\/u1\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1316_ ( .A(\u0\/u1\/_0099_ ), .B(\u0\/u1\/_0058_ ), .X(\u0\/u1\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1317_ ( .A(\u0\/u1\/_0533_ ), .Y(\u0\/u1\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u1/_1318_ ( .A_N(\u0\/u1\/_0529_ ), .B(\u0\/u1\/_0531_ ), .C(\u0\/u1\/_0534_ ), .D(\u0\/u1\/_0192_ ), .X(\u0\/u1\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1319_ ( .A(\u0\/u1\/_0434_ ), .B(\u0\/u1\/_0078_ ), .X(\u0\/u1\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u1/_1320_ ( .A1(\u0\/u1\/_0750_ ), .A2(\u0\/u1\/_0079_ ), .B1(\u0\/u1\/_0129_ ), .B2(\u0\/u1\/_0705_ ), .X(\u0\/u1\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1321_ ( .A1(\u0\/u1\/_0161_ ), .A2(\u0\/u1\/_0032_ ), .B1(\u0\/u1\/_0536_ ), .C1(\u0\/u1\/_0537_ ), .Y(\u0\/u1\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u1/_1322_ ( .A1(\u0\/u1\/_0746_ ), .A2(\u0\/u1\/_0162_ ), .B1(\u0\/u1\/_0079_ ), .B2(\u0\/u1\/_0043_ ), .X(\u0\/u1\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1323_ ( .A1(\u0\/u1\/_0093_ ), .A2(\u0\/u1\/_0029_ ), .B1(\u0\/u1\/_0240_ ), .C1(\u0\/u1\/_0539_ ), .Y(\u0\/u1\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1324_ ( .A(\u0\/u1\/_0434_ ), .B(\u0\/u1\/_0043_ ), .X(\u0\/u1\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u1/_1325_ ( .A1(\u0\/u1\/_0142_ ), .A2(\u0\/u1\/_0150_ ), .B1(\u0\/u1\/_0022_ ), .B2(\u0\/u1\/_0137_ ), .X(\u0\/u1\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1326_ ( .A1(\u0\/u1\/_0279_ ), .A2(\u0\/u1\/_0051_ ), .B1(\u0\/u1\/_0541_ ), .C1(\u0\/u1\/_0542_ ), .Y(\u0\/u1\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1327_ ( .A(\u0\/u1\/_0159_ ), .B(\u0\/u1\/_0035_ ), .X(\u0\/u1\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u1/_1328_ ( .A1(\u0\/u1\/_0271_ ), .A2(\u0\/u1\/_0434_ ), .B1(\u0\/u1\/_0027_ ), .X(\u0\/u1\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1329_ ( .A1(\u0\/u1\/_0091_ ), .A2(\u0\/u1\/_0128_ ), .B1(\u0\/u1\/_0545_ ), .C1(\u0\/u1\/_0546_ ), .Y(\u0\/u1\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1330_ ( .A(\u0\/u1\/_0538_ ), .B(\u0\/u1\/_0540_ ), .C(\u0\/u1\/_0544_ ), .D(\u0\/u1\/_0547_ ), .X(\u0\/u1\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1331_ ( .A(\u0\/u1\/_0099_ ), .B(\u0\/u1\/_0193_ ), .X(\u0\/u1\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u1/_1332_ ( .A(\u0\/u1\/_0549_ ), .B(\u0\/u1\/_0186_ ), .C(\u0\/u1\/_0187_ ), .Y(\u0\/u1\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1333_ ( .A(\u0\/u1\/_0062_ ), .B(\u0\/u1\/_0347_ ), .C(\u0\/u1\/_0749_ ), .D(\u0\/u1\/_0694_ ), .X(\u0\/u1\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1334_ ( .A1(\u0\/u1\/_0130_ ), .A2(\u0\/u1\/_0218_ ), .B1(\u0\/u1\/_0551_ ), .C1(\u0\/u1\/_0101_ ), .Y(\u0\/u1\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1335_ ( .A(\u0\/u1\/_0139_ ), .B(\u0\/u1\/_0640_ ), .Y(\u0\/u1\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1336_ ( .A1(\u0\/u1\/_0752_ ), .A2(\u0\/u1\/_0662_ ), .B1(\u0\/u1\/_0084_ ), .B2(\u0\/u1\/_0099_ ), .Y(\u0\/u1\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1337_ ( .A(\u0\/u1\/_0550_ ), .B(\u0\/u1\/_0552_ ), .C(\u0\/u1\/_0553_ ), .D(\u0\/u1\/_0555_ ), .X(\u0\/u1\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1338_ ( .A(\u0\/u1\/_0528_ ), .B(\u0\/u1\/_0535_ ), .C(\u0\/u1\/_0548_ ), .D(\u0\/u1\/_0556_ ), .X(\u0\/u1\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u1/_1339_ ( .A(\u0\/u1\/_0504_ ), .B(\u0\/u1\/_0519_ ), .C(\u0\/u1\/_0557_ ), .Y(\u0\/u1\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1340_ ( .A(\u0\/u1\/_0054_ ), .B(\u0\/u1\/_0507_ ), .X(\u0\/u1\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u1/_1341_ ( .A_N(\u0\/u1\/_0558_ ), .B(\u0\/u1\/_0408_ ), .C(\u0\/u1\/_0451_ ), .D(\u0\/u1\/_0452_ ), .X(\u0\/u1\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1342_ ( .A(\u0\/u1\/_0549_ ), .Y(\u0\/u1\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1343_ ( .A(\u0\/u1\/_0559_ ), .B(\u0\/u1\/_0403_ ), .C(\u0\/u1\/_0560_ ), .D(\u0\/u1\/_0371_ ), .X(\u0\/u1\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1344_ ( .A(\u0\/u1\/_0181_ ), .B(\u0\/u1\/_0178_ ), .X(\u0\/u1\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1345_ ( .A(\u0\/u1\/_0562_ ), .B(\u0\/u1\/_0552_ ), .C(\u0\/u1\/_0553_ ), .D(\u0\/u1\/_0555_ ), .X(\u0\/u1\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1346_ ( .A(\u0\/u1\/_0029_ ), .B(\u0\/u1\/_0020_ ), .Y(\u0\/u1\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1347_ ( .A(\u0\/u1\/_0051_ ), .B(\u0\/u1\/_0130_ ), .X(\u0\/u1\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1348_ ( .A(\u0\/u1\/_0566_ ), .Y(\u0\/u1\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1349_ ( .A(\u0\/u1\/_0159_ ), .B(\u0\/u1\/_0412_ ), .X(\u0\/u1\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1350_ ( .A1(\u0\/u1\/_0752_ ), .A2(\u0\/u1\/_0640_ ), .B1(\u0\/u1\/_0568_ ), .B2(\u0\/u1\/_0175_ ), .Y(\u0\/u1\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1351_ ( .A(\u0\/u1\/_0076_ ), .B(\u0\/u1\/_0565_ ), .C(\u0\/u1\/_0567_ ), .D(\u0\/u1\/_0569_ ), .X(\u0\/u1\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u1/_1352_ ( .A1(\u0\/u1\/_0035_ ), .A2(\u0\/u1\/_0142_ ), .B1(\u0\/u1\/_0161_ ), .X(\u0\/u1\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1353_ ( .A(\u0\/u1\/_0099_ ), .B(\u0\/u1\/_0662_ ), .Y(\u0\/u1\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u1/_1354_ ( .A(\u0\/u1\/_0420_ ), .B(\u0\/u1\/_0571_ ), .C_N(\u0\/u1\/_0572_ ), .Y(\u0\/u1\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1355_ ( .A(\u0\/u1\/_0051_ ), .B(\u0\/u1\/_0746_ ), .Y(\u0\/u1\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1356_ ( .A(\u0\/u1\/_0574_ ), .B(\u0\/u1\/_0319_ ), .C(\u0\/u1\/_0320_ ), .D(\u0\/u1\/_0411_ ), .X(\u0\/u1\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1357_ ( .A(\u0\/u1\/_0736_ ), .B(\u0\/u1\/_0035_ ), .Y(\u0\/u1\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1358_ ( .A(\u0\/u1\/_0736_ ), .B(\u0\/u1\/_0030_ ), .Y(\u0\/u1\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1359_ ( .A(\u0\/u1\/_0298_ ), .B(\u0\/u1\/_0208_ ), .C(\u0\/u1\/_0577_ ), .D(\u0\/u1\/_0578_ ), .X(\u0\/u1\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1360_ ( .A1(\u0\/u1\/_0020_ ), .A2(\u0\/u1\/_0137_ ), .B1(\u0\/u1\/_0261_ ), .B2(\u0\/u1\/_0128_ ), .Y(\u0\/u1\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1361_ ( .A(\u0\/u1\/_0573_ ), .B(\u0\/u1\/_0576_ ), .C(\u0\/u1\/_0579_ ), .D(\u0\/u1\/_0580_ ), .X(\u0\/u1\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1362_ ( .A(\u0\/u1\/_0561_ ), .B(\u0\/u1\/_0563_ ), .C(\u0\/u1\/_0570_ ), .D(\u0\/u1\/_0581_ ), .X(\u0\/u1\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1363_ ( .A(\u0\/u1\/_0128_ ), .B(\u0\/u1\/_0193_ ), .X(\u0\/u1\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1364_ ( .A(\u0\/u1\/_0082_ ), .B(\u0\/u1\/_0162_ ), .X(\u0\/u1\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u1/_1365_ ( .A(\u0\/u1\/_0583_ ), .B(\u0\/u1\/_0584_ ), .C_N(\u0\/u1\/_0437_ ), .Y(\u0\/u1\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u1/_1366_ ( .A(\u0\/u1\/_0150_ ), .B(\u0\/u1\/_0118_ ), .C(\u0\/u1\/_0380_ ), .Y(\u0\/u1\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u1/_1367_ ( .A_N(\u0\/u1\/_0182_ ), .B(\u0\/u1\/_0587_ ), .C(\u0\/u1\/_0323_ ), .X(\u0\/u1\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1368_ ( .A1(\u0\/u1\/_0575_ ), .A2(\u0\/u1\/_0153_ ), .B1(\u0\/u1\/_0727_ ), .B2(\u0\/u1\/_0058_ ), .Y(\u0\/u1\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1369_ ( .A1(\u0\/u1\/_0218_ ), .A2(\u0\/u1\/_0064_ ), .B1(\u0\/u1\/_0456_ ), .B2(\u0\/u1\/_0255_ ), .Y(\u0\/u1\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1370_ ( .A(\u0\/u1\/_0585_ ), .B(\u0\/u1\/_0588_ ), .C(\u0\/u1\/_0589_ ), .D(\u0\/u1\/_0590_ ), .X(\u0\/u1\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \u0/u1/_1371_ ( .A1(\u0\/u1\/_0091_ ), .A2(\u0\/u1\/_0139_ ), .B1(\u0\/u1\/_0250_ ), .Y(\u0\/u1\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1372_ ( .A1(\u0\/u1\/_0092_ ), .A2(\u0\/u1\/_0739_ ), .B1(\u0\/u1\/_0324_ ), .B2(\u0\/u1\/_0029_ ), .Y(\u0\/u1\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1373_ ( .A1(\u0\/u1\/_0144_ ), .A2(\u0\/u1\/_0153_ ), .B1(\u0\/u1\/_0683_ ), .B2(\u0\/u1\/_0056_ ), .Y(\u0\/u1\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1374_ ( .A1(\u0\/u1\/_0091_ ), .A2(\u0\/u1\/_0218_ ), .B1(\u0\/u1\/_0330_ ), .B2(\u0\/u1\/_0056_ ), .Y(\u0\/u1\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1375_ ( .A(\u0\/u1\/_0592_ ), .B(\u0\/u1\/_0593_ ), .C(\u0\/u1\/_0594_ ), .D(\u0\/u1\/_0595_ ), .X(\u0\/u1\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1376_ ( .A(\u0\/u1\/_0218_ ), .B(\u0\/u1\/_0144_ ), .Y(\u0\/u1\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1377_ ( .A(\u0\/u1\/_0312_ ), .B(\u0\/u1\/_0598_ ), .Y(\u0\/u1\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1378_ ( .A(\u0\/u1\/_0575_ ), .B(\u0\/u1\/_0147_ ), .Y(\u0\/u1\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1379_ ( .A1(\u0\/u1\/_0293_ ), .A2(\u0\/u1\/_0137_ ), .B1(\u0\/u1\/_0093_ ), .B2(\u0\/u1\/_0739_ ), .Y(\u0\/u1\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1380_ ( .A1(\u0\/u1\/_0734_ ), .A2(\u0\/u1\/_0531_ ), .B1(\u0\/u1\/_0600_ ), .C1(\u0\/u1\/_0601_ ), .Y(\u0\/u1\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1381_ ( .A1(\u0\/u1\/_0153_ ), .A2(\u0\/u1\/_0261_ ), .B1(\u0\/u1\/_0599_ ), .C1(\u0\/u1\/_0602_ ), .Y(\u0\/u1\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1382_ ( .A(\u0\/u1\/_0591_ ), .B(\u0\/u1\/_0596_ ), .C(\u0\/u1\/_0174_ ), .D(\u0\/u1\/_0603_ ), .X(\u0\/u1\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1383_ ( .A(\u0\/u1\/_0029_ ), .B(\u0\/u1\/_0144_ ), .Y(\u0\/u1\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1384_ ( .A(\u0\/u1\/_0113_ ), .B(\u0\/u1\/_0017_ ), .Y(\u0\/u1\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1385_ ( .A(\u0\/u1\/_0381_ ), .B(\u0\/u1\/_0605_ ), .C(\u0\/u1\/_0361_ ), .D(\u0\/u1\/_0606_ ), .X(\u0\/u1\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1386_ ( .A1(\u0\/u1\/_0016_ ), .A2(\u0\/u1\/_0727_ ), .B1(\u0\/u1\/_0733_ ), .Y(\u0\/u1\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1387_ ( .A1(\u0\/u1\/_0586_ ), .A2(\u0\/u1\/_0159_ ), .B1(\u0\/u1\/_0082_ ), .B2(\u0\/u1\/_0750_ ), .Y(\u0\/u1\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1388_ ( .A1(\u0\/u1\/_0142_ ), .A2(\u0\/u1\/_0162_ ), .B1(\u0\/u1\/_0079_ ), .B2(\u0\/u1\/_0054_ ), .Y(\u0\/u1\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1389_ ( .A(\u0\/u1\/_0610_ ), .B(\u0\/u1\/_0611_ ), .C(\u0\/u1\/_0105_ ), .D(\u0\/u1\/_0106_ ), .X(\u0\/u1\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1390_ ( .A1(\u0\/u1\/_0094_ ), .A2(\u0\/u1\/_0302_ ), .B1(\u0\/u1\/_0324_ ), .B2(\u0\/u1\/_0089_ ), .Y(\u0\/u1\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1391_ ( .A(\u0\/u1\/_0607_ ), .B(\u0\/u1\/_0609_ ), .C(\u0\/u1\/_0612_ ), .D(\u0\/u1\/_0613_ ), .X(\u0\/u1\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1392_ ( .A(\u0\/u1\/_0041_ ), .B(\u0\/u1\/_0170_ ), .X(\u0\/u1\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1393_ ( .A(\u0\/u1\/_0554_ ), .B(\u0\/u1\/_0027_ ), .X(\u0\/u1\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1394_ ( .A(\u0\/u1\/_0027_ ), .B(\u0\/u1\/_0261_ ), .Y(\u0\/u1\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u1/_1395_ ( .A_N(\u0\/u1\/_0616_ ), .B(\u0\/u1\/_0617_ ), .Y(\u0\/u1\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1396_ ( .A1(\u0\/u1\/_0147_ ), .A2(\u0\/u1\/_0302_ ), .B1(\u0\/u1\/_0342_ ), .C1(\u0\/u1\/_0618_ ), .Y(\u0\/u1\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1397_ ( .A(\u0\/u1\/_0614_ ), .B(\u0\/u1\/_0272_ ), .C(\u0\/u1\/_0615_ ), .D(\u0\/u1\/_0620_ ), .X(\u0\/u1\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u1/_1398_ ( .A(\u0\/u1\/_0582_ ), .B(\u0\/u1\/_0604_ ), .C(\u0\/u1\/_0621_ ), .Y(\u0\/u1\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1399_ ( .A1(\u0\/u1\/_0084_ ), .A2(\u0\/u1\/_0456_ ), .B1(\u0\/u1\/_0089_ ), .Y(\u0\/u1\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1400_ ( .A1(\u0\/u1\/_0144_ ), .A2(\u0\/u1\/_0608_ ), .A3(\u0\/u1\/_0330_ ), .B1(\u0\/u1\/_0089_ ), .Y(\u0\/u1\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1401_ ( .A1(\u0\/u1\/_0197_ ), .A2(\u0\/u1\/_0130_ ), .A3(\u0\/u1\/_0110_ ), .B1(\u0\/u1\/_0094_ ), .Y(\u0\/u1\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1402_ ( .A(\u0\/u1\/_0432_ ), .B(\u0\/u1\/_0622_ ), .C(\u0\/u1\/_0623_ ), .D(\u0\/u1\/_0624_ ), .X(\u0\/u1\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \u0/u1/_1403_ ( .A1(\u0\/u1\/_0554_ ), .A2(\u0\/u1\/_0017_ ), .A3(\u0\/u1\/_0022_ ), .B1(\u0\/u1\/_0161_ ), .X(\u0\/u1\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u1/_1404_ ( .A_N(\u0\/u1\/_0269_ ), .B(\u0\/u1\/_0170_ ), .X(\u0\/u1\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1405_ ( .A1(\u0\/u1\/_0109_ ), .A2(\u0\/u1\/_0064_ ), .A3(\u0\/u1\/_0733_ ), .B1(\u0\/u1\/_0355_ ), .Y(\u0\/u1\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u1/_1406_ ( .A_N(\u0\/u1\/_0626_ ), .B(\u0\/u1\/_0627_ ), .C(\u0\/u1\/_0353_ ), .D(\u0\/u1\/_0628_ ), .X(\u0\/u1\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1407_ ( .A1(\u0\/u1\/_0091_ ), .A2(\u0\/u1\/_0110_ ), .A3(\u0\/u1\/_0176_ ), .B1(\u0\/u1\/_0139_ ), .Y(\u0\/u1\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1408_ ( .A1(\u0\/u1\/_0020_ ), .A2(\u0\/u1\/_0261_ ), .B1(\u0\/u1\/_0147_ ), .Y(\u0\/u1\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1409_ ( .A(\u0\/u1\/_0631_ ), .B(\u0\/u1\/_0344_ ), .C(\u0\/u1\/_0421_ ), .D(\u0\/u1\/_0632_ ), .X(\u0\/u1\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u1/_1410_ ( .A1(\u0\/u1\/_0325_ ), .A2(\u0\/u1\/_0734_ ), .B1(\u0\/u1\/_0038_ ), .C1(\u0\/u1\/_0113_ ), .X(\u0\/u1\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1411_ ( .A1(\u0\/u1\/_0456_ ), .A2(\u0\/u1\/_0114_ ), .B1(\u0\/u1\/_0221_ ), .C1(\u0\/u1\/_0634_ ), .Y(\u0\/u1\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u1/_1412_ ( .A(\u0\/u1\/_0119_ ), .B_N(\u0\/u1\/_0111_ ), .Y(\u0\/u1\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1413_ ( .A1(\u0\/u1\/_0032_ ), .A2(\u0\/u1\/_0113_ ), .B1(\u0\/u1\/_0636_ ), .C1(\u0\/u1\/_0400_ ), .Y(\u0\/u1\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1414_ ( .A1(\u0\/u1\/_0731_ ), .A2(\u0\/u1\/_0293_ ), .A3(\u0\/u1\/_0251_ ), .B1(\u0\/u1\/_0099_ ), .Y(\u0\/u1\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1415_ ( .A(\u0\/u1\/_0189_ ), .B(\u0\/u1\/_0635_ ), .C(\u0\/u1\/_0637_ ), .D(\u0\/u1\/_0638_ ), .X(\u0\/u1\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1416_ ( .A(\u0\/u1\/_0625_ ), .B(\u0\/u1\/_0630_ ), .C(\u0\/u1\/_0633_ ), .D(\u0\/u1\/_0639_ ), .X(\u0\/u1\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1417_ ( .A(\u0\/u1\/_0746_ ), .B(\u0\/u1\/_0738_ ), .X(\u0\/u1\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1418_ ( .A(\u0\/u1\/_0736_ ), .B(\u0\/u1\/_0731_ ), .X(\u0\/u1\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u1/_1419_ ( .A_N(\u0\/u1\/_0643_ ), .B(\u0\/u1\/_0577_ ), .Y(\u0\/u1\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1420_ ( .A1(\u0\/u1\/_0084_ ), .A2(\u0\/u1\/_0739_ ), .B1(\u0\/u1\/_0642_ ), .C1(\u0\/u1\/_0644_ ), .Y(\u0\/u1\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1421_ ( .A1(\u0\/u1\/_0050_ ), .A2(\u0\/u1\/_0543_ ), .B1(\u0\/u1\/_0194_ ), .C1(\u0\/u1\/_0738_ ), .Y(\u0\/u1\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1422_ ( .A(\u0\/u1\/_0646_ ), .B(\u0\/u1\/_0232_ ), .C(\u0\/u1\/_0417_ ), .D(\u0\/u1\/_0578_ ), .X(\u0\/u1\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1423_ ( .A1(\u0\/u1\/_0064_ ), .A2(\u0\/u1\/_0733_ ), .B1(\u0\/u1\/_0727_ ), .Y(\u0\/u1\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1424_ ( .A1(\u0\/u1\/_0193_ ), .A2(\u0\/u1\/_0276_ ), .B1(\u0\/u1\/_0727_ ), .Y(\u0\/u1\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1425_ ( .A(\u0\/u1\/_0645_ ), .B(\u0\/u1\/_0647_ ), .C(\u0\/u1\/_0648_ ), .D(\u0\/u1\/_0649_ ), .X(\u0\/u1\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1426_ ( .A1(\u0\/u1\/_0325_ ), .A2(\u0\/u1\/_0734_ ), .B1(\u0\/u1\/_0038_ ), .C1(\u0\/u1\/_0029_ ), .Y(\u0\/u1\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1427_ ( .A1(\u0\/u1\/_0543_ ), .A2(\u0\/u1\/_0216_ ), .B1(\u0\/u1\/_0412_ ), .C1(\u0\/u1\/_0029_ ), .Y(\u0\/u1\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1428_ ( .A(\u0\/u1\/_0652_ ), .B(\u0\/u1\/_0653_ ), .X(\u0\/u1\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1429_ ( .A1(\u0\/u1\/_0733_ ), .A2(\u0\/u1\/_0748_ ), .A3(\u0\/u1\/_0324_ ), .B1(\u0\/u1\/_0016_ ), .Y(\u0\/u1\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1430_ ( .A1(\u0\/u1\/_0640_ ), .A2(\u0\/u1\/_0193_ ), .A3(\u0\/u1\/_0091_ ), .B1(\u0\/u1\/_0016_ ), .Y(\u0\/u1\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1431_ ( .A1(\u0\/u1\/_0102_ ), .A2(\u0\/u1\/_0301_ ), .B1(\w3\[11\] ), .C1(\u0\/u1\/_0029_ ), .Y(\u0\/u1\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1432_ ( .A(\u0\/u1\/_0654_ ), .B(\u0\/u1\/_0655_ ), .C(\u0\/u1\/_0656_ ), .D(\u0\/u1\/_0657_ ), .X(\u0\/u1\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1433_ ( .A1(\u0\/u1\/_0118_ ), .A2(\u0\/u1\/_0050_ ), .B1(\u0\/u1\/_0038_ ), .C1(\u0\/u1\/_0478_ ), .Y(\u0\/u1\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u1/_1434_ ( .A_N(\u0\/u1\/_0250_ ), .B(\u0\/u1\/_0465_ ), .C(\u0\/u1\/_0659_ ), .X(\u0\/u1\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1435_ ( .A1(\u0\/u1\/_0683_ ), .A2(\u0\/u1\/_0324_ ), .B1(\u0\/u1\/_0255_ ), .Y(\u0\/u1\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1436_ ( .A1(\u0\/u1\/_0032_ ), .A2(\u0\/u1\/_0193_ ), .A3(\u0\/u1\/_0047_ ), .B1(\u0\/u1\/_0255_ ), .Y(\u0\/u1\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1437_ ( .A1(\u0\/u1\/_0144_ ), .A2(\u0\/u1\/_0586_ ), .A3(\u0\/u1\/_0047_ ), .B1(\u0\/u1\/_0218_ ), .Y(\u0\/u1\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1438_ ( .A(\u0\/u1\/_0660_ ), .B(\u0\/u1\/_0661_ ), .C(\u0\/u1\/_0663_ ), .D(\u0\/u1\/_0664_ ), .X(\u0\/u1\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1439_ ( .A1(\u0\/u1\/_0091_ ), .A2(\u0\/u1\/_0276_ ), .B1(\u0\/u1\/_0060_ ), .Y(\u0\/u1\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1440_ ( .A1(\u0\/u1\/_0144_ ), .A2(\u0\/u1\/_0608_ ), .B1(\u0\/u1\/_0056_ ), .Y(\u0\/u1\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1441_ ( .A1(\u0\/u1\/_0412_ ), .A2(\u0\/u1\/_0038_ ), .B1(\u0\/u1\/_0102_ ), .C1(\u0\/u1\/_0060_ ), .Y(\u0\/u1\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1442_ ( .A1(\w3\[9\] ), .A2(\u0\/u1\/_0734_ ), .B1(\u0\/u1\/_0109_ ), .C1(\u0\/u1\/_0056_ ), .Y(\u0\/u1\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1443_ ( .A(\u0\/u1\/_0666_ ), .B(\u0\/u1\/_0667_ ), .C(\u0\/u1\/_0668_ ), .D(\u0\/u1\/_0669_ ), .X(\u0\/u1\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1444_ ( .A(\u0\/u1\/_0650_ ), .B(\u0\/u1\/_0658_ ), .C(\u0\/u1\/_0665_ ), .D(\u0\/u1\/_0670_ ), .X(\u0\/u1\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u1/_1445_ ( .A(\u0\/u1\/_0641_ ), .B(\u0\/u1\/_0174_ ), .C(\u0\/u1\/_0671_ ), .Y(\u0\/u1\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u1/_1446_ ( .A(\u0\/u1\/_0049_ ), .B(\u0\/u1\/_0618_ ), .C_N(\u0\/u1\/_0052_ ), .Y(\u0\/u1\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \u0/u1/_1447_ ( .A(\u0\/u1\/_0239_ ), .Y(\u0\/u1\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1448_ ( .A(\u0\/u1\/_0705_ ), .B(\u0\/u1\/_0032_ ), .Y(\u0\/u1\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1449_ ( .A1(\u0\/u1\/_0054_ ), .A2(\u0\/u1\/_0731_ ), .B1(\u0\/u1\/_0035_ ), .B2(\u0\/u1\/_0705_ ), .Y(\u0\/u1\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1450_ ( .A1(\u0\/u1\/_0304_ ), .A2(\u0\/u1\/_0731_ ), .B1(\u0\/u1\/_0047_ ), .B2(\u0\/u1\/_0750_ ), .Y(\u0\/u1\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1451_ ( .A(\u0\/u1\/_0674_ ), .B(\u0\/u1\/_0675_ ), .C(\u0\/u1\/_0676_ ), .D(\u0\/u1\/_0677_ ), .X(\u0\/u1\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u1/_1452_ ( .A_N(\u0\/u1\/_0584_ ), .B(\u0\/u1\/_0283_ ), .X(\u0\/u1\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1453_ ( .A(\u0\/u1\/_0673_ ), .B(\u0\/u1\/_0678_ ), .C(\u0\/u1\/_0679_ ), .D(\u0\/u1\/_0508_ ), .X(\u0\/u1\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1454_ ( .A1(\u0\/u1\/_0016_ ), .A2(\u0\/u1\/_0733_ ), .B1(\u0\/u1\/_0355_ ), .B2(\u0\/u1\/_0092_ ), .Y(\u0\/u1\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1455_ ( .A(\u0\/u1\/_0681_ ), .B(\u0\/u1\/_0034_ ), .X(\u0\/u1\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u1/_1456_ ( .A1(\u0\/u1\/_0330_ ), .A2(\u0\/u1\/_0139_ ), .B1(\u0\/u1\/_0324_ ), .B2(\u0\/u1\/_0089_ ), .X(\u0\/u1\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1457_ ( .A1(\u0\/u1\/_0146_ ), .A2(\u0\/u1\/_0147_ ), .B1(\u0\/u1\/_0133_ ), .C1(\u0\/u1\/_0684_ ), .Y(\u0\/u1\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1458_ ( .A(\u0\/u1\/_0113_ ), .B(\u0\/u1\/_0251_ ), .Y(\u0\/u1\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u1/_1459_ ( .A_N(\u0\/u1\/_0463_ ), .B(\u0\/u1\/_0686_ ), .C(\u0\/u1\/_0383_ ), .D(\u0\/u1\/_0464_ ), .X(\u0\/u1\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1460_ ( .A1(\u0\/u1\/_0051_ ), .A2(\u0\/u1\/_0293_ ), .B1(\u0\/u1\/_0084_ ), .B2(\u0\/u1\/_0705_ ), .Y(\u0\/u1\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1461_ ( .A1(\u0\/u1\/_0017_ ), .A2(\u0\/u1\/_0072_ ), .B1(\u0\/u1\/_0456_ ), .B2(\u0\/u1\/_0078_ ), .Y(\u0\/u1\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1462_ ( .A(\u0\/u1\/_0687_ ), .B(\u0\/u1\/_0236_ ), .C(\u0\/u1\/_0688_ ), .D(\u0\/u1\/_0689_ ), .X(\u0\/u1\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1463_ ( .A(\u0\/u1\/_0680_ ), .B(\u0\/u1\/_0682_ ), .C(\u0\/u1\/_0685_ ), .D(\u0\/u1\/_0690_ ), .X(\u0\/u1\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u1/_1464_ ( .A1(\u0\/u1\/_0532_ ), .A2(\u0\/u1\/_0380_ ), .B1(\u0\/u1\/_0102_ ), .C1(\u0\/u1\/_0355_ ), .X(\u0\/u1\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u1/_1465_ ( .A(\u0\/u1\/_0692_ ), .B(\u0\/u1\/_0338_ ), .C(\u0\/u1\/_0644_ ), .Y(\u0\/u1\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1466_ ( .A(\u0\/u1\/_0016_ ), .B(\u0\/u1\/_0020_ ), .Y(\u0\/u1\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1467_ ( .A1(\u0\/u1\/_0032_ ), .A2(\u0\/u1\/_0137_ ), .B1(\u0\/u1\/_0279_ ), .B2(\u0\/u1\/_0094_ ), .Y(\u0\/u1\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1468_ ( .A1(\u0\/u1\/_0575_ ), .A2(\u0\/u1\/_0153_ ), .B1(\u0\/u1\/_0161_ ), .B2(\u0\/u1\/_0293_ ), .Y(\u0\/u1\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1469_ ( .A(\u0\/u1\/_0259_ ), .B(\u0\/u1\/_0695_ ), .C(\u0\/u1\/_0696_ ), .D(\u0\/u1\/_0697_ ), .X(\u0\/u1\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u1/_1470_ ( .A1(\u0\/u1\/_0255_ ), .A2(\u0\/u1\/_0640_ ), .B1(\u0\/u1\/_0016_ ), .B2(\u0\/u1\/_0193_ ), .X(\u0\/u1\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1471_ ( .A1(\u0\/u1\/_0060_ ), .A2(\u0\/u1\/_0176_ ), .B1(\u0\/u1\/_0699_ ), .C1(\u0\/u1\/_0177_ ), .Y(\u0\/u1\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1472_ ( .A1(\u0\/u1\/_0091_ ), .A2(\u0\/u1\/_0218_ ), .B1(\u0\/u1\/_0092_ ), .B2(\u0\/u1\/_0705_ ), .Y(\u0\/u1\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u1/_1473_ ( .A1(\u0\/u1\/_0705_ ), .A2(\u0\/u1\/_0683_ ), .B1(\u0\/u1\/_0093_ ), .B2(\u0\/u1\/_0114_ ), .Y(\u0\/u1\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u1/_1474_ ( .A1(\u0\/u1\/_0683_ ), .A2(\u0\/u1\/_0084_ ), .B1(\u0\/u1\/_0094_ ), .Y(\u0\/u1\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u1/_1475_ ( .A1(\u0\/u1\/_0543_ ), .A2(\u0\/u1\/_0216_ ), .B1(\u0\/u1\/_0038_ ), .C1(\u0\/u1\/_0056_ ), .Y(\u0\/u1\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1476_ ( .A(\u0\/u1\/_0701_ ), .B(\u0\/u1\/_0702_ ), .C(\u0\/u1\/_0703_ ), .D(\u0\/u1\/_0704_ ), .X(\u0\/u1\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1477_ ( .A(\u0\/u1\/_0693_ ), .B(\u0\/u1\/_0698_ ), .C(\u0\/u1\/_0700_ ), .D(\u0\/u1\/_0706_ ), .X(\u0\/u1\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u1/_1478_ ( .A1(\u0\/u1\/_0113_ ), .A2(\u0\/u1\/_0640_ ), .B1(\u0\/u1\/_0099_ ), .B2(\u0\/u1\/_0058_ ), .X(\u0\/u1\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u1/_1479_ ( .A(\u0\/u1\/_0407_ ), .B(\u0\/u1\/_0708_ ), .C(\u0\/u1\/_0529_ ), .Y(\u0\/u1\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1480_ ( .A(\u0\/u1\/_0568_ ), .B(\u0\/u1\/_0175_ ), .Y(\u0\/u1\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u1/_1481_ ( .A1(\u0\/u1\/_0029_ ), .A2(\u0\/u1\/_0114_ ), .A3(\u0\/u1\/_0051_ ), .B1(\u0\/u1\/_0130_ ), .Y(\u0\/u1\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1482_ ( .A(\u0\/u1\/_0709_ ), .B(\u0\/u1\/_0550_ ), .C(\u0\/u1\/_0710_ ), .D(\u0\/u1\/_0711_ ), .X(\u0\/u1\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u1/_1483_ ( .A1(\u0\/u1\/_0114_ ), .A2(\u0\/u1\/_0064_ ), .B1(\u0\/u1\/_0261_ ), .B2(\u0\/u1\/_0089_ ), .X(\u0\/u1\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1484_ ( .A1(\u0\/u1\/_0355_ ), .A2(\u0\/u1\/_0261_ ), .B1(\u0\/u1\/_0198_ ), .C1(\u0\/u1\/_0713_ ), .Y(\u0\/u1\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1485_ ( .A(\u0\/u1\/_0586_ ), .B(\u0\/u1\/_0478_ ), .Y(\u0\/u1\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u1/_1486_ ( .A_N(\u0\/u1\/_0541_ ), .B(\u0\/u1\/_0267_ ), .C(\u0\/u1\/_0715_ ), .D(\u0\/u1\/_0320_ ), .X(\u0\/u1\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1487_ ( .A(\u0\/u1\/_0586_ ), .B(\u0\/u1\/_0070_ ), .Y(\u0\/u1\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u1/_1488_ ( .A_N(\u0\/u1\/_0211_ ), .B(\u0\/u1\/_0155_ ), .C(\u0\/u1\/_0202_ ), .D(\u0\/u1\/_0718_ ), .X(\u0\/u1\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u1/_1489_ ( .A(\u0\/u1\/_0150_ ), .B(\u0\/u1\/_0216_ ), .C(\u0\/u1\/_0380_ ), .Y(\u0\/u1\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \u0/u1/_1490_ ( .A(\u0\/u1\/_0411_ ), .B(\u0\/u1\/_0720_ ), .X(\u0\/u1\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u1/_1491_ ( .A1(\u0\/u1\/_0017_ ), .A2(\u0\/u1\/_0022_ ), .B1(\u0\/u1\/_0078_ ), .X(\u0\/u1\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u1/_1492_ ( .A1(\u0\/u1\/_0456_ ), .A2(\u0\/u1\/_0738_ ), .B1(\u0\/u1\/_0101_ ), .C1(\u0\/u1\/_0722_ ), .Y(\u0\/u1\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1493_ ( .A(\u0\/u1\/_0717_ ), .B(\u0\/u1\/_0719_ ), .C(\u0\/u1\/_0721_ ), .D(\u0\/u1\/_0723_ ), .X(\u0\/u1\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u1/_1494_ ( .A(\u0\/u1\/_0739_ ), .B(\u0\/u1\/_0193_ ), .Y(\u0\/u1\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1495_ ( .A(\u0\/u1\/_0344_ ), .B(\u0\/u1\/_0184_ ), .C(\u0\/u1\/_0449_ ), .D(\u0\/u1\/_0725_ ), .X(\u0\/u1\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \u0/u1/_1496_ ( .A(\u0\/u1\/_0712_ ), .B(\u0\/u1\/_0714_ ), .C(\u0\/u1\/_0724_ ), .D(\u0\/u1\/_0726_ ), .X(\u0\/u1\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u1/_1497_ ( .A(\u0\/u1\/_0691_ ), .B(\u0\/u1\/_0707_ ), .C(\u0\/u1\/_0728_ ), .Y(\u0\/u1\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u2/_0753_ ( .A(\w3\[2\] ), .B_N(\w3\[3\] ), .Y(\u0\/u2\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0755_ ( .A(\w3\[1\] ), .B(\w3\[0\] ), .X(\u0\/u2\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0756_ ( .A(\u0\/u2\/_0096_ ), .B(\u0\/u2\/_0118_ ), .X(\u0\/u2\/_0129_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0757_ ( .A(\w3\[7\] ), .B(\w3\[6\] ), .X(\u0\/u2\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_0758_ ( .A(\w3\[4\] ), .B(\w3\[5\] ), .Y(\u0\/u2\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0759_ ( .A(\u0\/u2\/_0140_ ), .B(\u0\/u2\/_0151_ ), .X(\u0\/u2\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0761_ ( .A(\u0\/u2\/_0129_ ), .B(\u0\/u2\/_0162_ ), .X(\u0\/u2\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0762_ ( .A(\u0\/u2\/_0096_ ), .X(\u0\/u2\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u2/_0763_ ( .A(\w3\[1\] ), .B_N(\w3\[0\] ), .Y(\u0\/u2\/_0205_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0764_ ( .A(\u0\/u2\/_0205_ ), .X(\u0\/u2\/_0216_ ) );
sky130_fd_sc_hd__and3_1 \u0/u2/_0765_ ( .A(\u0\/u2\/_0162_ ), .B(\u0\/u2\/_0194_ ), .C(\u0\/u2\/_0216_ ), .X(\u0\/u2\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \u0/u2/_0766_ ( .A(\u0\/u2\/_0183_ ), .SLEEP(\u0\/u2\/_0227_ ), .X(\u0\/u2\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u2/_0767_ ( .A(\w3\[0\] ), .B_N(\w3\[1\] ), .Y(\u0\/u2\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_0768_ ( .A(\w3\[2\] ), .B(\w3\[3\] ), .Y(\u0\/u2\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0769_ ( .A(\u0\/u2\/_0249_ ), .B(\u0\/u2\/_0260_ ), .X(\u0\/u2\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0771_ ( .A(\u0\/u2\/_0271_ ), .X(\u0\/u2\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0772_ ( .A(\u0\/u2\/_0162_ ), .X(\u0\/u2\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_0773_ ( .A(\u0\/u2\/_0293_ ), .B(\u0\/u2\/_0304_ ), .Y(\u0\/u2\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \u0/u2/_0774_ ( .A(\w3\[1\] ), .Y(\u0\/u2\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \u0/u2/_0776_ ( .A(\w3\[0\] ), .Y(\u0\/u2\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0777_ ( .A(\w3\[2\] ), .B(\w3\[3\] ), .X(\u0\/u2\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0779_ ( .A(\u0\/u2\/_0358_ ), .X(\u0\/u2\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_0780_ ( .A1(\u0\/u2\/_0325_ ), .A2(\u0\/u2\/_0347_ ), .B1(\u0\/u2\/_0380_ ), .C1(\u0\/u2\/_0304_ ), .Y(\u0\/u2\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u2/_0781_ ( .A_N(\u0\/u2\/_0238_ ), .B(\u0\/u2\/_0314_ ), .C(\u0\/u2\/_0391_ ), .X(\u0\/u2\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u2/_0782_ ( .A(\w3\[3\] ), .B_N(\w3\[2\] ), .Y(\u0\/u2\/_0412_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0783_ ( .A(\u0\/u2\/_0412_ ), .X(\u0\/u2\/_0423_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0784_ ( .A(\u0\/u2\/_0423_ ), .B(\u0\/u2\/_0205_ ), .X(\u0\/u2\/_0434_ ) );
sky130_fd_sc_hd__buf_2 \u0/u2/_0786_ ( .A(\u0\/u2\/_0434_ ), .X(\u0\/u2\/_0456_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u2/_0787_ ( .A(\w3\[5\] ), .B_N(\w3\[4\] ), .Y(\u0\/u2\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0788_ ( .A(\u0\/u2\/_0467_ ), .B(\u0\/u2\/_0140_ ), .X(\u0\/u2\/_0478_ ) );
sky130_fd_sc_hd__buf_2 \u0/u2/_0790_ ( .A(\u0\/u2\/_0478_ ), .X(\u0\/u2\/_0499_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_0791_ ( .A(\u0\/u2\/_0456_ ), .B(\u0\/u2\/_0499_ ), .Y(\u0\/u2\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_0792_ ( .A(\u0\/u2\/_0478_ ), .B(\u0\/u2\/_0271_ ), .Y(\u0\/u2\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0793_ ( .A(\u0\/u2\/_0194_ ), .X(\u0\/u2\/_0532_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0794_ ( .A(\u0\/u2\/_0249_ ), .X(\u0\/u2\/_0543_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0795_ ( .A(\u0\/u2\/_0543_ ), .B(\u0\/u2\/_0358_ ), .X(\u0\/u2\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0797_ ( .A(\u0\/u2\/_0554_ ), .X(\u0\/u2\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0798_ ( .A(\u0\/u2\/_0216_ ), .B(\u0\/u2\/_0358_ ), .X(\u0\/u2\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0800_ ( .A(\u0\/u2\/_0586_ ), .X(\u0\/u2\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_0801_ ( .A1(\u0\/u2\/_0532_ ), .A2(\u0\/u2\/_0575_ ), .A3(\u0\/u2\/_0608_ ), .B1(\u0\/u2\/_0499_ ), .Y(\u0\/u2\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_0802_ ( .A(\u0\/u2\/_0401_ ), .B(\u0\/u2\/_0510_ ), .C(\u0\/u2\/_0521_ ), .D(\u0\/u2\/_0619_ ), .X(\u0\/u2\/_0629_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0803_ ( .A(\u0\/u2\/_0358_ ), .B(\w3\[1\] ), .X(\u0\/u2\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0805_ ( .A(\u0\/u2\/_0205_ ), .B(\u0\/u2\/_0260_ ), .X(\u0\/u2\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0807_ ( .A(\u0\/u2\/_0662_ ), .X(\u0\/u2\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u2/_0808_ ( .A(\w3\[6\] ), .B_N(\w3\[7\] ), .Y(\u0\/u2\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0809_ ( .A(\u0\/u2\/_0467_ ), .B(\u0\/u2\/_0694_ ), .X(\u0\/u2\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0811_ ( .A(\u0\/u2\/_0705_ ), .X(\u0\/u2\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_0812_ ( .A1(\u0\/u2\/_0640_ ), .A2(\u0\/u2\/_0293_ ), .A3(\u0\/u2\/_0683_ ), .B1(\u0\/u2\/_0727_ ), .Y(\u0\/u2\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_0813_ ( .A(\w3\[1\] ), .B(\w3\[0\] ), .Y(\u0\/u2\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0814_ ( .A(\u0\/u2\/_0730_ ), .B(\u0\/u2\/_0260_ ), .X(\u0\/u2\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0816_ ( .A(\u0\/u2\/_0731_ ), .X(\u0\/u2\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0817_ ( .A(\w3\[0\] ), .X(\u0\/u2\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u2/_0818_ ( .A1(\u0\/u2\/_0325_ ), .A2(\u0\/u2\/_0734_ ), .B1(\u0\/u2\/_0423_ ), .X(\u0\/u2\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0819_ ( .A(\u0\/u2\/_0694_ ), .B(\u0\/u2\/_0151_ ), .X(\u0\/u2\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0821_ ( .A(\u0\/u2\/_0736_ ), .X(\u0\/u2\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0822_ ( .A(\u0\/u2\/_0738_ ), .X(\u0\/u2\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_0823_ ( .A1(\u0\/u2\/_0733_ ), .A2(\u0\/u2\/_0735_ ), .A3(\u0\/u2\/_0293_ ), .B1(\u0\/u2\/_0739_ ), .Y(\u0\/u2\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u2/_0824_ ( .A(\u0\/u2\/_0730_ ), .B_N(\u0\/u2\/_0358_ ), .Y(\u0\/u2\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_0825_ ( .A(\u0\/u2\/_0741_ ), .B(\u0\/u2\/_0739_ ), .Y(\u0\/u2\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_0827_ ( .A1(\u0\/u2\/_0118_ ), .A2(\u0\/u2\/_0216_ ), .B1(\u0\/u2\/_0532_ ), .C1(\u0\/u2\/_0739_ ), .Y(\u0\/u2\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_0828_ ( .A(\u0\/u2\/_0729_ ), .B(\u0\/u2\/_0740_ ), .C(\u0\/u2\/_0742_ ), .D(\u0\/u2\/_0744_ ), .X(\u0\/u2\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0829_ ( .A(\u0\/u2\/_0423_ ), .B(\u0\/u2\/_0730_ ), .X(\u0\/u2\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0831_ ( .A(\u0\/u2\/_0746_ ), .X(\u0\/u2\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u2/_0832_ ( .A(\w3\[4\] ), .B_N(\w3\[5\] ), .Y(\u0\/u2\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0833_ ( .A(\u0\/u2\/_0749_ ), .B(\u0\/u2\/_0694_ ), .X(\u0\/u2\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0835_ ( .A(\u0\/u2\/_0750_ ), .X(\u0\/u2\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0836_ ( .A(\u0\/u2\/_0752_ ), .X(\u0\/u2\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0837_ ( .A(\u0\/u2\/_0118_ ), .B(\u0\/u2\/_0358_ ), .X(\u0\/u2\/_0017_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0839_ ( .A(\u0\/u2\/_0752_ ), .B(\u0\/u2\/_0017_ ), .X(\u0\/u2\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0840_ ( .A(\u0\/u2\/_0358_ ), .B(\u0\/u2\/_0325_ ), .X(\u0\/u2\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0842_ ( .A(\u0\/u2\/_0096_ ), .B(\u0\/u2\/_0205_ ), .X(\u0\/u2\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u2/_0844_ ( .A1(\u0\/u2\/_0020_ ), .A2(\u0\/u2\/_0022_ ), .B1(\u0\/u2\/_0752_ ), .X(\u0\/u2\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_0845_ ( .A1(\u0\/u2\/_0748_ ), .A2(\u0\/u2\/_0016_ ), .B1(\u0\/u2\/_0019_ ), .C1(\u0\/u2\/_0024_ ), .Y(\u0\/u2\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0846_ ( .A(\w3\[4\] ), .B(\w3\[5\] ), .X(\u0\/u2\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0847_ ( .A(\u0\/u2\/_0694_ ), .B(\u0\/u2\/_0026_ ), .X(\u0\/u2\/_0027_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0850_ ( .A(\u0\/u2\/_0358_ ), .B(\u0\/u2\/_0730_ ), .X(\u0\/u2\/_0030_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0852_ ( .A(\u0\/u2\/_0030_ ), .X(\u0\/u2\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_0853_ ( .A(\u0\/u2\/_0247_ ), .B(\u0\/u2\/_0032_ ), .Y(\u0\/u2\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_0854_ ( .A(\u0\/u2\/_0247_ ), .B(\u0\/u2\/_0735_ ), .Y(\u0\/u2\/_0034_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0855_ ( .A(\u0\/u2\/_0118_ ), .B(\u0\/u2\/_0260_ ), .X(\u0\/u2\/_0035_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0857_ ( .A(\u0\/u2\/_0027_ ), .B(\u0\/u2\/_0035_ ), .X(\u0\/u2\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0858_ ( .A(\u0\/u2\/_0260_ ), .X(\u0\/u2\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_0859_ ( .A(\u0\/u2\/_0038_ ), .B(\u0\/u2\/_0347_ ), .Y(\u0\/u2\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u2/_0860_ ( .A_N(\u0\/u2\/_0039_ ), .B(\u0\/u2\/_0027_ ), .X(\u0\/u2\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_0861_ ( .A(\u0\/u2\/_0037_ ), .B(\u0\/u2\/_0040_ ), .Y(\u0\/u2\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_0862_ ( .A(\u0\/u2\/_0025_ ), .B(\u0\/u2\/_0033_ ), .C(\u0\/u2\/_0034_ ), .D(\u0\/u2\/_0041_ ), .X(\u0\/u2\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0863_ ( .A(\u0\/u2\/_0749_ ), .B(\u0\/u2\/_0140_ ), .X(\u0\/u2\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \u0/u2/_0865_ ( .A(\w3\[0\] ), .B(\w3\[2\] ), .C(\w3\[3\] ), .X(\u0\/u2\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0866_ ( .A(\u0\/u2\/_0043_ ), .B(\u0\/u2\/_0045_ ), .X(\u0\/u2\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0867_ ( .A(\u0\/u2\/_0096_ ), .B(\u0\/u2\/_0543_ ), .X(\u0\/u2\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0869_ ( .A(\u0\/u2\/_0047_ ), .B(\u0\/u2\/_0043_ ), .X(\u0\/u2\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0870_ ( .A(\u0\/u2\/_0730_ ), .X(\u0\/u2\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0871_ ( .A(\u0\/u2\/_0043_ ), .X(\u0\/u2\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_0872_ ( .A1(\u0\/u2\/_0118_ ), .A2(\u0\/u2\/_0050_ ), .B1(\u0\/u2\/_0194_ ), .C1(\u0\/u2\/_0051_ ), .Y(\u0\/u2\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u2/_0873_ ( .A(\u0\/u2\/_0046_ ), .B(\u0\/u2\/_0049_ ), .C_N(\u0\/u2\/_0052_ ), .Y(\u0\/u2\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0874_ ( .A(\u0\/u2\/_0026_ ), .B(\u0\/u2\/_0140_ ), .X(\u0\/u2\/_0054_ ) );
sky130_fd_sc_hd__buf_2 \u0/u2/_0876_ ( .A(\u0\/u2\/_0054_ ), .X(\u0\/u2\/_0056_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_0877_ ( .A1(\u0\/u2\/_0532_ ), .A2(\u0\/u2\/_0575_ ), .B1(\u0\/u2\/_0056_ ), .Y(\u0\/u2\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0878_ ( .A(\u0\/u2\/_0423_ ), .B(\u0\/u2\/_0325_ ), .X(\u0\/u2\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0880_ ( .A(\u0\/u2\/_0051_ ), .X(\u0\/u2\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_0881_ ( .A1(\u0\/u2\/_0731_ ), .A2(\u0\/u2\/_0035_ ), .A3(\u0\/u2\/_0058_ ), .B1(\u0\/u2\/_0060_ ), .Y(\u0\/u2\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0882_ ( .A(\u0\/u2\/_0260_ ), .B(\w3\[1\] ), .X(\u0\/u2\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0884_ ( .A(\u0\/u2\/_0062_ ), .X(\u0\/u2\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_0885_ ( .A1(\u0\/u2\/_0064_ ), .A2(\u0\/u2\/_0748_ ), .A3(\u0\/u2\/_0683_ ), .B1(\u0\/u2\/_0056_ ), .Y(\u0\/u2\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_0886_ ( .A(\u0\/u2\/_0053_ ), .B(\u0\/u2\/_0057_ ), .C(\u0\/u2\/_0061_ ), .D(\u0\/u2\/_0065_ ), .X(\u0\/u2\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_0887_ ( .A(\u0\/u2\/_0629_ ), .B(\u0\/u2\/_0745_ ), .C(\u0\/u2\/_0042_ ), .D(\u0\/u2\/_0066_ ), .X(\u0\/u2\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u2/_0889_ ( .A(\w3\[7\] ), .B_N(\w3\[6\] ), .Y(\u0\/u2\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0890_ ( .A(\u0\/u2\/_0069_ ), .B(\u0\/u2\/_0151_ ), .X(\u0\/u2\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0892_ ( .A(\u0\/u2\/_0070_ ), .X(\u0\/u2\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_0893_ ( .A1(\u0\/u2\/_0129_ ), .A2(\u0\/u2\/_0586_ ), .B1(\u0\/u2\/_0072_ ), .Y(\u0\/u2\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_0894_ ( .A1(\u0\/u2\/_0380_ ), .A2(\u0\/u2\/_0347_ ), .B1(\u0\/u2\/_0194_ ), .B2(\u0\/u2\/_0216_ ), .Y(\u0\/u2\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u2/_0895_ ( .A(\u0\/u2\/_0074_ ), .B_N(\u0\/u2\/_0070_ ), .Y(\u0\/u2\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u2/_0896_ ( .A(\u0\/u2\/_0073_ ), .SLEEP(\u0\/u2\/_0075_ ), .X(\u0\/u2\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0897_ ( .A(\u0\/u2\/_0467_ ), .B(\u0\/u2\/_0069_ ), .X(\u0\/u2\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0898_ ( .A(\u0\/u2\/_0077_ ), .X(\u0\/u2\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0899_ ( .A(\u0\/u2\/_0412_ ), .B(\u0\/u2\/_0118_ ), .X(\u0\/u2\/_0079_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0901_ ( .A(\u0\/u2\/_0078_ ), .B(\u0\/u2\/_0079_ ), .X(\u0\/u2\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0902_ ( .A(\u0\/u2\/_0412_ ), .B(\u0\/u2\/_0249_ ), .X(\u0\/u2\/_0082_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0905_ ( .A(\u0\/u2\/_0280_ ), .B(\u0\/u2\/_0078_ ), .X(\u0\/u2\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u2/_0906_ ( .A1(\w3\[0\] ), .A2(\u0\/u2\/_0325_ ), .B1(\u0\/u2\/_0260_ ), .Y(\u0\/u2\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u2/_0907_ ( .A_N(\u0\/u2\/_0086_ ), .B(\u0\/u2\/_0078_ ), .X(\u0\/u2\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u2/_0908_ ( .A(\u0\/u2\/_0081_ ), .B(\u0\/u2\/_0085_ ), .C(\u0\/u2\/_0087_ ), .Y(\u0\/u2\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0909_ ( .A(\u0\/u2\/_0072_ ), .X(\u0\/u2\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_0910_ ( .A1(\u0\/u2\/_0733_ ), .A2(\u0\/u2\/_0748_ ), .A3(\u0\/u2\/_0683_ ), .B1(\u0\/u2\/_0089_ ), .Y(\u0\/u2\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0911_ ( .A(\u0\/u2\/_0129_ ), .X(\u0\/u2\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0912_ ( .A(\u0\/u2\/_0017_ ), .X(\u0\/u2\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0913_ ( .A(\u0\/u2\/_0022_ ), .X(\u0\/u2\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0914_ ( .A(\u0\/u2\/_0078_ ), .X(\u0\/u2\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_0915_ ( .A1(\u0\/u2\/_0091_ ), .A2(\u0\/u2\/_0092_ ), .A3(\u0\/u2\/_0093_ ), .B1(\u0\/u2\/_0094_ ), .Y(\u0\/u2\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_0916_ ( .A(\u0\/u2\/_0076_ ), .B(\u0\/u2\/_0088_ ), .C(\u0\/u2\/_0090_ ), .D(\u0\/u2\/_0095_ ), .X(\u0\/u2\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0917_ ( .A(\u0\/u2\/_0069_ ), .B(\u0\/u2\/_0026_ ), .X(\u0\/u2\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \u0/u2/_0918_ ( .A(\u0\/u2\/_0098_ ), .X(\u0\/u2\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0919_ ( .A(\u0\/u2\/_0434_ ), .B(\u0\/u2\/_0099_ ), .X(\u0\/u2\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0920_ ( .A(\u0\/u2\/_0079_ ), .B(\u0\/u2\/_0098_ ), .X(\u0\/u2\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0921_ ( .A(\u0\/u2\/_0325_ ), .X(\u0\/u2\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_0922_ ( .A1(\u0\/u2\/_0102_ ), .A2(\u0\/u2\/_0734_ ), .B1(\u0\/u2\/_0038_ ), .C1(\u0\/u2\/_0099_ ), .Y(\u0\/u2\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u2/_0923_ ( .A(\u0\/u2\/_0100_ ), .B(\u0\/u2\/_0101_ ), .C_N(\u0\/u2\/_0103_ ), .Y(\u0\/u2\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_0924_ ( .A1(\u0\/u2\/_0554_ ), .A2(\u0\/u2\/_0586_ ), .B1(\u0\/u2\/_0099_ ), .Y(\u0\/u2\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_0925_ ( .A(\u0\/u2\/_0129_ ), .B(\u0\/u2\/_0099_ ), .Y(\u0\/u2\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0926_ ( .A(\u0\/u2\/_0105_ ), .B(\u0\/u2\/_0106_ ), .X(\u0\/u2\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0927_ ( .A(\u0\/u2\/_0423_ ), .X(\u0\/u2\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0928_ ( .A(\u0\/u2\/_0260_ ), .B(\w3\[0\] ), .X(\u0\/u2\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0929_ ( .A(\u0\/u2\/_0069_ ), .B(\u0\/u2\/_0749_ ), .X(\u0\/u2\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0931_ ( .A(\u0\/u2\/_0111_ ), .X(\u0\/u2\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0932_ ( .A(\u0\/u2\/_0113_ ), .X(\u0\/u2\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_0933_ ( .A1(\u0\/u2\/_0109_ ), .A2(\u0\/u2\/_0110_ ), .B1(\u0\/u2\/_0114_ ), .Y(\u0\/u2\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_0934_ ( .A(\u0\/u2\/_0022_ ), .Y(\u0\/u2\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_0935_ ( .A(\u0\/u2\/_0554_ ), .Y(\u0\/u2\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u2/_0936_ ( .A1(\u0\/u2\/_0050_ ), .A2(\u0\/u2\/_0118_ ), .B1(\u0\/u2\/_0194_ ), .Y(\u0\/u2\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_0937_ ( .A(\u0\/u2\/_0113_ ), .Y(\u0\/u2\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \u0/u2/_0938_ ( .A1(\u0\/u2\/_0116_ ), .A2(\u0\/u2\/_0117_ ), .A3(\u0\/u2\/_0119_ ), .B1(\u0\/u2\/_0120_ ), .X(\u0\/u2\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_0939_ ( .A(\u0\/u2\/_0104_ ), .B(\u0\/u2\/_0108_ ), .C(\u0\/u2\/_0115_ ), .D(\u0\/u2\/_0121_ ), .X(\u0\/u2\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_0940_ ( .A(\w3\[7\] ), .B(\w3\[6\] ), .Y(\u0\/u2\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0941_ ( .A(\u0\/u2\/_0749_ ), .B(\u0\/u2\/_0123_ ), .X(\u0\/u2\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0943_ ( .A(\u0\/u2\/_0082_ ), .B(\u0\/u2\/_0124_ ), .X(\u0\/u2\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_0944_ ( .A(\u0\/u2\/_0271_ ), .B(\u0\/u2\/_0124_ ), .Y(\u0\/u2\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0945_ ( .A(\u0\/u2\/_0124_ ), .X(\u0\/u2\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0946_ ( .A(\u0\/u2\/_0260_ ), .B(\u0\/u2\/_0325_ ), .X(\u0\/u2\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_0948_ ( .A(\u0\/u2\/_0128_ ), .B(\u0\/u2\/_0130_ ), .Y(\u0\/u2\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_0949_ ( .A(\u0\/u2\/_0127_ ), .B(\u0\/u2\/_0132_ ), .Y(\u0\/u2\/_0133_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_0951_ ( .A(\u0\/u2\/_0456_ ), .B(\u0\/u2\/_0128_ ), .Y(\u0\/u2\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u2/_0952_ ( .A(\u0\/u2\/_0126_ ), .B(\u0\/u2\/_0133_ ), .C_N(\u0\/u2\/_0135_ ), .Y(\u0\/u2\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0953_ ( .A(\u0\/u2\/_0026_ ), .B(\u0\/u2\/_0123_ ), .X(\u0\/u2\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0955_ ( .A(\u0\/u2\/_0137_ ), .X(\u0\/u2\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_0956_ ( .A1(\u0\/u2\/_0110_ ), .A2(\u0\/u2\/_0293_ ), .A3(\u0\/u2\/_0280_ ), .B1(\u0\/u2\/_0139_ ), .Y(\u0\/u2\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0957_ ( .A(\u0\/u2\/_0096_ ), .B(\u0\/u2\/_0730_ ), .X(\u0\/u2\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0959_ ( .A(\u0\/u2\/_0142_ ), .X(\u0\/u2\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_0960_ ( .A1(\u0\/u2\/_0020_ ), .A2(\u0\/u2\/_0144_ ), .A3(\u0\/u2\/_0017_ ), .B1(\u0\/u2\/_0139_ ), .Y(\u0\/u2\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u2/_0961_ ( .A(\w3\[2\] ), .B(\u0\/u2\/_0050_ ), .C_N(\w3\[3\] ), .Y(\u0\/u2\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0962_ ( .A(\u0\/u2\/_0128_ ), .X(\u0\/u2\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_0963_ ( .A1(\u0\/u2\/_0146_ ), .A2(\u0\/u2\/_0032_ ), .A3(\u0\/u2\/_0640_ ), .B1(\u0\/u2\/_0147_ ), .Y(\u0\/u2\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_0964_ ( .A(\u0\/u2\/_0136_ ), .B(\u0\/u2\/_0141_ ), .C(\u0\/u2\/_0145_ ), .D(\u0\/u2\/_0148_ ), .X(\u0\/u2\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0965_ ( .A(\u0\/u2\/_0123_ ), .B(\u0\/u2\/_0151_ ), .X(\u0\/u2\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0967_ ( .A(\u0\/u2\/_0150_ ), .X(\u0\/u2\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0968_ ( .A(\u0\/u2\/_0150_ ), .B(\u0\/u2\/_0062_ ), .X(\u0\/u2\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_0969_ ( .A(\u0\/u2\/_0079_ ), .B(\u0\/u2\/_0150_ ), .Y(\u0\/u2\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u2/_0970_ ( .A(\u0\/u2\/_0150_ ), .B(\u0\/u2\/_0423_ ), .C(\u0\/u2\/_0543_ ), .Y(\u0\/u2\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_0971_ ( .A(\u0\/u2\/_0155_ ), .B(\u0\/u2\/_0156_ ), .Y(\u0\/u2\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_0972_ ( .A1(\u0\/u2\/_0153_ ), .A2(\u0\/u2\/_0456_ ), .B1(\u0\/u2\/_0154_ ), .C1(\u0\/u2\/_0157_ ), .Y(\u0\/u2\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0973_ ( .A(\u0\/u2\/_0467_ ), .B(\u0\/u2\/_0123_ ), .X(\u0\/u2\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_0975_ ( .A(\u0\/u2\/_0159_ ), .X(\u0\/u2\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u2/_0976_ ( .A_N(\u0\/u2\/_0119_ ), .B(\u0\/u2\/_0161_ ), .X(\u0\/u2\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_0977_ ( .A(\u0\/u2\/_0163_ ), .Y(\u0\/u2\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_0978_ ( .A1(\u0\/u2\/_0146_ ), .A2(\u0\/u2\/_0575_ ), .A3(\u0\/u2\/_0608_ ), .B1(\u0\/u2\/_0153_ ), .Y(\u0\/u2\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_0979_ ( .A1(\u0\/u2\/_0062_ ), .A2(\u0\/u2\/_0280_ ), .A3(\u0\/u2\/_0456_ ), .B1(\u0\/u2\/_0161_ ), .Y(\u0\/u2\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_0980_ ( .A(\u0\/u2\/_0158_ ), .B(\u0\/u2\/_0164_ ), .C(\u0\/u2\/_0165_ ), .D(\u0\/u2\/_0166_ ), .X(\u0\/u2\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_0981_ ( .A(\u0\/u2\/_0097_ ), .B(\u0\/u2\/_0122_ ), .C(\u0\/u2\/_0149_ ), .D(\u0\/u2\/_0167_ ), .X(\u0\/u2\/_0168_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0982_ ( .A(\u0\/u2\/_0662_ ), .B(\u0\/u2\/_0150_ ), .X(\u0\/u2\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_0983_ ( .A(\u0\/u2\/_0154_ ), .B(\u0\/u2\/_0169_ ), .Y(\u0\/u2\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \u0/u2/_0984_ ( .A(\u0\/u2\/_0123_ ), .B(\u0\/u2\/_0151_ ), .C(\u0\/u2\/_0038_ ), .X(\u0\/u2\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0985_ ( .A(\u0\/u2\/_0170_ ), .B(\u0\/u2\/_0171_ ), .X(\u0\/u2\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_0986_ ( .A(\u0\/u2\/_0172_ ), .Y(\u0\/u2\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u2/_0987_ ( .A(\u0\/u2\/_0067_ ), .B(\u0\/u2\/_0168_ ), .C(\u0\/u2\/_0174_ ), .Y(\u0\/u2\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/u2/_0988_ ( .A(\w3\[1\] ), .B(\w3\[0\] ), .Y(\u0\/u2\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_0989_ ( .A(\u0\/u2\/_0175_ ), .B(\u0\/u2\/_0358_ ), .X(\u0\/u2\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0990_ ( .A(\u0\/u2\/_0176_ ), .B(\u0\/u2\/_0478_ ), .X(\u0\/u2\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_0991_ ( .A(\u0\/u2\/_0280_ ), .B(\u0\/u2\/_0113_ ), .Y(\u0\/u2\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0992_ ( .A(\u0\/u2\/_0111_ ), .B(\u0\/u2\/_0062_ ), .X(\u0\/u2\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0993_ ( .A(\u0\/u2\/_0111_ ), .B(\u0\/u2\/_0662_ ), .X(\u0\/u2\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_0994_ ( .A(\u0\/u2\/_0179_ ), .B(\u0\/u2\/_0180_ ), .Y(\u0\/u2\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0995_ ( .A(\u0\/u2\/_0054_ ), .B(\u0\/u2\/_0058_ ), .X(\u0\/u2\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_0996_ ( .A(\u0\/u2\/_0182_ ), .Y(\u0\/u2\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u2/_0997_ ( .A_N(\u0\/u2\/_0177_ ), .B(\u0\/u2\/_0178_ ), .C(\u0\/u2\/_0181_ ), .D(\u0\/u2\/_0184_ ), .X(\u0\/u2\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0998_ ( .A(\u0\/u2\/_0098_ ), .B(\u0\/u2\/_0741_ ), .X(\u0\/u2\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_0999_ ( .A(\u0\/u2\/_0047_ ), .B(\u0\/u2\/_0098_ ), .X(\u0\/u2\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \u0/u2/_1000_ ( .A(\u0\/u2\/_0186_ ), .B(\u0\/u2\/_0187_ ), .X(\u0\/u2\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1001_ ( .A(\u0\/u2\/_0188_ ), .Y(\u0\/u2\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1002_ ( .A(\u0\/u2\/_0738_ ), .B(\u0\/u2\/_0735_ ), .X(\u0\/u2\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1003_ ( .A(\u0\/u2\/_0271_ ), .B(\u0\/u2\/_0736_ ), .X(\u0\/u2\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_1004_ ( .A(\u0\/u2\/_0190_ ), .B(\u0\/u2\/_0191_ ), .Y(\u0\/u2\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_1005_ ( .A(\u0\/u2\/_0096_ ), .B(\u0\/u2\/_0325_ ), .X(\u0\/u2\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1006_ ( .A1(\u0\/u2\/_0193_ ), .A2(\u0\/u2\/_0176_ ), .B1(\u0\/u2\/_0043_ ), .Y(\u0\/u2\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1007_ ( .A(\u0\/u2\/_0185_ ), .B(\u0\/u2\/_0189_ ), .C(\u0\/u2\/_0192_ ), .D(\u0\/u2\/_0195_ ), .X(\u0\/u2\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u2/_1008_ ( .A_N(\w3\[3\] ), .B(\u0\/u2\/_0734_ ), .C(\w3\[2\] ), .X(\u0\/u2\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1009_ ( .A(\u0\/u2\/_0137_ ), .B(\u0\/u2\/_0197_ ), .X(\u0\/u2\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_1010_ ( .A(\u0\/u2\/_0198_ ), .B(\u0\/u2\/_0040_ ), .Y(\u0\/u2\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1011_ ( .A(\u0\/u2\/_0293_ ), .B(\u0\/u2\/_0137_ ), .X(\u0\/u2\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1012_ ( .A(\u0\/u2\/_0200_ ), .Y(\u0\/u2\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1013_ ( .A(\u0\/u2\/_0137_ ), .B(\u0\/u2\/_0110_ ), .Y(\u0\/u2\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1014_ ( .A(\u0\/u2\/_0139_ ), .B(\u0\/u2\/_0020_ ), .Y(\u0\/u2\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1015_ ( .A(\u0\/u2\/_0199_ ), .B(\u0\/u2\/_0201_ ), .C(\u0\/u2\/_0202_ ), .D(\u0\/u2\/_0203_ ), .X(\u0\/u2\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u2/_1016_ ( .A1(\u0\/u2\/_0532_ ), .A2(\u0\/u2\/_0109_ ), .B1(\u0\/u2\/_0102_ ), .C1(\u0\/u2\/_0727_ ), .X(\u0\/u2\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1017_ ( .A(\u0\/u2\/_0022_ ), .B(\u0\/u2\/_0078_ ), .Y(\u0\/u2\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1018_ ( .A(\u0\/u2\/_0078_ ), .B(\u0\/u2\/_0142_ ), .Y(\u0\/u2\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1019_ ( .A(\u0\/u2\/_0207_ ), .B(\u0\/u2\/_0208_ ), .Y(\u0\/u2\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1020_ ( .A1(\u0\/u2\/_0094_ ), .A2(\u0\/u2\/_0176_ ), .B1(\u0\/u2\/_0206_ ), .C1(\u0\/u2\/_0209_ ), .Y(\u0\/u2\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1021_ ( .A(\u0\/u2\/_0662_ ), .B(\u0\/u2\/_0070_ ), .X(\u0\/u2\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u2/_1022_ ( .A(\u0\/u2\/_0731_ ), .B(\u0\/u2\/_0123_ ), .C(\u0\/u2\/_0749_ ), .Y(\u0\/u2\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u2/_1023_ ( .A(\u0\/u2\/_0731_ ), .B(\u0\/u2\/_0467_ ), .C(\u0\/u2\/_0069_ ), .Y(\u0\/u2\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u2/_1024_ ( .A_N(\u0\/u2\/_0211_ ), .B(\u0\/u2\/_0127_ ), .C(\u0\/u2\/_0212_ ), .D(\u0\/u2\/_0213_ ), .X(\u0\/u2\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1025_ ( .A(\u0\/u2\/_0137_ ), .Y(\u0\/u2\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1026_ ( .A(\u0\/u2\/_0128_ ), .B(\u0\/u2\/_0035_ ), .Y(\u0\/u2\/_0217_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1028_ ( .A1(\u0\/u2\/_0159_ ), .A2(\u0\/u2\/_0746_ ), .B1(\u0\/u2\/_0434_ ), .B2(\u0\/u2\/_0499_ ), .Y(\u0\/u2\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u2/_1029_ ( .A1(\u0\/u2\/_0116_ ), .A2(\u0\/u2\/_0215_ ), .B1(\u0\/u2\/_0217_ ), .C1(\u0\/u2\/_0219_ ), .X(\u0\/u2\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1030_ ( .A(\u0\/u2\/_0113_ ), .B(\u0\/u2\/_0746_ ), .X(\u0\/u2\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u2/_1031_ ( .A1(\u0\/u2\/_0098_ ), .A2(\u0\/u2\/_0746_ ), .B1(\u0\/u2\/_0434_ ), .B2(\u0\/u2\/_0750_ ), .X(\u0\/u2\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1032_ ( .A1(\u0\/u2\/_0047_ ), .A2(\u0\/u2\/_0113_ ), .B1(\u0\/u2\/_0221_ ), .C1(\u0\/u2\/_0222_ ), .Y(\u0\/u2\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u2/_1033_ ( .A1(\u0\/u2\/_0129_ ), .A2(\u0\/u2\/_0162_ ), .B1(\u0\/u2\/_0271_ ), .B2(\u0\/u2\/_0705_ ), .X(\u0\/u2\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1034_ ( .A1(\u0\/u2\/_0093_ ), .A2(\u0\/u2\/_0738_ ), .B1(\u0\/u2\/_0081_ ), .C1(\u0\/u2\/_0224_ ), .Y(\u0\/u2\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1035_ ( .A(\u0\/u2\/_0214_ ), .B(\u0\/u2\/_0220_ ), .C(\u0\/u2\/_0223_ ), .D(\u0\/u2\/_0225_ ), .X(\u0\/u2\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1036_ ( .A(\u0\/u2\/_0196_ ), .B(\u0\/u2\/_0204_ ), .C(\u0\/u2\/_0210_ ), .D(\u0\/u2\/_0226_ ), .X(\u0\/u2\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1037_ ( .A(\u0\/u2\/_0111_ ), .B(\u0\/u2\/_0554_ ), .X(\u0\/u2\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1038_ ( .A(\u0\/u2\/_0229_ ), .Y(\u0\/u2\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1039_ ( .A(\u0\/u2\/_0111_ ), .B(\u0\/u2\/_0129_ ), .Y(\u0\/u2\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1040_ ( .A(\u0\/u2\/_0017_ ), .B(\u0\/u2\/_0738_ ), .Y(\u0\/u2\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1041_ ( .A(\u0\/u2\/_0030_ ), .B(\u0\/u2\/_0304_ ), .Y(\u0\/u2\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1042_ ( .A(\u0\/u2\/_0230_ ), .B(\u0\/u2\/_0231_ ), .C(\u0\/u2\/_0232_ ), .D(\u0\/u2\/_0233_ ), .X(\u0\/u2\/_0234_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1043_ ( .A(\u0\/u2\/_0047_ ), .B(\u0\/u2\/_0478_ ), .X(\u0\/u2\/_0235_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u2/_1044_ ( .A1(\u0\/u2\/_0129_ ), .A2(\u0\/u2\/_0554_ ), .B1(\u0\/u2\/_0137_ ), .Y(\u0\/u2\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u2/_1045_ ( .A(\u0\/u2\/_0235_ ), .B(\u0\/u2\/_0049_ ), .C_N(\u0\/u2\/_0236_ ), .Y(\u0\/u2\/_0237_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1046_ ( .A(\u0\/u2\/_0047_ ), .B(\u0\/u2\/_0077_ ), .X(\u0\/u2\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1047_ ( .A(\u0\/u2\/_0070_ ), .B(\u0\/u2\/_0035_ ), .X(\u0\/u2\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u2/_1048_ ( .A1(\u0\/u2\/_0047_ ), .A2(\u0\/u2\/_0736_ ), .B1(\u0\/u2\/_0022_ ), .B2(\u0\/u2\/_0099_ ), .X(\u0\/u2\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u2/_1049_ ( .A(\u0\/u2\/_0239_ ), .B(\u0\/u2\/_0240_ ), .C(\u0\/u2\/_0241_ ), .Y(\u0\/u2\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1050_ ( .A(\u0\/u2\/_0554_ ), .B(\u0\/u2\/_0072_ ), .X(\u0\/u2\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u2/_1051_ ( .A1(\u0\/u2\/_0142_ ), .A2(\u0\/u2\/_0137_ ), .B1(\u0\/u2\/_0159_ ), .B2(\u0\/u2\/_0082_ ), .X(\u0\/u2\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1052_ ( .A1(\u0\/u2\/_0608_ ), .A2(\u0\/u2\/_0072_ ), .B1(\u0\/u2\/_0243_ ), .C1(\u0\/u2\/_0244_ ), .Y(\u0\/u2\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1053_ ( .A(\u0\/u2\/_0234_ ), .B(\u0\/u2\/_0237_ ), .C(\u0\/u2\/_0242_ ), .D(\u0\/u2\/_0245_ ), .X(\u0\/u2\/_0246_ ) );
sky130_fd_sc_hd__buf_2 \u0/u2/_1054_ ( .A(\u0\/u2\/_0027_ ), .X(\u0\/u2\/_0247_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u2/_1055_ ( .A1(\u0\/u2\/_0554_ ), .A2(\u0\/u2\/_0586_ ), .B1(\u0\/u2\/_0247_ ), .X(\u0\/u2\/_0248_ ) );
sky130_fd_sc_hd__and2_1 \u0/u2/_1056_ ( .A(\u0\/u2\/_0082_ ), .B(\u0\/u2\/_0478_ ), .X(\u0\/u2\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_1057_ ( .A(\u0\/u2\/_0079_ ), .X(\u0\/u2\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1058_ ( .A(\u0\/u2\/_0251_ ), .B(\u0\/u2\/_0478_ ), .X(\u0\/u2\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_1059_ ( .A(\u0\/u2\/_0250_ ), .B(\u0\/u2\/_0252_ ), .Y(\u0\/u2\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1060_ ( .A(\u0\/u2\/_0016_ ), .B(\u0\/u2\/_0064_ ), .Y(\u0\/u2\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_1061_ ( .A(\u0\/u2\/_0304_ ), .X(\u0\/u2\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1062_ ( .A(\u0\/u2\/_0255_ ), .B(\u0\/u2\/_0640_ ), .Y(\u0\/u2\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u2/_1063_ ( .A_N(\u0\/u2\/_0248_ ), .B(\u0\/u2\/_0253_ ), .C(\u0\/u2\/_0254_ ), .D(\u0\/u2\/_0256_ ), .X(\u0\/u2\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1064_ ( .A(\u0\/u2\/_0099_ ), .B(\u0\/u2\/_0110_ ), .X(\u0\/u2\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \u0/u2/_1065_ ( .A1(\u0\/u2\/_0161_ ), .A2(\u0\/u2\/_0130_ ), .B1(\u0\/u2\/_0258_ ), .Y(\u0\/u2\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1066_ ( .A(\u0\/u2\/_0194_ ), .B(\w3\[1\] ), .X(\u0\/u2\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1068_ ( .A(\u0\/u2\/_0261_ ), .B(\u0\/u2\/_0153_ ), .Y(\u0\/u2\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u2/_1069_ ( .A_N(\u0\/u2\/_0154_ ), .B(\u0\/u2\/_0259_ ), .C(\u0\/u2\/_0263_ ), .X(\u0\/u2\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1070_ ( .A(\u0\/u2\/_0246_ ), .B(\u0\/u2\/_0174_ ), .C(\u0\/u2\/_0257_ ), .D(\u0\/u2\/_0264_ ), .X(\u0\/u2\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u2/_1071_ ( .A1(\u0\/u2\/_0261_ ), .A2(\u0\/u2\/_0554_ ), .B1(\u0\/u2\/_0159_ ), .X(\u0\/u2\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1072_ ( .A(\u0\/u2\/_0746_ ), .B(\u0\/u2\/_0150_ ), .Y(\u0\/u2\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1073_ ( .A(\u0\/u2\/_0175_ ), .Y(\u0\/u2\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \u0/u2/_1074_ ( .A(\u0\/u2\/_0423_ ), .B(\u0\/u2\/_0123_ ), .C(\u0\/u2\/_0151_ ), .X(\u0\/u2\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1075_ ( .A(\u0\/u2\/_0268_ ), .B(\u0\/u2\/_0269_ ), .Y(\u0\/u2\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u2/_1076_ ( .A_N(\u0\/u2\/_0266_ ), .B(\u0\/u2\/_0267_ ), .C(\u0\/u2\/_0270_ ), .X(\u0\/u2\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1077_ ( .A(\u0\/u2\/_0554_ ), .B(\u0\/u2\/_0150_ ), .X(\u0\/u2\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1078_ ( .A(\u0\/u2\/_0273_ ), .Y(\u0\/u2\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1079_ ( .A1(\u0\/u2\/_0734_ ), .A2(\u0\/u2\/_0325_ ), .B1(\u0\/u2\/_0380_ ), .Y(\u0\/u2\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1080_ ( .A(\u0\/u2\/_0275_ ), .Y(\u0\/u2\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1081_ ( .A(\u0\/u2\/_0276_ ), .B(\u0\/u2\/_0153_ ), .Y(\u0\/u2\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \u0/u2/_1082_ ( .A(\u0\/u2\/_0272_ ), .B(\u0\/u2\/_0274_ ), .C(\u0\/u2\/_0277_ ), .X(\u0\/u2\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_1083_ ( .A(\u0\/u2\/_0035_ ), .X(\u0\/u2\/_0279_ ) );
sky130_fd_sc_hd__buf_2 \u0/u2/_1084_ ( .A(\u0\/u2\/_0082_ ), .X(\u0\/u2\/_0280_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1085_ ( .A1(\u0\/u2\/_0499_ ), .A2(\u0\/u2\/_0279_ ), .B1(\u0\/u2\/_0280_ ), .B2(\u0\/u2\/_0060_ ), .Y(\u0\/u2\/_0281_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1086_ ( .A1(\u0\/u2\/_0251_ ), .A2(\u0\/u2\/_0434_ ), .B1(\u0\/u2\/_0304_ ), .Y(\u0\/u2\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1087_ ( .A(\u0\/u2\/_0091_ ), .B(\u0\/u2\/_0056_ ), .Y(\u0\/u2\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1088_ ( .A1(\u0\/u2\/_0118_ ), .A2(\u0\/u2\/_0050_ ), .B1(\u0\/u2\/_0038_ ), .C1(\u0\/u2\/_0255_ ), .Y(\u0\/u2\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1089_ ( .A(\u0\/u2\/_0281_ ), .B(\u0\/u2\/_0283_ ), .C(\u0\/u2\/_0284_ ), .D(\u0\/u2\/_0285_ ), .X(\u0\/u2\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1090_ ( .A(\u0\/u2\/_0082_ ), .B(\u0\/u2\/_0027_ ), .X(\u0\/u2\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1091_ ( .A(\u0\/u2\/_0129_ ), .B(\u0\/u2\/_0027_ ), .X(\u0\/u2\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_1092_ ( .A(\u0\/u2\/_0287_ ), .B(\u0\/u2\/_0288_ ), .Y(\u0\/u2\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1093_ ( .A1(\u0\/u2\/_0752_ ), .A2(\u0\/u2\/_0683_ ), .B1(\u0\/u2\/_0093_ ), .B2(\u0\/u2\/_0247_ ), .Y(\u0\/u2\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1094_ ( .A1(\u0\/u2\/_0092_ ), .A2(\u0\/u2\/_0575_ ), .B1(\u0\/u2\/_0056_ ), .Y(\u0\/u2\/_0291_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1096_ ( .A1(\u0\/u2\/_0499_ ), .A2(\u0\/u2\/_0662_ ), .B1(\u0\/u2\/_0280_ ), .B2(\u0\/u2\/_0056_ ), .Y(\u0\/u2\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1097_ ( .A(\u0\/u2\/_0289_ ), .B(\u0\/u2\/_0290_ ), .C(\u0\/u2\/_0291_ ), .D(\u0\/u2\/_0294_ ), .X(\u0\/u2\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1098_ ( .A(\u0\/u2\/_0750_ ), .B(\u0\/u2\/_0193_ ), .X(\u0\/u2\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1099_ ( .A(\u0\/u2\/_0705_ ), .B(\u0\/u2\/_0380_ ), .X(\u0\/u2\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1100_ ( .A(\u0\/u2\/_0752_ ), .B(\u0\/u2\/_0129_ ), .Y(\u0\/u2\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u2/_1101_ ( .A(\u0\/u2\/_0296_ ), .B(\u0\/u2\/_0297_ ), .C_N(\u0\/u2\/_0298_ ), .Y(\u0\/u2\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1102_ ( .A(\u0\/u2\/_0089_ ), .B(\u0\/u2\/_0532_ ), .Y(\u0\/u2\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1103_ ( .A(\w3\[2\] ), .Y(\u0\/u2\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u2/_1104_ ( .A(\u0\/u2\/_0301_ ), .B(\w3\[3\] ), .C(\u0\/u2\/_0118_ ), .Y(\u0\/u2\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1105_ ( .A(\u0\/u2\/_0072_ ), .B(\u0\/u2\/_0302_ ), .X(\u0\/u2\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1106_ ( .A(\u0\/u2\/_0303_ ), .Y(\u0\/u2\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1107_ ( .A(\u0\/u2\/_0147_ ), .B(\u0\/u2\/_0302_ ), .Y(\u0\/u2\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1108_ ( .A(\u0\/u2\/_0299_ ), .B(\u0\/u2\/_0300_ ), .C(\u0\/u2\/_0305_ ), .D(\u0\/u2\/_0306_ ), .X(\u0\/u2\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1109_ ( .A(\u0\/u2\/_0278_ ), .B(\u0\/u2\/_0286_ ), .C(\u0\/u2\/_0295_ ), .D(\u0\/u2\/_0307_ ), .X(\u0\/u2\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u2/_1110_ ( .A(\u0\/u2\/_0228_ ), .B(\u0\/u2\/_0265_ ), .C(\u0\/u2\/_0308_ ), .Y(\u0\/u2\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1111_ ( .A(\u0\/u2\/_0235_ ), .Y(\u0\/u2\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1112_ ( .A(\u0\/u2\/_0478_ ), .B(\u0\/u2\/_0640_ ), .X(\u0\/u2\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1113_ ( .A(\u0\/u2\/_0310_ ), .Y(\u0\/u2\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1114_ ( .A(\u0\/u2\/_0022_ ), .B(\u0\/u2\/_0499_ ), .Y(\u0\/u2\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1115_ ( .A(\u0\/u2\/_0499_ ), .B(\u0\/u2\/_0032_ ), .Y(\u0\/u2\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1116_ ( .A(\u0\/u2\/_0309_ ), .B(\u0\/u2\/_0311_ ), .C(\u0\/u2\/_0312_ ), .D(\u0\/u2\/_0313_ ), .X(\u0\/u2\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1117_ ( .A(\u0\/u2\/_0499_ ), .B(\u0\/u2\/_0064_ ), .Y(\u0\/u2\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1118_ ( .A(\u0\/u2\/_0499_ ), .B(\u0\/u2\/_0683_ ), .Y(\u0\/u2\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1119_ ( .A(\u0\/u2\/_0315_ ), .B(\u0\/u2\/_0316_ ), .C(\u0\/u2\/_0317_ ), .D(\u0\/u2\/_0253_ ), .X(\u0\/u2\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1120_ ( .A(\u0\/u2\/_0047_ ), .B(\u0\/u2\/_0304_ ), .Y(\u0\/u2\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1121_ ( .A(\u0\/u2\/_0586_ ), .B(\u0\/u2\/_0162_ ), .Y(\u0\/u2\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1122_ ( .A(\u0\/u2\/_0319_ ), .B(\u0\/u2\/_0320_ ), .Y(\u0\/u2\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_1123_ ( .A(\u0\/u2\/_0321_ ), .B(\u0\/u2\/_0238_ ), .Y(\u0\/u2\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1124_ ( .A(\u0\/u2\/_0304_ ), .B(\u0\/u2\/_0062_ ), .Y(\u0\/u2\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_1125_ ( .A(\u0\/u2\/_0251_ ), .X(\u0\/u2\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1126_ ( .A1(\u0\/u2\/_0324_ ), .A2(\u0\/u2\/_0280_ ), .B1(\u0\/u2\/_0255_ ), .Y(\u0\/u2\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1127_ ( .A1(\u0\/u2\/_0050_ ), .A2(\u0\/u2\/_0216_ ), .B1(\u0\/u2\/_0109_ ), .C1(\u0\/u2\/_0255_ ), .Y(\u0\/u2\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1128_ ( .A(\u0\/u2\/_0322_ ), .B(\u0\/u2\/_0323_ ), .C(\u0\/u2\/_0326_ ), .D(\u0\/u2\/_0327_ ), .X(\u0\/u2\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1129_ ( .A1(\u0\/u2\/_0733_ ), .A2(\u0\/u2\/_0279_ ), .A3(\u0\/u2\/_0058_ ), .B1(\u0\/u2\/_0056_ ), .Y(\u0\/u2\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_1130_ ( .A(\u0\/u2\/_0047_ ), .X(\u0\/u2\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1131_ ( .A(\u0\/u2\/_0330_ ), .B(\u0\/u2\/_0056_ ), .Y(\u0\/u2\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1132_ ( .A(\u0\/u2\/_0054_ ), .B(\u0\/u2\/_0045_ ), .Y(\u0\/u2\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1133_ ( .A(\u0\/u2\/_0329_ ), .B(\u0\/u2\/_0331_ ), .C(\u0\/u2\/_0284_ ), .D(\u0\/u2\/_0332_ ), .X(\u0\/u2\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u2/_1134_ ( .A1(\u0\/u2\/_0543_ ), .A2(\u0\/u2\/_0216_ ), .B1(\u0\/u2\/_0532_ ), .C1(\u0\/u2\/_0060_ ), .X(\u0\/u2\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1135_ ( .A(\u0\/u2\/_0280_ ), .B(\u0\/u2\/_0060_ ), .Y(\u0\/u2\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1136_ ( .A(\u0\/u2\/_0324_ ), .B(\u0\/u2\/_0060_ ), .Y(\u0\/u2\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1137_ ( .A(\u0\/u2\/_0335_ ), .B(\u0\/u2\/_0337_ ), .Y(\u0\/u2\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1138_ ( .A1(\u0\/u2\/_0276_ ), .A2(\u0\/u2\/_0060_ ), .B1(\u0\/u2\/_0334_ ), .C1(\u0\/u2\/_0338_ ), .Y(\u0\/u2\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1139_ ( .A(\u0\/u2\/_0318_ ), .B(\u0\/u2\/_0328_ ), .C(\u0\/u2\/_0333_ ), .D(\u0\/u2\/_0339_ ), .X(\u0\/u2\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u2/_1140_ ( .A1(\u0\/u2\/_0746_ ), .A2(\u0\/u2\/_0456_ ), .B1(\u0\/u2\/_0128_ ), .X(\u0\/u2\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u2/_1141_ ( .A_N(\u0\/u2\/_0086_ ), .B(\u0\/u2\/_0128_ ), .X(\u0\/u2\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1142_ ( .A(\u0\/u2\/_0079_ ), .B(\u0\/u2\/_0124_ ), .X(\u0\/u2\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_1143_ ( .A(\u0\/u2\/_0126_ ), .B(\u0\/u2\/_0343_ ), .Y(\u0\/u2\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u2/_1144_ ( .A(\u0\/u2\/_0341_ ), .B(\u0\/u2\/_0342_ ), .C_N(\u0\/u2\/_0344_ ), .Y(\u0\/u2\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1146_ ( .A1(\u0\/u2\/_0193_ ), .A2(\u0\/u2\/_0092_ ), .A3(\u0\/u2\/_0330_ ), .B1(\u0\/u2\/_0147_ ), .Y(\u0\/u2\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1147_ ( .A1(\u0\/u2\/_0130_ ), .A2(\u0\/u2\/_0280_ ), .A3(\u0\/u2\/_0456_ ), .B1(\u0\/u2\/_0139_ ), .Y(\u0\/u2\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1148_ ( .A1(\u0\/u2\/_0144_ ), .A2(\u0\/u2\/_0608_ ), .A3(\u0\/u2\/_0092_ ), .B1(\u0\/u2\/_0139_ ), .Y(\u0\/u2\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1149_ ( .A(\u0\/u2\/_0345_ ), .B(\u0\/u2\/_0348_ ), .C(\u0\/u2\/_0349_ ), .D(\u0\/u2\/_0350_ ), .X(\u0\/u2\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \u0/u2/_1150_ ( .A(\u0\/u2\/_0150_ ), .B(\u0\/u2\/_0194_ ), .C(\u0\/u2\/_0543_ ), .X(\u0\/u2\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u2/_1151_ ( .A(\u0\/u2\/_0277_ ), .SLEEP(\u0\/u2\/_0352_ ), .X(\u0\/u2\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \u0/u2/_1152_ ( .A1(\u0\/u2\/_0268_ ), .A2(\u0\/u2\/_0171_ ), .B1(\u0\/u2\/_0157_ ), .Y(\u0\/u2\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u2/_1153_ ( .A(\u0\/u2\/_0161_ ), .X(\u0\/u2\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1154_ ( .A1(\u0\/u2\/_0279_ ), .A2(\u0\/u2\/_0280_ ), .B1(\u0\/u2\/_0355_ ), .Y(\u0\/u2\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1155_ ( .A1(\u0\/u2\/_0020_ ), .A2(\u0\/u2\/_0193_ ), .A3(\u0\/u2\/_0091_ ), .B1(\u0\/u2\/_0355_ ), .Y(\u0\/u2\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1156_ ( .A(\u0\/u2\/_0353_ ), .B(\u0\/u2\/_0354_ ), .C(\u0\/u2\/_0356_ ), .D(\u0\/u2\/_0357_ ), .X(\u0\/u2\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1157_ ( .A(\u0\/u2\/_0111_ ), .B(\u0\/u2\/_0586_ ), .X(\u0\/u2\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1158_ ( .A(\u0\/u2\/_0360_ ), .Y(\u0\/u2\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u2/_1159_ ( .A1(\u0\/u2\/_0119_ ), .A2(\u0\/u2\/_0120_ ), .B1(\u0\/u2\/_0230_ ), .C1(\u0\/u2\/_0361_ ), .X(\u0\/u2\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1160_ ( .A1(\u0\/u2\/_0662_ ), .A2(\u0\/u2\/_0251_ ), .A3(\u0\/u2\/_0456_ ), .B1(\u0\/u2\/_0114_ ), .Y(\u0\/u2\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1162_ ( .A1(\u0\/u2\/_0035_ ), .A2(\u0\/u2\/_0251_ ), .A3(\u0\/u2\/_0456_ ), .B1(\u0\/u2\/_0099_ ), .Y(\u0\/u2\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1163_ ( .A1(\u0\/u2\/_0193_ ), .A2(\u0\/u2\/_0608_ ), .B1(\u0\/u2\/_0099_ ), .Y(\u0\/u2\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1164_ ( .A(\u0\/u2\/_0362_ ), .B(\u0\/u2\/_0363_ ), .C(\u0\/u2\/_0365_ ), .D(\u0\/u2\/_0366_ ), .X(\u0\/u2\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1165_ ( .A1(\u0\/u2\/_0575_ ), .A2(\u0\/u2\/_0092_ ), .A3(\u0\/u2\/_0330_ ), .B1(\u0\/u2\/_0089_ ), .Y(\u0\/u2\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1166_ ( .A1(\u0\/u2\/_0586_ ), .A2(\u0\/u2\/_0017_ ), .A3(\u0\/u2\/_0330_ ), .B1(\u0\/u2\/_0094_ ), .Y(\u0\/u2\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u2/_1167_ ( .A1(\u0\/u2\/_0293_ ), .A2(\u0\/u2\/_0456_ ), .B1(\u0\/u2\/_0089_ ), .Y(\u0\/u2\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1168_ ( .A1(\u0\/u2\/_0279_ ), .A2(\u0\/u2\/_0456_ ), .B1(\u0\/u2\/_0094_ ), .Y(\u0\/u2\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1169_ ( .A(\u0\/u2\/_0368_ ), .B(\u0\/u2\/_0370_ ), .C(\u0\/u2\/_0371_ ), .D(\u0\/u2\/_0372_ ), .X(\u0\/u2\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1170_ ( .A(\u0\/u2\/_0351_ ), .B(\u0\/u2\/_0359_ ), .C(\u0\/u2\/_0367_ ), .D(\u0\/u2\/_0373_ ), .X(\u0\/u2\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1171_ ( .A1(\u0\/u2\/_0102_ ), .A2(\u0\/u2\/_0347_ ), .B1(\u0\/u2\/_0109_ ), .C1(\u0\/u2\/_0247_ ), .Y(\u0\/u2\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1172_ ( .A1(\u0\/u2\/_0102_ ), .A2(\u0\/u2\/_0347_ ), .B1(\u0\/u2\/_0532_ ), .C1(\u0\/u2\/_0247_ ), .Y(\u0\/u2\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1173_ ( .A1(\u0\/u2\/_0050_ ), .A2(\u0\/u2\/_0543_ ), .B1(\u0\/u2\/_0380_ ), .C1(\u0\/u2\/_0247_ ), .Y(\u0\/u2\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1174_ ( .A(\u0\/u2\/_0041_ ), .B(\u0\/u2\/_0375_ ), .C(\u0\/u2\/_0376_ ), .D(\u0\/u2\/_0377_ ), .X(\u0\/u2\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1175_ ( .A(\u0\/u2\/_0047_ ), .B(\u0\/u2\/_0750_ ), .X(\u0\/u2\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1176_ ( .A(\u0\/u2\/_0379_ ), .Y(\u0\/u2\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1177_ ( .A(\u0\/u2\/_0016_ ), .B(\u0\/u2\/_0608_ ), .Y(\u0\/u2\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1178_ ( .A(\u0\/u2\/_0752_ ), .B(\u0\/u2\/_0554_ ), .Y(\u0\/u2\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1179_ ( .A1(\w3\[1\] ), .A2(\u0\/u2\/_0734_ ), .B1(\u0\/u2\/_0109_ ), .C1(\u0\/u2\/_0016_ ), .Y(\u0\/u2\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1180_ ( .A(\u0\/u2\/_0381_ ), .B(\u0\/u2\/_0382_ ), .C(\u0\/u2\/_0383_ ), .D(\u0\/u2\/_0384_ ), .X(\u0\/u2\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \u0/u2/_1181_ ( .A(\u0\/u2\/_0086_ ), .B_N(\u0\/u2\/_0736_ ), .X(\u0\/u2\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1182_ ( .A1(\u0\/u2\/_0748_ ), .A2(\u0\/u2\/_0456_ ), .B1(\u0\/u2\/_0739_ ), .Y(\u0\/u2\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1183_ ( .A1(\u0\/u2\/_0118_ ), .A2(\u0\/u2\/_0543_ ), .B1(\u0\/u2\/_0109_ ), .C1(\u0\/u2\/_0739_ ), .Y(\u0\/u2\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1184_ ( .A1(\u0\/u2\/_0102_ ), .A2(\u0\/u2\/_0301_ ), .B1(\w3\[3\] ), .C1(\u0\/u2\/_0739_ ), .Y(\u0\/u2\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1185_ ( .A(\u0\/u2\/_0386_ ), .B(\u0\/u2\/_0387_ ), .C(\u0\/u2\/_0388_ ), .D(\u0\/u2\/_0389_ ), .X(\u0\/u2\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1186_ ( .A(\u0\/u2\/_0020_ ), .Y(\u0\/u2\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1187_ ( .A(\u0\/u2\/_0727_ ), .Y(\u0\/u2\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1188_ ( .A(\u0\/u2\/_0727_ ), .B(\u0\/u2\/_0064_ ), .Y(\u0\/u2\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1189_ ( .A1(\u0\/u2\/_0102_ ), .A2(\u0\/u2\/_0734_ ), .B1(\u0\/u2\/_0532_ ), .C1(\u0\/u2\/_0727_ ), .Y(\u0\/u2\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u2/_1190_ ( .A1(\u0\/u2\/_0392_ ), .A2(\u0\/u2\/_0393_ ), .B1(\u0\/u2\/_0394_ ), .C1(\u0\/u2\/_0395_ ), .X(\u0\/u2\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1191_ ( .A(\u0\/u2\/_0378_ ), .B(\u0\/u2\/_0385_ ), .C(\u0\/u2\/_0390_ ), .D(\u0\/u2\/_0396_ ), .X(\u0\/u2\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u2/_1192_ ( .A(\u0\/u2\/_0340_ ), .B(\u0\/u2\/_0374_ ), .C(\u0\/u2\/_0397_ ), .Y(\u0\/u2\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1193_ ( .A(\u0\/u2\/_0077_ ), .B(\u0\/u2\/_0129_ ), .X(\u0\/u2\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_1194_ ( .A(\u0\/u2\/_0398_ ), .B(\u0\/u2\/_0239_ ), .Y(\u0\/u2\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1195_ ( .A(\u0\/u2\/_0022_ ), .B(\u0\/u2\/_0111_ ), .X(\u0\/u2\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u2/_1196_ ( .A_N(\u0\/u2\/_0400_ ), .B(\u0\/u2\/_0231_ ), .Y(\u0\/u2\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u2/_1197_ ( .A(\u0\/u2\/_0399_ ), .SLEEP(\u0\/u2\/_0402_ ), .X(\u0\/u2\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_1198_ ( .A(\u0\/u2\/_0746_ ), .B(\u0\/u2\/_0251_ ), .Y(\u0\/u2\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u2/_1199_ ( .A_N(\u0\/u2\/_0404_ ), .B(\u0\/u2\/_0752_ ), .Y(\u0\/u2\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \u0/u2/_1200_ ( .A(\u0\/u2\/_0467_ ), .B(\u0\/u2\/_0194_ ), .C(\u0\/u2\/_0694_ ), .X(\u0\/u2\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u2/_1201_ ( .A_N(\u0\/u2\/_0175_ ), .B(\u0\/u2\/_0406_ ), .X(\u0\/u2\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1202_ ( .A(\u0\/u2\/_0407_ ), .Y(\u0\/u2\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1203_ ( .A1(\u0\/u2\/_0094_ ), .A2(\u0\/u2\/_0197_ ), .B1(\u0\/u2\/_0114_ ), .B2(\u0\/u2\/_0640_ ), .Y(\u0\/u2\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1204_ ( .A(\u0\/u2\/_0403_ ), .B(\u0\/u2\/_0405_ ), .C(\u0\/u2\/_0408_ ), .D(\u0\/u2\/_0409_ ), .X(\u0\/u2\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1205_ ( .A(\u0\/u2\/_0030_ ), .B(\u0\/u2\/_0150_ ), .Y(\u0\/u2\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u2/_1206_ ( .A_N(\u0\/u2\/_0169_ ), .B(\u0\/u2\/_0289_ ), .C(\u0\/u2\/_0411_ ), .X(\u0\/u2\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u2/_1207_ ( .A1(\u0\/u2\/_0467_ ), .A2(\u0\/u2\/_0151_ ), .B1(\u0\/u2\/_0140_ ), .C1(\u0\/u2\/_0129_ ), .X(\u0\/u2\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1208_ ( .A1(\u0\/u2\/_0608_ ), .A2(\u0\/u2\/_0099_ ), .B1(\u0\/u2\/_0037_ ), .C1(\u0\/u2\/_0414_ ), .Y(\u0\/u2\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1209_ ( .A(\u0\/u2\/_0738_ ), .Y(\u0\/u2\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1210_ ( .A(\u0\/u2\/_0586_ ), .B(\u0\/u2\/_0736_ ), .Y(\u0\/u2\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1211_ ( .A1(\u0\/u2\/_0194_ ), .A2(\u0\/u2\/_0038_ ), .B1(\u0\/u2\/_0118_ ), .C1(\u0\/u2\/_0153_ ), .Y(\u0\/u2\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u2/_1212_ ( .A1(\u0\/u2\/_0416_ ), .A2(\u0\/u2\/_0117_ ), .B1(\u0\/u2\/_0417_ ), .C1(\u0\/u2\/_0418_ ), .X(\u0\/u2\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1213_ ( .A(\u0\/u2\/_0077_ ), .B(\u0\/u2\/_0035_ ), .X(\u0\/u2\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1214_ ( .A(\u0\/u2\/_0662_ ), .B(\u0\/u2\/_0124_ ), .Y(\u0\/u2\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1215_ ( .A(\u0\/u2\/_0030_ ), .B(\u0\/u2\/_0137_ ), .Y(\u0\/u2\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1216_ ( .A(\u0\/u2\/_0072_ ), .B(\u0\/u2\/_0731_ ), .Y(\u0\/u2\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u2/_1217_ ( .A_N(\u0\/u2\/_0420_ ), .B(\u0\/u2\/_0421_ ), .C(\u0\/u2\/_0422_ ), .D(\u0\/u2\/_0424_ ), .X(\u0\/u2\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1218_ ( .A(\u0\/u2\/_0413_ ), .B(\u0\/u2\/_0415_ ), .C(\u0\/u2\/_0419_ ), .D(\u0\/u2\/_0425_ ), .X(\u0\/u2\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u2/_1219_ ( .A(\u0\/u2\/_0355_ ), .B(\u0\/u2\/_0102_ ), .C(\u0\/u2\/_0109_ ), .Y(\u0\/u2\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1220_ ( .A(\u0\/u2\/_0077_ ), .B(\u0\/u2\/_0017_ ), .X(\u0\/u2\/_0428_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1221_ ( .A(\u0\/u2\/_0077_ ), .B(\u0\/u2\/_0554_ ), .X(\u0\/u2\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u2/_1222_ ( .A1(\u0\/u2\/_0050_ ), .A2(\u0\/u2\/_0216_ ), .B1(\u0\/u2\/_0380_ ), .C1(\u0\/u2\/_0078_ ), .X(\u0\/u2\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u2/_1223_ ( .A(\u0\/u2\/_0428_ ), .B(\u0\/u2\/_0429_ ), .C(\u0\/u2\/_0430_ ), .Y(\u0\/u2\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u2/_1224_ ( .A_N(\u0\/u2\/_0209_ ), .B(\u0\/u2\/_0431_ ), .X(\u0\/u2\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u2/_1225_ ( .A1(\u0\/u2\/_0215_ ), .A2(\u0\/u2\/_0404_ ), .B1(\u0\/u2\/_0427_ ), .C1(\u0\/u2\/_0432_ ), .X(\u0\/u2\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1226_ ( .A(\u0\/u2\/_0043_ ), .B(\u0\/u2\/_0058_ ), .Y(\u0\/u2\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1227_ ( .A(\u0\/u2\/_0195_ ), .B(\u0\/u2\/_0233_ ), .C(\u0\/u2\/_0320_ ), .D(\u0\/u2\/_0435_ ), .X(\u0\/u2\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1228_ ( .A(\u0\/u2\/_0261_ ), .B(\u0\/u2\/_0738_ ), .Y(\u0\/u2\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1229_ ( .A1(\u0\/u2\/_0499_ ), .A2(\u0\/u2\/_0640_ ), .B1(\u0\/u2\/_0261_ ), .B2(\u0\/u2\/_0056_ ), .Y(\u0\/u2\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1230_ ( .A(\u0\/u2\/_0436_ ), .B(\u0\/u2\/_0394_ ), .C(\u0\/u2\/_0437_ ), .D(\u0\/u2\/_0438_ ), .X(\u0\/u2\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1231_ ( .A(\u0\/u2\/_0410_ ), .B(\u0\/u2\/_0426_ ), .C(\u0\/u2\/_0433_ ), .D(\u0\/u2\/_0439_ ), .X(\u0\/u2\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u2/_1232_ ( .A(\u0\/u2\/_0135_ ), .SLEEP(\u0\/u2\/_0273_ ), .X(\u0\/u2\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1233_ ( .A1(\u0\/u2\/_0279_ ), .A2(\u0\/u2\/_0456_ ), .B1(\u0\/u2\/_0099_ ), .Y(\u0\/u2\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1234_ ( .A(\u0\/u2\/_0441_ ), .B(\u0\/u2\/_0164_ ), .C(\u0\/u2\/_0270_ ), .D(\u0\/u2\/_0442_ ), .X(\u0\/u2\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1235_ ( .A(\u0\/u2\/_0051_ ), .B(\u0\/u2\/_0662_ ), .Y(\u0\/u2\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1236_ ( .A(\u0\/u2\/_0051_ ), .B(\u0\/u2\/_0271_ ), .Y(\u0\/u2\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1237_ ( .A(\u0\/u2\/_0444_ ), .B(\u0\/u2\/_0446_ ), .X(\u0\/u2\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1238_ ( .A(\u0\/u2\/_0193_ ), .B(\u0\/u2\/_0304_ ), .X(\u0\/u2\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1239_ ( .A(\u0\/u2\/_0448_ ), .Y(\u0\/u2\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1240_ ( .A(\u0\/u2\/_0162_ ), .B(\u0\/u2\/_0130_ ), .X(\u0\/u2\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1241_ ( .A(\u0\/u2\/_0450_ ), .Y(\u0\/u2\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1242_ ( .A1(\u0\/u2\/_0129_ ), .A2(\u0\/u2\/_0554_ ), .B1(\u0\/u2\/_0043_ ), .Y(\u0\/u2\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1243_ ( .A(\u0\/u2\/_0447_ ), .B(\u0\/u2\/_0449_ ), .C(\u0\/u2\/_0451_ ), .D(\u0\/u2\/_0452_ ), .X(\u0\/u2\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1244_ ( .A(\u0\/u2\/_0056_ ), .B(\u0\/u2\/_0064_ ), .Y(\u0\/u2\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u2/_1245_ ( .A_N(\u0\/u2\/_0248_ ), .B(\u0\/u2\/_0454_ ), .C(\u0\/u2\/_0254_ ), .D(\u0\/u2\/_0256_ ), .X(\u0\/u2\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1246_ ( .A1(\u0\/u2\/_0330_ ), .A2(\u0\/u2\/_0099_ ), .B1(\u0\/u2\/_0456_ ), .B2(\u0\/u2\/_0705_ ), .Y(\u0\/u2\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1247_ ( .A1(\u0\/u2\/_0748_ ), .A2(\u0\/u2\/_0738_ ), .B1(\u0\/u2\/_0092_ ), .B2(\u0\/u2\/_0752_ ), .Y(\u0\/u2\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1248_ ( .A1(\u0\/u2\/_0072_ ), .A2(\u0\/u2\/_0035_ ), .B1(\u0\/u2\/_0748_ ), .B2(\u0\/u2\/_0056_ ), .Y(\u0\/u2\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1249_ ( .A1(\u0\/u2\/_0748_ ), .A2(\u0\/u2\/_0251_ ), .B1(\u0\/u2\/_0247_ ), .Y(\u0\/u2\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1250_ ( .A(\u0\/u2\/_0457_ ), .B(\u0\/u2\/_0458_ ), .C(\u0\/u2\/_0459_ ), .D(\u0\/u2\/_0460_ ), .X(\u0\/u2\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1251_ ( .A(\u0\/u2\/_0443_ ), .B(\u0\/u2\/_0453_ ), .C(\u0\/u2\/_0455_ ), .D(\u0\/u2\/_0461_ ), .X(\u0\/u2\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1252_ ( .A(\u0\/u2\/_0705_ ), .B(\u0\/u2\/_0079_ ), .X(\u0\/u2\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1253_ ( .A(\u0\/u2\/_0586_ ), .B(\u0\/u2\/_0124_ ), .Y(\u0\/u2\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1254_ ( .A(\u0\/u2\/_0499_ ), .B(\u0\/u2\/_0746_ ), .Y(\u0\/u2\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u2/_1255_ ( .A_N(\u0\/u2\/_0463_ ), .B(\u0\/u2\/_0464_ ), .C(\u0\/u2\/_0465_ ), .X(\u0\/u2\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u2/_1256_ ( .A1(\u0\/u2\/_0271_ ), .A2(\u0\/u2\/_0072_ ), .B1(\u0\/u2\/_0142_ ), .B2(\u0\/u2\/_0027_ ), .X(\u0\/u2\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1257_ ( .A1(\u0\/u2\/_0144_ ), .A2(\u0\/u2\/_0099_ ), .B1(\u0\/u2\/_0360_ ), .C1(\u0\/u2\/_0468_ ), .Y(\u0\/u2\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u2/_1258_ ( .A1(\u0\/u2\/_0662_ ), .A2(\u0\/u2\/_0251_ ), .B1(\u0\/u2\/_0499_ ), .X(\u0\/u2\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1259_ ( .A1(\u0\/u2\/_0575_ ), .A2(\u0\/u2\/_0056_ ), .B1(\u0\/u2\/_0379_ ), .C1(\u0\/u2\/_0470_ ), .Y(\u0\/u2\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1260_ ( .A(\u0\/u2\/_0466_ ), .B(\u0\/u2\/_0469_ ), .C(\u0\/u2\/_0471_ ), .D(\u0\/u2\/_0305_ ), .X(\u0\/u2\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u2/_1261_ ( .A1(\u0\/u2\/_0247_ ), .A2(\u0\/u2\/_0683_ ), .B1(\u0\/u2\/_0324_ ), .B2(\u0\/u2\/_0056_ ), .X(\u0\/u2\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1262_ ( .A(\u0\/u2\/_0280_ ), .B(\u0\/u2\/_0099_ ), .X(\u0\/u2\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \u0/u2/_1263_ ( .A1(\u0\/u2\/_0092_ ), .A2(\u0\/u2\/_0247_ ), .B1(\u0\/u2\/_0474_ ), .X(\u0\/u2\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u2/_1264_ ( .A(\u0\/u2\/_0075_ ), .B(\u0\/u2\/_0473_ ), .C(\u0\/u2\/_0475_ ), .Y(\u0\/u2\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1265_ ( .A1(\u0\/u2\/_0279_ ), .A2(\u0\/u2\/_0255_ ), .B1(\u0\/u2\/_0280_ ), .B2(\u0\/u2\/_0060_ ), .Y(\u0\/u2\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1266_ ( .A1(\u0\/u2\/_0093_ ), .A2(\u0\/u2\/_0056_ ), .B1(\u0\/u2\/_0456_ ), .B2(\u0\/u2\/_0114_ ), .Y(\u0\/u2\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1267_ ( .A1(\u0\/u2\/_0161_ ), .A2(\u0\/u2\/_0032_ ), .B1(\u0\/u2\/_0324_ ), .B2(\u0\/u2\/_0147_ ), .Y(\u0\/u2\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1268_ ( .A1(\u0\/u2\/_0054_ ), .A2(\u0\/u2\/_0731_ ), .B1(\u0\/u2\/_0748_ ), .B2(\u0\/u2\/_0304_ ), .Y(\u0\/u2\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1269_ ( .A(\u0\/u2\/_0477_ ), .B(\u0\/u2\/_0479_ ), .C(\u0\/u2\/_0480_ ), .D(\u0\/u2\/_0481_ ), .X(\u0\/u2\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1270_ ( .A(\u0\/u2\/_0161_ ), .B(\u0\/u2\/_0064_ ), .Y(\u0\/u2\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u2/_1271_ ( .A(\u0\/u2\/_0731_ ), .B(\u0\/u2\/_0123_ ), .C(\u0\/u2\/_0467_ ), .Y(\u0\/u2\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1272_ ( .A(\u0\/u2\/_0483_ ), .B(\u0\/u2\/_0484_ ), .Y(\u0\/u2\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1273_ ( .A(\u0\/u2\/_0297_ ), .Y(\u0\/u2\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u2/_1274_ ( .A_N(\u0\/u2\/_0485_ ), .B(\u0\/u2\/_0181_ ), .C(\u0\/u2\/_0486_ ), .D(\u0\/u2\/_0386_ ), .X(\u0\/u2\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1275_ ( .A(\u0\/u2\/_0472_ ), .B(\u0\/u2\/_0476_ ), .C(\u0\/u2\/_0482_ ), .D(\u0\/u2\/_0487_ ), .X(\u0\/u2\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u2/_1276_ ( .A(\u0\/u2\/_0440_ ), .B(\u0\/u2\/_0462_ ), .C(\u0\/u2\/_0488_ ), .Y(\u0\/u2\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1277_ ( .A(\u0\/u2\/_0403_ ), .B(\u0\/u2\/_0230_ ), .C(\u0\/u2\/_0451_ ), .D(\u0\/u2\/_0361_ ), .X(\u0\/u2\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1278_ ( .A1(\u0\/u2\/_0118_ ), .A2(\u0\/u2\/_0050_ ), .B1(\u0\/u2\/_0109_ ), .C1(\u0\/u2\/_0139_ ), .Y(\u0\/u2\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1279_ ( .A(\u0\/u2\/_0447_ ), .B(\u0\/u2\/_0437_ ), .C(\u0\/u2\/_0491_ ), .D(\u0\/u2\/_0427_ ), .X(\u0\/u2\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1280_ ( .A1(\u0\/u2\/_0280_ ), .A2(\u0\/u2\/_0255_ ), .B1(\u0\/u2\/_0608_ ), .B2(\u0\/u2\/_0247_ ), .Y(\u0\/u2\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1281_ ( .A1(\u0\/u2\/_0144_ ), .A2(\u0\/u2\/_0147_ ), .B1(\u0\/u2\/_0355_ ), .B2(\u0\/u2\/_0093_ ), .Y(\u0\/u2\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1282_ ( .A1(\u0\/u2\/_0705_ ), .A2(\u0\/u2\/_0279_ ), .B1(\u0\/u2\/_0330_ ), .B2(\u0\/u2\/_0247_ ), .Y(\u0\/u2\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1283_ ( .A1(\u0\/u2\/_0279_ ), .A2(\u0\/u2\/_0280_ ), .B1(\u0\/u2\/_0114_ ), .Y(\u0\/u2\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1284_ ( .A(\u0\/u2\/_0493_ ), .B(\u0\/u2\/_0494_ ), .C(\u0\/u2\/_0495_ ), .D(\u0\/u2\/_0496_ ), .X(\u0\/u2\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1285_ ( .A1(\u0\/u2\/_0456_ ), .A2(\u0\/u2\/_0137_ ), .B1(\u0\/u2\/_0355_ ), .B2(\u0\/u2\/_0575_ ), .Y(\u0\/u2\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1286_ ( .A1(\u0\/u2\/_0099_ ), .A2(\u0\/u2\/_0733_ ), .B1(\u0\/u2\/_0093_ ), .B2(\u0\/u2\/_0499_ ), .Y(\u0\/u2\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1287_ ( .A(\u0\/u2\/_0147_ ), .B(\u0\/u2\/_0640_ ), .Y(\u0\/u2\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1288_ ( .A1(\u0\/u2\/_0153_ ), .A2(\u0\/u2\/_0056_ ), .B1(\u0\/u2\/_0748_ ), .Y(\u0\/u2\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1289_ ( .A(\u0\/u2\/_0498_ ), .B(\u0\/u2\/_0500_ ), .C(\u0\/u2\/_0501_ ), .D(\u0\/u2\/_0502_ ), .X(\u0\/u2\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1290_ ( .A(\u0\/u2\/_0490_ ), .B(\u0\/u2\/_0492_ ), .C(\u0\/u2\/_0497_ ), .D(\u0\/u2\/_0503_ ), .X(\u0\/u2\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u2/_1291_ ( .A_N(\u0\/u2\/_0275_ ), .B(\u0\/u2\/_0705_ ), .X(\u0\/u2\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1292_ ( .A(\u0\/u2\/_0505_ ), .Y(\u0\/u2\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1293_ ( .A(\u0\/u2\/_0380_ ), .B(\u0\/u2\/_0347_ ), .X(\u0\/u2\/_0507_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1294_ ( .A1(\u0\/u2\/_0507_ ), .A2(\u0\/u2\/_0093_ ), .B1(\u0\/u2\/_0056_ ), .Y(\u0\/u2\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1295_ ( .A(\u0\/u2\/_0322_ ), .B(\u0\/u2\/_0277_ ), .C(\u0\/u2\/_0506_ ), .D(\u0\/u2\/_0508_ ), .X(\u0\/u2\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1296_ ( .A(\u0\/u2\/_0280_ ), .B(\u0\/u2\/_0705_ ), .X(\u0\/u2\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1297_ ( .A1(\u0\/u2\/_0733_ ), .A2(\u0\/u2\/_0114_ ), .B1(\u0\/u2\/_0429_ ), .C1(\u0\/u2\/_0511_ ), .Y(\u0\/u2\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_1298_ ( .A(\u0\/u2\/_0019_ ), .B(\u0\/u2\/_0024_ ), .Y(\u0\/u2\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1299_ ( .A(\u0\/u2\/_0512_ ), .B(\u0\/u2\/_0513_ ), .C(\u0\/u2\/_0742_ ), .D(\u0\/u2\/_0306_ ), .X(\u0\/u2\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1300_ ( .A1(\u0\/u2\/_0532_ ), .A2(\u0\/u2\/_0089_ ), .B1(\u0\/u2\/_0154_ ), .C1(\u0\/u2\/_0169_ ), .Y(\u0\/u2\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u2/_1301_ ( .A1(\u0\/u2\/_0749_ ), .A2(\u0\/u2\/_0026_ ), .B1(\u0\/u2\/_0069_ ), .C1(\u0\/u2\/_0032_ ), .X(\u0\/u2\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u2/_1302_ ( .A1(\u0\/u2\/_0324_ ), .A2(\u0\/u2\/_0355_ ), .B1(\u0\/u2\/_0330_ ), .B2(\u0\/u2\/_0727_ ), .X(\u0\/u2\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u2/_1303_ ( .A(\u0\/u2\/_0133_ ), .B(\u0\/u2\/_0516_ ), .C(\u0\/u2\/_0517_ ), .Y(\u0\/u2\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1304_ ( .A(\u0\/u2\/_0509_ ), .B(\u0\/u2\/_0514_ ), .C(\u0\/u2\/_0515_ ), .D(\u0\/u2\/_0518_ ), .X(\u0\/u2\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1305_ ( .A(\u0\/u2\/_0746_ ), .B(\u0\/u2\/_0072_ ), .Y(\u0\/u2\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1306_ ( .A1(\u0\/u2\/_0082_ ), .A2(\u0\/u2\/_0070_ ), .B1(\u0\/u2\/_0043_ ), .B2(\u0\/u2\/_0193_ ), .Y(\u0\/u2\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1307_ ( .A(\u0\/u2\/_0311_ ), .B(\u0\/u2\/_0520_ ), .C(\u0\/u2\/_0332_ ), .D(\u0\/u2\/_0522_ ), .X(\u0\/u2\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1308_ ( .A(\u0\/u2\/_0129_ ), .B(\u0\/u2\/_0499_ ), .X(\u0\/u2\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_1309_ ( .A(\u0\/u2\/_0235_ ), .B(\u0\/u2\/_0524_ ), .Y(\u0\/u2\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u2/_1310_ ( .A(\u0\/u2\/_0081_ ), .B(\u0\/u2\/_0085_ ), .Y(\u0\/u2\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1311_ ( .A1(\u0\/u2\/_0051_ ), .A2(\u0\/u2\/_0045_ ), .B1(\u0\/u2\/_0130_ ), .B2(\u0\/u2\/_0094_ ), .Y(\u0\/u2\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1312_ ( .A(\u0\/u2\/_0523_ ), .B(\u0\/u2\/_0525_ ), .C(\u0\/u2\/_0526_ ), .D(\u0\/u2\/_0527_ ), .X(\u0\/u2\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u2/_1313_ ( .A_N(\u0\/u2\/_0250_ ), .B(\u0\/u2\/_0521_ ), .Y(\u0\/u2\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1314_ ( .A(\u0\/u2\/_0128_ ), .B(\u0\/u2\/_0020_ ), .X(\u0\/u2\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1315_ ( .A(\u0\/u2\/_0530_ ), .Y(\u0\/u2\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1316_ ( .A(\u0\/u2\/_0099_ ), .B(\u0\/u2\/_0058_ ), .X(\u0\/u2\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1317_ ( .A(\u0\/u2\/_0533_ ), .Y(\u0\/u2\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u2/_1318_ ( .A_N(\u0\/u2\/_0529_ ), .B(\u0\/u2\/_0531_ ), .C(\u0\/u2\/_0534_ ), .D(\u0\/u2\/_0192_ ), .X(\u0\/u2\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1319_ ( .A(\u0\/u2\/_0434_ ), .B(\u0\/u2\/_0078_ ), .X(\u0\/u2\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u2/_1320_ ( .A1(\u0\/u2\/_0750_ ), .A2(\u0\/u2\/_0079_ ), .B1(\u0\/u2\/_0129_ ), .B2(\u0\/u2\/_0705_ ), .X(\u0\/u2\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1321_ ( .A1(\u0\/u2\/_0161_ ), .A2(\u0\/u2\/_0032_ ), .B1(\u0\/u2\/_0536_ ), .C1(\u0\/u2\/_0537_ ), .Y(\u0\/u2\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u2/_1322_ ( .A1(\u0\/u2\/_0746_ ), .A2(\u0\/u2\/_0162_ ), .B1(\u0\/u2\/_0079_ ), .B2(\u0\/u2\/_0043_ ), .X(\u0\/u2\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1323_ ( .A1(\u0\/u2\/_0093_ ), .A2(\u0\/u2\/_0247_ ), .B1(\u0\/u2\/_0240_ ), .C1(\u0\/u2\/_0539_ ), .Y(\u0\/u2\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1324_ ( .A(\u0\/u2\/_0434_ ), .B(\u0\/u2\/_0043_ ), .X(\u0\/u2\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u2/_1325_ ( .A1(\u0\/u2\/_0142_ ), .A2(\u0\/u2\/_0150_ ), .B1(\u0\/u2\/_0022_ ), .B2(\u0\/u2\/_0137_ ), .X(\u0\/u2\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1326_ ( .A1(\u0\/u2\/_0279_ ), .A2(\u0\/u2\/_0051_ ), .B1(\u0\/u2\/_0541_ ), .C1(\u0\/u2\/_0542_ ), .Y(\u0\/u2\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1327_ ( .A(\u0\/u2\/_0159_ ), .B(\u0\/u2\/_0035_ ), .X(\u0\/u2\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u2/_1328_ ( .A1(\u0\/u2\/_0271_ ), .A2(\u0\/u2\/_0434_ ), .B1(\u0\/u2\/_0027_ ), .X(\u0\/u2\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1329_ ( .A1(\u0\/u2\/_0091_ ), .A2(\u0\/u2\/_0128_ ), .B1(\u0\/u2\/_0545_ ), .C1(\u0\/u2\/_0546_ ), .Y(\u0\/u2\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1330_ ( .A(\u0\/u2\/_0538_ ), .B(\u0\/u2\/_0540_ ), .C(\u0\/u2\/_0544_ ), .D(\u0\/u2\/_0547_ ), .X(\u0\/u2\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1331_ ( .A(\u0\/u2\/_0099_ ), .B(\u0\/u2\/_0193_ ), .X(\u0\/u2\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u2/_1332_ ( .A(\u0\/u2\/_0549_ ), .B(\u0\/u2\/_0186_ ), .C(\u0\/u2\/_0187_ ), .Y(\u0\/u2\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1333_ ( .A(\u0\/u2\/_0062_ ), .B(\u0\/u2\/_0347_ ), .C(\u0\/u2\/_0749_ ), .D(\u0\/u2\/_0694_ ), .X(\u0\/u2\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1334_ ( .A1(\u0\/u2\/_0130_ ), .A2(\u0\/u2\/_0499_ ), .B1(\u0\/u2\/_0551_ ), .C1(\u0\/u2\/_0101_ ), .Y(\u0\/u2\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1335_ ( .A(\u0\/u2\/_0139_ ), .B(\u0\/u2\/_0640_ ), .Y(\u0\/u2\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1336_ ( .A1(\u0\/u2\/_0752_ ), .A2(\u0\/u2\/_0662_ ), .B1(\u0\/u2\/_0280_ ), .B2(\u0\/u2\/_0099_ ), .Y(\u0\/u2\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1337_ ( .A(\u0\/u2\/_0550_ ), .B(\u0\/u2\/_0552_ ), .C(\u0\/u2\/_0553_ ), .D(\u0\/u2\/_0555_ ), .X(\u0\/u2\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1338_ ( .A(\u0\/u2\/_0528_ ), .B(\u0\/u2\/_0535_ ), .C(\u0\/u2\/_0548_ ), .D(\u0\/u2\/_0556_ ), .X(\u0\/u2\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u2/_1339_ ( .A(\u0\/u2\/_0504_ ), .B(\u0\/u2\/_0519_ ), .C(\u0\/u2\/_0557_ ), .Y(\u0\/u2\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1340_ ( .A(\u0\/u2\/_0054_ ), .B(\u0\/u2\/_0507_ ), .X(\u0\/u2\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u2/_1341_ ( .A_N(\u0\/u2\/_0558_ ), .B(\u0\/u2\/_0408_ ), .C(\u0\/u2\/_0451_ ), .D(\u0\/u2\/_0452_ ), .X(\u0\/u2\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1342_ ( .A(\u0\/u2\/_0549_ ), .Y(\u0\/u2\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1343_ ( .A(\u0\/u2\/_0559_ ), .B(\u0\/u2\/_0403_ ), .C(\u0\/u2\/_0560_ ), .D(\u0\/u2\/_0371_ ), .X(\u0\/u2\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1344_ ( .A(\u0\/u2\/_0181_ ), .B(\u0\/u2\/_0178_ ), .X(\u0\/u2\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1345_ ( .A(\u0\/u2\/_0562_ ), .B(\u0\/u2\/_0552_ ), .C(\u0\/u2\/_0553_ ), .D(\u0\/u2\/_0555_ ), .X(\u0\/u2\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1346_ ( .A(\u0\/u2\/_0247_ ), .B(\u0\/u2\/_0020_ ), .Y(\u0\/u2\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1347_ ( .A(\u0\/u2\/_0051_ ), .B(\u0\/u2\/_0130_ ), .X(\u0\/u2\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1348_ ( .A(\u0\/u2\/_0566_ ), .Y(\u0\/u2\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1349_ ( .A(\u0\/u2\/_0159_ ), .B(\u0\/u2\/_0423_ ), .X(\u0\/u2\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1350_ ( .A1(\u0\/u2\/_0752_ ), .A2(\u0\/u2\/_0640_ ), .B1(\u0\/u2\/_0568_ ), .B2(\u0\/u2\/_0175_ ), .Y(\u0\/u2\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1351_ ( .A(\u0\/u2\/_0076_ ), .B(\u0\/u2\/_0565_ ), .C(\u0\/u2\/_0567_ ), .D(\u0\/u2\/_0569_ ), .X(\u0\/u2\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u2/_1352_ ( .A1(\u0\/u2\/_0035_ ), .A2(\u0\/u2\/_0142_ ), .B1(\u0\/u2\/_0161_ ), .X(\u0\/u2\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1353_ ( .A(\u0\/u2\/_0099_ ), .B(\u0\/u2\/_0662_ ), .Y(\u0\/u2\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u2/_1354_ ( .A(\u0\/u2\/_0420_ ), .B(\u0\/u2\/_0571_ ), .C_N(\u0\/u2\/_0572_ ), .Y(\u0\/u2\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1355_ ( .A(\u0\/u2\/_0051_ ), .B(\u0\/u2\/_0746_ ), .Y(\u0\/u2\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1356_ ( .A(\u0\/u2\/_0574_ ), .B(\u0\/u2\/_0319_ ), .C(\u0\/u2\/_0320_ ), .D(\u0\/u2\/_0411_ ), .X(\u0\/u2\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1357_ ( .A(\u0\/u2\/_0736_ ), .B(\u0\/u2\/_0035_ ), .Y(\u0\/u2\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1358_ ( .A(\u0\/u2\/_0736_ ), .B(\u0\/u2\/_0030_ ), .Y(\u0\/u2\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1359_ ( .A(\u0\/u2\/_0298_ ), .B(\u0\/u2\/_0208_ ), .C(\u0\/u2\/_0577_ ), .D(\u0\/u2\/_0578_ ), .X(\u0\/u2\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1360_ ( .A1(\u0\/u2\/_0020_ ), .A2(\u0\/u2\/_0137_ ), .B1(\u0\/u2\/_0261_ ), .B2(\u0\/u2\/_0128_ ), .Y(\u0\/u2\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1361_ ( .A(\u0\/u2\/_0573_ ), .B(\u0\/u2\/_0576_ ), .C(\u0\/u2\/_0579_ ), .D(\u0\/u2\/_0580_ ), .X(\u0\/u2\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1362_ ( .A(\u0\/u2\/_0561_ ), .B(\u0\/u2\/_0563_ ), .C(\u0\/u2\/_0570_ ), .D(\u0\/u2\/_0581_ ), .X(\u0\/u2\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1363_ ( .A(\u0\/u2\/_0128_ ), .B(\u0\/u2\/_0193_ ), .X(\u0\/u2\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1364_ ( .A(\u0\/u2\/_0082_ ), .B(\u0\/u2\/_0162_ ), .X(\u0\/u2\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u2/_1365_ ( .A(\u0\/u2\/_0583_ ), .B(\u0\/u2\/_0584_ ), .C_N(\u0\/u2\/_0437_ ), .Y(\u0\/u2\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u2/_1366_ ( .A(\u0\/u2\/_0150_ ), .B(\u0\/u2\/_0118_ ), .C(\u0\/u2\/_0380_ ), .Y(\u0\/u2\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u2/_1367_ ( .A_N(\u0\/u2\/_0182_ ), .B(\u0\/u2\/_0587_ ), .C(\u0\/u2\/_0323_ ), .X(\u0\/u2\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1368_ ( .A1(\u0\/u2\/_0575_ ), .A2(\u0\/u2\/_0153_ ), .B1(\u0\/u2\/_0727_ ), .B2(\u0\/u2\/_0058_ ), .Y(\u0\/u2\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1369_ ( .A1(\u0\/u2\/_0499_ ), .A2(\u0\/u2\/_0064_ ), .B1(\u0\/u2\/_0456_ ), .B2(\u0\/u2\/_0255_ ), .Y(\u0\/u2\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1370_ ( .A(\u0\/u2\/_0585_ ), .B(\u0\/u2\/_0588_ ), .C(\u0\/u2\/_0589_ ), .D(\u0\/u2\/_0590_ ), .X(\u0\/u2\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \u0/u2/_1371_ ( .A1(\u0\/u2\/_0091_ ), .A2(\u0\/u2\/_0139_ ), .B1(\u0\/u2\/_0250_ ), .Y(\u0\/u2\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1372_ ( .A1(\u0\/u2\/_0092_ ), .A2(\u0\/u2\/_0739_ ), .B1(\u0\/u2\/_0324_ ), .B2(\u0\/u2\/_0247_ ), .Y(\u0\/u2\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1373_ ( .A1(\u0\/u2\/_0144_ ), .A2(\u0\/u2\/_0153_ ), .B1(\u0\/u2\/_0683_ ), .B2(\u0\/u2\/_0056_ ), .Y(\u0\/u2\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1374_ ( .A1(\u0\/u2\/_0091_ ), .A2(\u0\/u2\/_0499_ ), .B1(\u0\/u2\/_0330_ ), .B2(\u0\/u2\/_0056_ ), .Y(\u0\/u2\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1375_ ( .A(\u0\/u2\/_0592_ ), .B(\u0\/u2\/_0593_ ), .C(\u0\/u2\/_0594_ ), .D(\u0\/u2\/_0595_ ), .X(\u0\/u2\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1376_ ( .A(\u0\/u2\/_0499_ ), .B(\u0\/u2\/_0144_ ), .Y(\u0\/u2\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1377_ ( .A(\u0\/u2\/_0312_ ), .B(\u0\/u2\/_0598_ ), .Y(\u0\/u2\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1378_ ( .A(\u0\/u2\/_0575_ ), .B(\u0\/u2\/_0147_ ), .Y(\u0\/u2\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1379_ ( .A1(\u0\/u2\/_0293_ ), .A2(\u0\/u2\/_0137_ ), .B1(\u0\/u2\/_0093_ ), .B2(\u0\/u2\/_0739_ ), .Y(\u0\/u2\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1380_ ( .A1(\u0\/u2\/_0734_ ), .A2(\u0\/u2\/_0531_ ), .B1(\u0\/u2\/_0600_ ), .C1(\u0\/u2\/_0601_ ), .Y(\u0\/u2\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1381_ ( .A1(\u0\/u2\/_0153_ ), .A2(\u0\/u2\/_0261_ ), .B1(\u0\/u2\/_0599_ ), .C1(\u0\/u2\/_0602_ ), .Y(\u0\/u2\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1382_ ( .A(\u0\/u2\/_0591_ ), .B(\u0\/u2\/_0596_ ), .C(\u0\/u2\/_0174_ ), .D(\u0\/u2\/_0603_ ), .X(\u0\/u2\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1383_ ( .A(\u0\/u2\/_0247_ ), .B(\u0\/u2\/_0144_ ), .Y(\u0\/u2\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1384_ ( .A(\u0\/u2\/_0113_ ), .B(\u0\/u2\/_0017_ ), .Y(\u0\/u2\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1385_ ( .A(\u0\/u2\/_0381_ ), .B(\u0\/u2\/_0605_ ), .C(\u0\/u2\/_0361_ ), .D(\u0\/u2\/_0606_ ), .X(\u0\/u2\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1386_ ( .A1(\u0\/u2\/_0016_ ), .A2(\u0\/u2\/_0727_ ), .B1(\u0\/u2\/_0733_ ), .Y(\u0\/u2\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1387_ ( .A1(\u0\/u2\/_0586_ ), .A2(\u0\/u2\/_0159_ ), .B1(\u0\/u2\/_0082_ ), .B2(\u0\/u2\/_0750_ ), .Y(\u0\/u2\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1388_ ( .A1(\u0\/u2\/_0142_ ), .A2(\u0\/u2\/_0162_ ), .B1(\u0\/u2\/_0079_ ), .B2(\u0\/u2\/_0054_ ), .Y(\u0\/u2\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1389_ ( .A(\u0\/u2\/_0610_ ), .B(\u0\/u2\/_0611_ ), .C(\u0\/u2\/_0105_ ), .D(\u0\/u2\/_0106_ ), .X(\u0\/u2\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1390_ ( .A1(\u0\/u2\/_0094_ ), .A2(\u0\/u2\/_0302_ ), .B1(\u0\/u2\/_0324_ ), .B2(\u0\/u2\/_0089_ ), .Y(\u0\/u2\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1391_ ( .A(\u0\/u2\/_0607_ ), .B(\u0\/u2\/_0609_ ), .C(\u0\/u2\/_0612_ ), .D(\u0\/u2\/_0613_ ), .X(\u0\/u2\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1392_ ( .A(\u0\/u2\/_0041_ ), .B(\u0\/u2\/_0170_ ), .X(\u0\/u2\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1393_ ( .A(\u0\/u2\/_0554_ ), .B(\u0\/u2\/_0027_ ), .X(\u0\/u2\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1394_ ( .A(\u0\/u2\/_0027_ ), .B(\u0\/u2\/_0261_ ), .Y(\u0\/u2\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u2/_1395_ ( .A_N(\u0\/u2\/_0616_ ), .B(\u0\/u2\/_0617_ ), .Y(\u0\/u2\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1396_ ( .A1(\u0\/u2\/_0147_ ), .A2(\u0\/u2\/_0302_ ), .B1(\u0\/u2\/_0342_ ), .C1(\u0\/u2\/_0618_ ), .Y(\u0\/u2\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1397_ ( .A(\u0\/u2\/_0614_ ), .B(\u0\/u2\/_0272_ ), .C(\u0\/u2\/_0615_ ), .D(\u0\/u2\/_0620_ ), .X(\u0\/u2\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u2/_1398_ ( .A(\u0\/u2\/_0582_ ), .B(\u0\/u2\/_0604_ ), .C(\u0\/u2\/_0621_ ), .Y(\u0\/u2\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1399_ ( .A1(\u0\/u2\/_0280_ ), .A2(\u0\/u2\/_0456_ ), .B1(\u0\/u2\/_0089_ ), .Y(\u0\/u2\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1400_ ( .A1(\u0\/u2\/_0144_ ), .A2(\u0\/u2\/_0608_ ), .A3(\u0\/u2\/_0330_ ), .B1(\u0\/u2\/_0089_ ), .Y(\u0\/u2\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1401_ ( .A1(\u0\/u2\/_0197_ ), .A2(\u0\/u2\/_0130_ ), .A3(\u0\/u2\/_0110_ ), .B1(\u0\/u2\/_0094_ ), .Y(\u0\/u2\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1402_ ( .A(\u0\/u2\/_0432_ ), .B(\u0\/u2\/_0622_ ), .C(\u0\/u2\/_0623_ ), .D(\u0\/u2\/_0624_ ), .X(\u0\/u2\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \u0/u2/_1403_ ( .A1(\u0\/u2\/_0554_ ), .A2(\u0\/u2\/_0017_ ), .A3(\u0\/u2\/_0022_ ), .B1(\u0\/u2\/_0161_ ), .X(\u0\/u2\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u2/_1404_ ( .A_N(\u0\/u2\/_0269_ ), .B(\u0\/u2\/_0170_ ), .X(\u0\/u2\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1405_ ( .A1(\u0\/u2\/_0109_ ), .A2(\u0\/u2\/_0064_ ), .A3(\u0\/u2\/_0733_ ), .B1(\u0\/u2\/_0355_ ), .Y(\u0\/u2\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u2/_1406_ ( .A_N(\u0\/u2\/_0626_ ), .B(\u0\/u2\/_0627_ ), .C(\u0\/u2\/_0353_ ), .D(\u0\/u2\/_0628_ ), .X(\u0\/u2\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1407_ ( .A1(\u0\/u2\/_0091_ ), .A2(\u0\/u2\/_0110_ ), .A3(\u0\/u2\/_0176_ ), .B1(\u0\/u2\/_0139_ ), .Y(\u0\/u2\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1408_ ( .A1(\u0\/u2\/_0020_ ), .A2(\u0\/u2\/_0261_ ), .B1(\u0\/u2\/_0147_ ), .Y(\u0\/u2\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1409_ ( .A(\u0\/u2\/_0631_ ), .B(\u0\/u2\/_0344_ ), .C(\u0\/u2\/_0421_ ), .D(\u0\/u2\/_0632_ ), .X(\u0\/u2\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u2/_1410_ ( .A1(\u0\/u2\/_0325_ ), .A2(\u0\/u2\/_0734_ ), .B1(\u0\/u2\/_0038_ ), .C1(\u0\/u2\/_0113_ ), .X(\u0\/u2\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1411_ ( .A1(\u0\/u2\/_0456_ ), .A2(\u0\/u2\/_0114_ ), .B1(\u0\/u2\/_0221_ ), .C1(\u0\/u2\/_0634_ ), .Y(\u0\/u2\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u2/_1412_ ( .A(\u0\/u2\/_0119_ ), .B_N(\u0\/u2\/_0111_ ), .Y(\u0\/u2\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1413_ ( .A1(\u0\/u2\/_0032_ ), .A2(\u0\/u2\/_0113_ ), .B1(\u0\/u2\/_0636_ ), .C1(\u0\/u2\/_0400_ ), .Y(\u0\/u2\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1414_ ( .A1(\u0\/u2\/_0731_ ), .A2(\u0\/u2\/_0293_ ), .A3(\u0\/u2\/_0251_ ), .B1(\u0\/u2\/_0099_ ), .Y(\u0\/u2\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1415_ ( .A(\u0\/u2\/_0189_ ), .B(\u0\/u2\/_0635_ ), .C(\u0\/u2\/_0637_ ), .D(\u0\/u2\/_0638_ ), .X(\u0\/u2\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1416_ ( .A(\u0\/u2\/_0625_ ), .B(\u0\/u2\/_0630_ ), .C(\u0\/u2\/_0633_ ), .D(\u0\/u2\/_0639_ ), .X(\u0\/u2\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1417_ ( .A(\u0\/u2\/_0746_ ), .B(\u0\/u2\/_0738_ ), .X(\u0\/u2\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1418_ ( .A(\u0\/u2\/_0736_ ), .B(\u0\/u2\/_0731_ ), .X(\u0\/u2\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u2/_1419_ ( .A_N(\u0\/u2\/_0643_ ), .B(\u0\/u2\/_0577_ ), .Y(\u0\/u2\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1420_ ( .A1(\u0\/u2\/_0280_ ), .A2(\u0\/u2\/_0739_ ), .B1(\u0\/u2\/_0642_ ), .C1(\u0\/u2\/_0644_ ), .Y(\u0\/u2\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1421_ ( .A1(\u0\/u2\/_0050_ ), .A2(\u0\/u2\/_0543_ ), .B1(\u0\/u2\/_0194_ ), .C1(\u0\/u2\/_0738_ ), .Y(\u0\/u2\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1422_ ( .A(\u0\/u2\/_0646_ ), .B(\u0\/u2\/_0232_ ), .C(\u0\/u2\/_0417_ ), .D(\u0\/u2\/_0578_ ), .X(\u0\/u2\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1423_ ( .A1(\u0\/u2\/_0064_ ), .A2(\u0\/u2\/_0733_ ), .B1(\u0\/u2\/_0727_ ), .Y(\u0\/u2\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1424_ ( .A1(\u0\/u2\/_0193_ ), .A2(\u0\/u2\/_0276_ ), .B1(\u0\/u2\/_0727_ ), .Y(\u0\/u2\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1425_ ( .A(\u0\/u2\/_0645_ ), .B(\u0\/u2\/_0647_ ), .C(\u0\/u2\/_0648_ ), .D(\u0\/u2\/_0649_ ), .X(\u0\/u2\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1426_ ( .A1(\u0\/u2\/_0325_ ), .A2(\u0\/u2\/_0734_ ), .B1(\u0\/u2\/_0038_ ), .C1(\u0\/u2\/_0247_ ), .Y(\u0\/u2\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1427_ ( .A1(\u0\/u2\/_0543_ ), .A2(\u0\/u2\/_0216_ ), .B1(\u0\/u2\/_0423_ ), .C1(\u0\/u2\/_0247_ ), .Y(\u0\/u2\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1428_ ( .A(\u0\/u2\/_0652_ ), .B(\u0\/u2\/_0653_ ), .X(\u0\/u2\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1429_ ( .A1(\u0\/u2\/_0733_ ), .A2(\u0\/u2\/_0748_ ), .A3(\u0\/u2\/_0324_ ), .B1(\u0\/u2\/_0016_ ), .Y(\u0\/u2\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1430_ ( .A1(\u0\/u2\/_0640_ ), .A2(\u0\/u2\/_0193_ ), .A3(\u0\/u2\/_0091_ ), .B1(\u0\/u2\/_0016_ ), .Y(\u0\/u2\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1431_ ( .A1(\u0\/u2\/_0102_ ), .A2(\u0\/u2\/_0301_ ), .B1(\w3\[3\] ), .C1(\u0\/u2\/_0247_ ), .Y(\u0\/u2\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1432_ ( .A(\u0\/u2\/_0654_ ), .B(\u0\/u2\/_0655_ ), .C(\u0\/u2\/_0656_ ), .D(\u0\/u2\/_0657_ ), .X(\u0\/u2\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1433_ ( .A1(\u0\/u2\/_0118_ ), .A2(\u0\/u2\/_0050_ ), .B1(\u0\/u2\/_0038_ ), .C1(\u0\/u2\/_0478_ ), .Y(\u0\/u2\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u2/_1434_ ( .A_N(\u0\/u2\/_0250_ ), .B(\u0\/u2\/_0465_ ), .C(\u0\/u2\/_0659_ ), .X(\u0\/u2\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1435_ ( .A1(\u0\/u2\/_0683_ ), .A2(\u0\/u2\/_0324_ ), .B1(\u0\/u2\/_0255_ ), .Y(\u0\/u2\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1436_ ( .A1(\u0\/u2\/_0032_ ), .A2(\u0\/u2\/_0193_ ), .A3(\u0\/u2\/_0047_ ), .B1(\u0\/u2\/_0255_ ), .Y(\u0\/u2\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1437_ ( .A1(\u0\/u2\/_0144_ ), .A2(\u0\/u2\/_0586_ ), .A3(\u0\/u2\/_0047_ ), .B1(\u0\/u2\/_0499_ ), .Y(\u0\/u2\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1438_ ( .A(\u0\/u2\/_0660_ ), .B(\u0\/u2\/_0661_ ), .C(\u0\/u2\/_0663_ ), .D(\u0\/u2\/_0664_ ), .X(\u0\/u2\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1439_ ( .A1(\u0\/u2\/_0091_ ), .A2(\u0\/u2\/_0276_ ), .B1(\u0\/u2\/_0060_ ), .Y(\u0\/u2\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1440_ ( .A1(\u0\/u2\/_0144_ ), .A2(\u0\/u2\/_0608_ ), .B1(\u0\/u2\/_0056_ ), .Y(\u0\/u2\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1441_ ( .A1(\u0\/u2\/_0423_ ), .A2(\u0\/u2\/_0038_ ), .B1(\u0\/u2\/_0102_ ), .C1(\u0\/u2\/_0060_ ), .Y(\u0\/u2\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1442_ ( .A1(\w3\[1\] ), .A2(\u0\/u2\/_0734_ ), .B1(\u0\/u2\/_0109_ ), .C1(\u0\/u2\/_0056_ ), .Y(\u0\/u2\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1443_ ( .A(\u0\/u2\/_0666_ ), .B(\u0\/u2\/_0667_ ), .C(\u0\/u2\/_0668_ ), .D(\u0\/u2\/_0669_ ), .X(\u0\/u2\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1444_ ( .A(\u0\/u2\/_0650_ ), .B(\u0\/u2\/_0658_ ), .C(\u0\/u2\/_0665_ ), .D(\u0\/u2\/_0670_ ), .X(\u0\/u2\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u2/_1445_ ( .A(\u0\/u2\/_0641_ ), .B(\u0\/u2\/_0174_ ), .C(\u0\/u2\/_0671_ ), .Y(\u0\/u2\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u2/_1446_ ( .A(\u0\/u2\/_0049_ ), .B(\u0\/u2\/_0618_ ), .C_N(\u0\/u2\/_0052_ ), .Y(\u0\/u2\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \u0/u2/_1447_ ( .A(\u0\/u2\/_0239_ ), .Y(\u0\/u2\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1448_ ( .A(\u0\/u2\/_0705_ ), .B(\u0\/u2\/_0032_ ), .Y(\u0\/u2\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1449_ ( .A1(\u0\/u2\/_0054_ ), .A2(\u0\/u2\/_0731_ ), .B1(\u0\/u2\/_0035_ ), .B2(\u0\/u2\/_0705_ ), .Y(\u0\/u2\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1450_ ( .A1(\u0\/u2\/_0304_ ), .A2(\u0\/u2\/_0731_ ), .B1(\u0\/u2\/_0047_ ), .B2(\u0\/u2\/_0750_ ), .Y(\u0\/u2\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1451_ ( .A(\u0\/u2\/_0674_ ), .B(\u0\/u2\/_0675_ ), .C(\u0\/u2\/_0676_ ), .D(\u0\/u2\/_0677_ ), .X(\u0\/u2\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u2/_1452_ ( .A_N(\u0\/u2\/_0584_ ), .B(\u0\/u2\/_0283_ ), .X(\u0\/u2\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1453_ ( .A(\u0\/u2\/_0673_ ), .B(\u0\/u2\/_0678_ ), .C(\u0\/u2\/_0679_ ), .D(\u0\/u2\/_0508_ ), .X(\u0\/u2\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1454_ ( .A1(\u0\/u2\/_0016_ ), .A2(\u0\/u2\/_0733_ ), .B1(\u0\/u2\/_0355_ ), .B2(\u0\/u2\/_0092_ ), .Y(\u0\/u2\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1455_ ( .A(\u0\/u2\/_0681_ ), .B(\u0\/u2\/_0034_ ), .X(\u0\/u2\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u2/_1456_ ( .A1(\u0\/u2\/_0330_ ), .A2(\u0\/u2\/_0139_ ), .B1(\u0\/u2\/_0324_ ), .B2(\u0\/u2\/_0089_ ), .X(\u0\/u2\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1457_ ( .A1(\u0\/u2\/_0146_ ), .A2(\u0\/u2\/_0147_ ), .B1(\u0\/u2\/_0133_ ), .C1(\u0\/u2\/_0684_ ), .Y(\u0\/u2\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1458_ ( .A(\u0\/u2\/_0113_ ), .B(\u0\/u2\/_0251_ ), .Y(\u0\/u2\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u2/_1459_ ( .A_N(\u0\/u2\/_0463_ ), .B(\u0\/u2\/_0686_ ), .C(\u0\/u2\/_0383_ ), .D(\u0\/u2\/_0464_ ), .X(\u0\/u2\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1460_ ( .A1(\u0\/u2\/_0051_ ), .A2(\u0\/u2\/_0293_ ), .B1(\u0\/u2\/_0280_ ), .B2(\u0\/u2\/_0705_ ), .Y(\u0\/u2\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1461_ ( .A1(\u0\/u2\/_0017_ ), .A2(\u0\/u2\/_0072_ ), .B1(\u0\/u2\/_0456_ ), .B2(\u0\/u2\/_0078_ ), .Y(\u0\/u2\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1462_ ( .A(\u0\/u2\/_0687_ ), .B(\u0\/u2\/_0236_ ), .C(\u0\/u2\/_0688_ ), .D(\u0\/u2\/_0689_ ), .X(\u0\/u2\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1463_ ( .A(\u0\/u2\/_0680_ ), .B(\u0\/u2\/_0682_ ), .C(\u0\/u2\/_0685_ ), .D(\u0\/u2\/_0690_ ), .X(\u0\/u2\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u2/_1464_ ( .A1(\u0\/u2\/_0532_ ), .A2(\u0\/u2\/_0380_ ), .B1(\u0\/u2\/_0102_ ), .C1(\u0\/u2\/_0355_ ), .X(\u0\/u2\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u2/_1465_ ( .A(\u0\/u2\/_0692_ ), .B(\u0\/u2\/_0338_ ), .C(\u0\/u2\/_0644_ ), .Y(\u0\/u2\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1466_ ( .A(\u0\/u2\/_0016_ ), .B(\u0\/u2\/_0020_ ), .Y(\u0\/u2\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1467_ ( .A1(\u0\/u2\/_0032_ ), .A2(\u0\/u2\/_0137_ ), .B1(\u0\/u2\/_0279_ ), .B2(\u0\/u2\/_0094_ ), .Y(\u0\/u2\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1468_ ( .A1(\u0\/u2\/_0575_ ), .A2(\u0\/u2\/_0153_ ), .B1(\u0\/u2\/_0161_ ), .B2(\u0\/u2\/_0293_ ), .Y(\u0\/u2\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1469_ ( .A(\u0\/u2\/_0259_ ), .B(\u0\/u2\/_0695_ ), .C(\u0\/u2\/_0696_ ), .D(\u0\/u2\/_0697_ ), .X(\u0\/u2\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u2/_1470_ ( .A1(\u0\/u2\/_0255_ ), .A2(\u0\/u2\/_0640_ ), .B1(\u0\/u2\/_0016_ ), .B2(\u0\/u2\/_0193_ ), .X(\u0\/u2\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1471_ ( .A1(\u0\/u2\/_0060_ ), .A2(\u0\/u2\/_0176_ ), .B1(\u0\/u2\/_0699_ ), .C1(\u0\/u2\/_0177_ ), .Y(\u0\/u2\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1472_ ( .A1(\u0\/u2\/_0091_ ), .A2(\u0\/u2\/_0499_ ), .B1(\u0\/u2\/_0092_ ), .B2(\u0\/u2\/_0705_ ), .Y(\u0\/u2\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u2/_1473_ ( .A1(\u0\/u2\/_0705_ ), .A2(\u0\/u2\/_0683_ ), .B1(\u0\/u2\/_0093_ ), .B2(\u0\/u2\/_0114_ ), .Y(\u0\/u2\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u2/_1474_ ( .A1(\u0\/u2\/_0683_ ), .A2(\u0\/u2\/_0280_ ), .B1(\u0\/u2\/_0094_ ), .Y(\u0\/u2\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u2/_1475_ ( .A1(\u0\/u2\/_0543_ ), .A2(\u0\/u2\/_0216_ ), .B1(\u0\/u2\/_0038_ ), .C1(\u0\/u2\/_0056_ ), .Y(\u0\/u2\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1476_ ( .A(\u0\/u2\/_0701_ ), .B(\u0\/u2\/_0702_ ), .C(\u0\/u2\/_0703_ ), .D(\u0\/u2\/_0704_ ), .X(\u0\/u2\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1477_ ( .A(\u0\/u2\/_0693_ ), .B(\u0\/u2\/_0698_ ), .C(\u0\/u2\/_0700_ ), .D(\u0\/u2\/_0706_ ), .X(\u0\/u2\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u2/_1478_ ( .A1(\u0\/u2\/_0113_ ), .A2(\u0\/u2\/_0640_ ), .B1(\u0\/u2\/_0099_ ), .B2(\u0\/u2\/_0058_ ), .X(\u0\/u2\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u2/_1479_ ( .A(\u0\/u2\/_0407_ ), .B(\u0\/u2\/_0708_ ), .C(\u0\/u2\/_0529_ ), .Y(\u0\/u2\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1480_ ( .A(\u0\/u2\/_0568_ ), .B(\u0\/u2\/_0175_ ), .Y(\u0\/u2\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u2/_1481_ ( .A1(\u0\/u2\/_0247_ ), .A2(\u0\/u2\/_0114_ ), .A3(\u0\/u2\/_0051_ ), .B1(\u0\/u2\/_0130_ ), .Y(\u0\/u2\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1482_ ( .A(\u0\/u2\/_0709_ ), .B(\u0\/u2\/_0550_ ), .C(\u0\/u2\/_0710_ ), .D(\u0\/u2\/_0711_ ), .X(\u0\/u2\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u2/_1483_ ( .A1(\u0\/u2\/_0114_ ), .A2(\u0\/u2\/_0064_ ), .B1(\u0\/u2\/_0261_ ), .B2(\u0\/u2\/_0089_ ), .X(\u0\/u2\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1484_ ( .A1(\u0\/u2\/_0355_ ), .A2(\u0\/u2\/_0261_ ), .B1(\u0\/u2\/_0198_ ), .C1(\u0\/u2\/_0713_ ), .Y(\u0\/u2\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1485_ ( .A(\u0\/u2\/_0586_ ), .B(\u0\/u2\/_0478_ ), .Y(\u0\/u2\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u2/_1486_ ( .A_N(\u0\/u2\/_0541_ ), .B(\u0\/u2\/_0267_ ), .C(\u0\/u2\/_0715_ ), .D(\u0\/u2\/_0320_ ), .X(\u0\/u2\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1487_ ( .A(\u0\/u2\/_0586_ ), .B(\u0\/u2\/_0070_ ), .Y(\u0\/u2\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u2/_1488_ ( .A_N(\u0\/u2\/_0211_ ), .B(\u0\/u2\/_0155_ ), .C(\u0\/u2\/_0202_ ), .D(\u0\/u2\/_0718_ ), .X(\u0\/u2\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u2/_1489_ ( .A(\u0\/u2\/_0150_ ), .B(\u0\/u2\/_0216_ ), .C(\u0\/u2\/_0380_ ), .Y(\u0\/u2\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \u0/u2/_1490_ ( .A(\u0\/u2\/_0411_ ), .B(\u0\/u2\/_0720_ ), .X(\u0\/u2\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u2/_1491_ ( .A1(\u0\/u2\/_0017_ ), .A2(\u0\/u2\/_0022_ ), .B1(\u0\/u2\/_0078_ ), .X(\u0\/u2\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u2/_1492_ ( .A1(\u0\/u2\/_0456_ ), .A2(\u0\/u2\/_0738_ ), .B1(\u0\/u2\/_0101_ ), .C1(\u0\/u2\/_0722_ ), .Y(\u0\/u2\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1493_ ( .A(\u0\/u2\/_0717_ ), .B(\u0\/u2\/_0719_ ), .C(\u0\/u2\/_0721_ ), .D(\u0\/u2\/_0723_ ), .X(\u0\/u2\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u2/_1494_ ( .A(\u0\/u2\/_0739_ ), .B(\u0\/u2\/_0193_ ), .Y(\u0\/u2\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1495_ ( .A(\u0\/u2\/_0344_ ), .B(\u0\/u2\/_0184_ ), .C(\u0\/u2\/_0449_ ), .D(\u0\/u2\/_0725_ ), .X(\u0\/u2\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \u0/u2/_1496_ ( .A(\u0\/u2\/_0712_ ), .B(\u0\/u2\/_0714_ ), .C(\u0\/u2\/_0724_ ), .D(\u0\/u2\/_0726_ ), .X(\u0\/u2\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u2/_1497_ ( .A(\u0\/u2\/_0691_ ), .B(\u0\/u2\/_0707_ ), .C(\u0\/u2\/_0728_ ), .Y(\u0\/u2\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u3/_0753_ ( .A(\w3\[26\] ), .B_N(\w3\[27\] ), .Y(\u0\/u3\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_0755_ ( .A(\w3\[25\] ), .B(\w3\[24\] ), .X(\u0\/u3\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_0756_ ( .A(\u0\/u3\/_0096_ ), .B(\u0\/u3\/_0118_ ), .X(\u0\/u3\/_0129_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0757_ ( .A(\u0\/u3\/_0007_ ), .B(\w3\[30\] ), .X(\u0\/u3\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_0758_ ( .A(\w3\[28\] ), .B(\w3\[29\] ), .Y(\u0\/u3\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0759_ ( .A(\u0\/u3\/_0140_ ), .B(\u0\/u3\/_0151_ ), .X(\u0\/u3\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0761_ ( .A(\u0\/u3\/_0129_ ), .B(\u0\/u3\/_0162_ ), .X(\u0\/u3\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0762_ ( .A(\u0\/u3\/_0096_ ), .X(\u0\/u3\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u3/_0763_ ( .A(\w3\[25\] ), .B_N(\w3\[24\] ), .Y(\u0\/u3\/_0205_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0764_ ( .A(\u0\/u3\/_0205_ ), .X(\u0\/u3\/_0216_ ) );
sky130_fd_sc_hd__and3_1 \u0/u3/_0765_ ( .A(\u0\/u3\/_0162_ ), .B(\u0\/u3\/_0194_ ), .C(\u0\/u3\/_0216_ ), .X(\u0\/u3\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \u0/u3/_0766_ ( .A(\u0\/u3\/_0183_ ), .SLEEP(\u0\/u3\/_0227_ ), .X(\u0\/u3\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u3/_0767_ ( .A(\w3\[24\] ), .B_N(\w3\[25\] ), .Y(\u0\/u3\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_0768_ ( .A(\w3\[26\] ), .B(\w3\[27\] ), .Y(\u0\/u3\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0769_ ( .A(\u0\/u3\/_0249_ ), .B(\u0\/u3\/_0260_ ), .X(\u0\/u3\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0771_ ( .A(\u0\/u3\/_0271_ ), .X(\u0\/u3\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0772_ ( .A(\u0\/u3\/_0162_ ), .X(\u0\/u3\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_0773_ ( .A(\u0\/u3\/_0293_ ), .B(\u0\/u3\/_0304_ ), .Y(\u0\/u3\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \u0/u3/_0774_ ( .A(\w3\[25\] ), .Y(\u0\/u3\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \u0/u3/_0776_ ( .A(\w3\[24\] ), .Y(\u0\/u3\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0777_ ( .A(\w3\[26\] ), .B(\w3\[27\] ), .X(\u0\/u3\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0779_ ( .A(\u0\/u3\/_0358_ ), .X(\u0\/u3\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_0780_ ( .A1(\u0\/u3\/_0325_ ), .A2(\u0\/u3\/_0347_ ), .B1(\u0\/u3\/_0380_ ), .C1(\u0\/u3\/_0304_ ), .Y(\u0\/u3\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u3/_0781_ ( .A_N(\u0\/u3\/_0238_ ), .B(\u0\/u3\/_0314_ ), .C(\u0\/u3\/_0391_ ), .X(\u0\/u3\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u3/_0782_ ( .A(\w3\[27\] ), .B_N(\w3\[26\] ), .Y(\u0\/u3\/_0412_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0784_ ( .A(\u0\/u3\/_0412_ ), .B(\u0\/u3\/_0205_ ), .X(\u0\/u3\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u3/_0787_ ( .A(\w3\[29\] ), .B_N(\w3\[28\] ), .Y(\u0\/u3\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0788_ ( .A(\u0\/u3\/_0467_ ), .B(\u0\/u3\/_0140_ ), .X(\u0\/u3\/_0478_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_0791_ ( .A(\u0\/u3\/_0134_ ), .B(\u0\/u3\/_0218_ ), .Y(\u0\/u3\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_0792_ ( .A(\u0\/u3\/_0478_ ), .B(\u0\/u3\/_0271_ ), .Y(\u0\/u3\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0793_ ( .A(\u0\/u3\/_0194_ ), .X(\u0\/u3\/_0532_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_0795_ ( .A(\u0\/u3\/_0249_ ), .B(\u0\/u3\/_0358_ ), .X(\u0\/u3\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0797_ ( .A(\u0\/u3\/_0554_ ), .X(\u0\/u3\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_0798_ ( .A(\u0\/u3\/_0216_ ), .B(\u0\/u3\/_0358_ ), .X(\u0\/u3\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0800_ ( .A(\u0\/u3\/_0586_ ), .X(\u0\/u3\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_0801_ ( .A1(\u0\/u3\/_0532_ ), .A2(\u0\/u3\/_0575_ ), .A3(\u0\/u3\/_0608_ ), .B1(\u0\/u3\/_0218_ ), .Y(\u0\/u3\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_0802_ ( .A(\u0\/u3\/_0401_ ), .B(\u0\/u3\/_0510_ ), .C(\u0\/u3\/_0521_ ), .D(\u0\/u3\/_0619_ ), .X(\u0\/u3\/_0629_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0803_ ( .A(\u0\/u3\/_0358_ ), .B(\w3\[25\] ), .X(\u0\/u3\/_0640_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_0805_ ( .A(\u0\/u3\/_0205_ ), .B(\u0\/u3\/_0260_ ), .X(\u0\/u3\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0807_ ( .A(\u0\/u3\/_0662_ ), .X(\u0\/u3\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u3/_0808_ ( .A(\w3\[30\] ), .B_N(\u0\/u3\/_0007_ ), .Y(\u0\/u3\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_0809_ ( .A(\u0\/u3\/_0467_ ), .B(\u0\/u3\/_0694_ ), .X(\u0\/u3\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0811_ ( .A(\u0\/u3\/_0705_ ), .X(\u0\/u3\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_0812_ ( .A1(\u0\/u3\/_0640_ ), .A2(\u0\/u3\/_0293_ ), .A3(\u0\/u3\/_0683_ ), .B1(\u0\/u3\/_0727_ ), .Y(\u0\/u3\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_0813_ ( .A(\w3\[25\] ), .B(\w3\[24\] ), .Y(\u0\/u3\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0814_ ( .A(\u0\/u3\/_0730_ ), .B(\u0\/u3\/_0260_ ), .X(\u0\/u3\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0816_ ( .A(\u0\/u3\/_0731_ ), .X(\u0\/u3\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0817_ ( .A(\w3\[24\] ), .X(\u0\/u3\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u3/_0818_ ( .A1(\u0\/u3\/_0325_ ), .A2(\u0\/u3\/_0734_ ), .B1(\u0\/u3\/_0412_ ), .X(\u0\/u3\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0819_ ( .A(\u0\/u3\/_0694_ ), .B(\u0\/u3\/_0151_ ), .X(\u0\/u3\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0821_ ( .A(\u0\/u3\/_0736_ ), .X(\u0\/u3\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0822_ ( .A(\u0\/u3\/_0738_ ), .X(\u0\/u3\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_0823_ ( .A1(\u0\/u3\/_0733_ ), .A2(\u0\/u3\/_0735_ ), .A3(\u0\/u3\/_0293_ ), .B1(\u0\/u3\/_0739_ ), .Y(\u0\/u3\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u3/_0824_ ( .A(\u0\/u3\/_0730_ ), .B_N(\u0\/u3\/_0358_ ), .Y(\u0\/u3\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_0825_ ( .A(\u0\/u3\/_0741_ ), .B(\u0\/u3\/_0739_ ), .Y(\u0\/u3\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_0827_ ( .A1(\u0\/u3\/_0118_ ), .A2(\u0\/u3\/_0216_ ), .B1(\u0\/u3\/_0532_ ), .C1(\u0\/u3\/_0739_ ), .Y(\u0\/u3\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_0828_ ( .A(\u0\/u3\/_0729_ ), .B(\u0\/u3\/_0740_ ), .C(\u0\/u3\/_0742_ ), .D(\u0\/u3\/_0744_ ), .X(\u0\/u3\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0829_ ( .A(\u0\/u3\/_0412_ ), .B(\u0\/u3\/_0730_ ), .X(\u0\/u3\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0831_ ( .A(\u0\/u3\/_0746_ ), .X(\u0\/u3\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u3/_0832_ ( .A(\w3\[28\] ), .B_N(\w3\[29\] ), .Y(\u0\/u3\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0833_ ( .A(\u0\/u3\/_0749_ ), .B(\u0\/u3\/_0694_ ), .X(\u0\/u3\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0835_ ( .A(\u0\/u3\/_0750_ ), .X(\u0\/u3\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0836_ ( .A(\u0\/u3\/_0752_ ), .X(\u0\/u3\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0837_ ( .A(\u0\/u3\/_0118_ ), .B(\u0\/u3\/_0358_ ), .X(\u0\/u3\/_0017_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0839_ ( .A(\u0\/u3\/_0752_ ), .B(\u0\/u3\/_0017_ ), .X(\u0\/u3\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0840_ ( .A(\u0\/u3\/_0358_ ), .B(\u0\/u3\/_0325_ ), .X(\u0\/u3\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0842_ ( .A(\u0\/u3\/_0096_ ), .B(\u0\/u3\/_0205_ ), .X(\u0\/u3\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u3/_0844_ ( .A1(\u0\/u3\/_0020_ ), .A2(\u0\/u3\/_0022_ ), .B1(\u0\/u3\/_0752_ ), .X(\u0\/u3\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_0845_ ( .A1(\u0\/u3\/_0748_ ), .A2(\u0\/u3\/_0016_ ), .B1(\u0\/u3\/_0019_ ), .C1(\u0\/u3\/_0024_ ), .Y(\u0\/u3\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_0846_ ( .A(\w3\[28\] ), .B(\w3\[29\] ), .X(\u0\/u3\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0847_ ( .A(\u0\/u3\/_0694_ ), .B(\u0\/u3\/_0026_ ), .X(\u0\/u3\/_0027_ ) );
sky130_fd_sc_hd__buf_2 \u0/u3/_0849_ ( .A(\u0\/u3\/_0027_ ), .X(\u0\/u3\/_0029_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0850_ ( .A(\u0\/u3\/_0358_ ), .B(\u0\/u3\/_0730_ ), .X(\u0\/u3\/_0030_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0852_ ( .A(\u0\/u3\/_0030_ ), .X(\u0\/u3\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_0853_ ( .A(\u0\/u3\/_0029_ ), .B(\u0\/u3\/_0032_ ), .Y(\u0\/u3\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_0854_ ( .A(\u0\/u3\/_0029_ ), .B(\u0\/u3\/_0735_ ), .Y(\u0\/u3\/_0034_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_0855_ ( .A(\u0\/u3\/_0118_ ), .B(\u0\/u3\/_0260_ ), .X(\u0\/u3\/_0035_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0857_ ( .A(\u0\/u3\/_0027_ ), .B(\u0\/u3\/_0035_ ), .X(\u0\/u3\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0858_ ( .A(\u0\/u3\/_0260_ ), .X(\u0\/u3\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_0859_ ( .A(\u0\/u3\/_0038_ ), .B(\u0\/u3\/_0347_ ), .Y(\u0\/u3\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u3/_0860_ ( .A_N(\u0\/u3\/_0039_ ), .B(\u0\/u3\/_0027_ ), .X(\u0\/u3\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_0861_ ( .A(\u0\/u3\/_0037_ ), .B(\u0\/u3\/_0040_ ), .Y(\u0\/u3\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_0862_ ( .A(\u0\/u3\/_0025_ ), .B(\u0\/u3\/_0033_ ), .C(\u0\/u3\/_0034_ ), .D(\u0\/u3\/_0041_ ), .X(\u0\/u3\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0863_ ( .A(\u0\/u3\/_0749_ ), .B(\u0\/u3\/_0140_ ), .X(\u0\/u3\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \u0/u3/_0865_ ( .A(\w3\[24\] ), .B(\w3\[26\] ), .C(\w3\[27\] ), .X(\u0\/u3\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0866_ ( .A(\u0\/u3\/_0043_ ), .B(\u0\/u3\/_0045_ ), .X(\u0\/u3\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0867_ ( .A(\u0\/u3\/_0096_ ), .B(\u0\/u3\/_0249_ ), .X(\u0\/u3\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0869_ ( .A(\u0\/u3\/_0047_ ), .B(\u0\/u3\/_0043_ ), .X(\u0\/u3\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0870_ ( .A(\u0\/u3\/_0730_ ), .X(\u0\/u3\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0871_ ( .A(\u0\/u3\/_0043_ ), .X(\u0\/u3\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_0872_ ( .A1(\u0\/u3\/_0118_ ), .A2(\u0\/u3\/_0050_ ), .B1(\u0\/u3\/_0194_ ), .C1(\u0\/u3\/_0051_ ), .Y(\u0\/u3\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u3/_0873_ ( .A(\u0\/u3\/_0046_ ), .B(\u0\/u3\/_0049_ ), .C_N(\u0\/u3\/_0052_ ), .Y(\u0\/u3\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0874_ ( .A(\u0\/u3\/_0026_ ), .B(\u0\/u3\/_0140_ ), .X(\u0\/u3\/_0054_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_0877_ ( .A1(\u0\/u3\/_0532_ ), .A2(\u0\/u3\/_0575_ ), .B1(\u0\/u3\/_0292_ ), .Y(\u0\/u3\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0878_ ( .A(\u0\/u3\/_0412_ ), .B(\u0\/u3\/_0325_ ), .X(\u0\/u3\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0880_ ( .A(\u0\/u3\/_0051_ ), .X(\u0\/u3\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_0881_ ( .A1(\u0\/u3\/_0731_ ), .A2(\u0\/u3\/_0035_ ), .A3(\u0\/u3\/_0058_ ), .B1(\u0\/u3\/_0060_ ), .Y(\u0\/u3\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0882_ ( .A(\u0\/u3\/_0260_ ), .B(\w3\[25\] ), .X(\u0\/u3\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0884_ ( .A(\u0\/u3\/_0062_ ), .X(\u0\/u3\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_0885_ ( .A1(\u0\/u3\/_0064_ ), .A2(\u0\/u3\/_0748_ ), .A3(\u0\/u3\/_0683_ ), .B1(\u0\/u3\/_0292_ ), .Y(\u0\/u3\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_0886_ ( .A(\u0\/u3\/_0053_ ), .B(\u0\/u3\/_0057_ ), .C(\u0\/u3\/_0061_ ), .D(\u0\/u3\/_0065_ ), .X(\u0\/u3\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_0887_ ( .A(\u0\/u3\/_0629_ ), .B(\u0\/u3\/_0745_ ), .C(\u0\/u3\/_0042_ ), .D(\u0\/u3\/_0066_ ), .X(\u0\/u3\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u3/_0889_ ( .A(\u0\/u3\/_0007_ ), .B_N(\w3\[30\] ), .Y(\u0\/u3\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0890_ ( .A(\u0\/u3\/_0069_ ), .B(\u0\/u3\/_0151_ ), .X(\u0\/u3\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0892_ ( .A(\u0\/u3\/_0070_ ), .X(\u0\/u3\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_0893_ ( .A1(\u0\/u3\/_0129_ ), .A2(\u0\/u3\/_0586_ ), .B1(\u0\/u3\/_0072_ ), .Y(\u0\/u3\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_0894_ ( .A1(\u0\/u3\/_0380_ ), .A2(\u0\/u3\/_0347_ ), .B1(\u0\/u3\/_0194_ ), .B2(\u0\/u3\/_0216_ ), .Y(\u0\/u3\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u3/_0895_ ( .A(\u0\/u3\/_0074_ ), .B_N(\u0\/u3\/_0070_ ), .Y(\u0\/u3\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u3/_0896_ ( .A(\u0\/u3\/_0073_ ), .SLEEP(\u0\/u3\/_0075_ ), .X(\u0\/u3\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_0897_ ( .A(\u0\/u3\/_0467_ ), .B(\u0\/u3\/_0069_ ), .X(\u0\/u3\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0898_ ( .A(\u0\/u3\/_0077_ ), .X(\u0\/u3\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0899_ ( .A(\u0\/u3\/_0412_ ), .B(\u0\/u3\/_0118_ ), .X(\u0\/u3\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0901_ ( .A(\u0\/u3\/_0078_ ), .B(\u0\/u3\/_0079_ ), .X(\u0\/u3\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0902_ ( .A(\u0\/u3\/_0412_ ), .B(\u0\/u3\/_0249_ ), .X(\u0\/u3\/_0082_ ) );
sky130_fd_sc_hd__buf_2 \u0/u3/_0904_ ( .A(\u0\/u3\/_0082_ ), .X(\u0\/u3\/_0084_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0905_ ( .A(\u0\/u3\/_0084_ ), .B(\u0\/u3\/_0078_ ), .X(\u0\/u3\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u3/_0906_ ( .A1(\w3\[24\] ), .A2(\u0\/u3\/_0325_ ), .B1(\u0\/u3\/_0260_ ), .Y(\u0\/u3\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u3/_0907_ ( .A_N(\u0\/u3\/_0086_ ), .B(\u0\/u3\/_0078_ ), .X(\u0\/u3\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u3/_0908_ ( .A(\u0\/u3\/_0081_ ), .B(\u0\/u3\/_0085_ ), .C(\u0\/u3\/_0087_ ), .Y(\u0\/u3\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0909_ ( .A(\u0\/u3\/_0072_ ), .X(\u0\/u3\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_0910_ ( .A1(\u0\/u3\/_0733_ ), .A2(\u0\/u3\/_0748_ ), .A3(\u0\/u3\/_0683_ ), .B1(\u0\/u3\/_0089_ ), .Y(\u0\/u3\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0911_ ( .A(\u0\/u3\/_0129_ ), .X(\u0\/u3\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0912_ ( .A(\u0\/u3\/_0017_ ), .X(\u0\/u3\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0913_ ( .A(\u0\/u3\/_0022_ ), .X(\u0\/u3\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0914_ ( .A(\u0\/u3\/_0078_ ), .X(\u0\/u3\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_0915_ ( .A1(\u0\/u3\/_0091_ ), .A2(\u0\/u3\/_0092_ ), .A3(\u0\/u3\/_0093_ ), .B1(\u0\/u3\/_0094_ ), .Y(\u0\/u3\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_0916_ ( .A(\u0\/u3\/_0076_ ), .B(\u0\/u3\/_0088_ ), .C(\u0\/u3\/_0090_ ), .D(\u0\/u3\/_0095_ ), .X(\u0\/u3\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_0917_ ( .A(\u0\/u3\/_0069_ ), .B(\u0\/u3\/_0026_ ), .X(\u0\/u3\/_0098_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0919_ ( .A(\u0\/u3\/_0434_ ), .B(\u0\/u3\/_0364_ ), .X(\u0\/u3\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0920_ ( .A(\u0\/u3\/_0079_ ), .B(\u0\/u3\/_0098_ ), .X(\u0\/u3\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0921_ ( .A(\u0\/u3\/_0325_ ), .X(\u0\/u3\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_0922_ ( .A1(\u0\/u3\/_0102_ ), .A2(\u0\/u3\/_0734_ ), .B1(\u0\/u3\/_0038_ ), .C1(\u0\/u3\/_0364_ ), .Y(\u0\/u3\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u3/_0923_ ( .A(\u0\/u3\/_0100_ ), .B(\u0\/u3\/_0101_ ), .C_N(\u0\/u3\/_0103_ ), .Y(\u0\/u3\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_0924_ ( .A1(\u0\/u3\/_0554_ ), .A2(\u0\/u3\/_0586_ ), .B1(\u0\/u3\/_0364_ ), .Y(\u0\/u3\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_0925_ ( .A(\u0\/u3\/_0129_ ), .B(\u0\/u3\/_0364_ ), .Y(\u0\/u3\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0926_ ( .A(\u0\/u3\/_0105_ ), .B(\u0\/u3\/_0106_ ), .X(\u0\/u3\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0927_ ( .A(\u0\/u3\/_0412_ ), .X(\u0\/u3\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_0928_ ( .A(\u0\/u3\/_0260_ ), .B(\w3\[24\] ), .X(\u0\/u3\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0929_ ( .A(\u0\/u3\/_0069_ ), .B(\u0\/u3\/_0749_ ), .X(\u0\/u3\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0931_ ( .A(\u0\/u3\/_0111_ ), .X(\u0\/u3\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0932_ ( .A(\u0\/u3\/_0113_ ), .X(\u0\/u3\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_0933_ ( .A1(\u0\/u3\/_0109_ ), .A2(\u0\/u3\/_0110_ ), .B1(\u0\/u3\/_0114_ ), .Y(\u0\/u3\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_0934_ ( .A(\u0\/u3\/_0022_ ), .Y(\u0\/u3\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_0935_ ( .A(\u0\/u3\/_0554_ ), .Y(\u0\/u3\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u3/_0936_ ( .A1(\u0\/u3\/_0050_ ), .A2(\u0\/u3\/_0118_ ), .B1(\u0\/u3\/_0194_ ), .Y(\u0\/u3\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_0937_ ( .A(\u0\/u3\/_0113_ ), .Y(\u0\/u3\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \u0/u3/_0938_ ( .A1(\u0\/u3\/_0116_ ), .A2(\u0\/u3\/_0117_ ), .A3(\u0\/u3\/_0119_ ), .B1(\u0\/u3\/_0120_ ), .X(\u0\/u3\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_0939_ ( .A(\u0\/u3\/_0104_ ), .B(\u0\/u3\/_0108_ ), .C(\u0\/u3\/_0115_ ), .D(\u0\/u3\/_0121_ ), .X(\u0\/u3\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_0940_ ( .A(\u0\/u3\/_0007_ ), .B(\w3\[30\] ), .Y(\u0\/u3\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0941_ ( .A(\u0\/u3\/_0749_ ), .B(\u0\/u3\/_0123_ ), .X(\u0\/u3\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0943_ ( .A(\u0\/u3\/_0082_ ), .B(\u0\/u3\/_0124_ ), .X(\u0\/u3\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_0944_ ( .A(\u0\/u3\/_0271_ ), .B(\u0\/u3\/_0124_ ), .Y(\u0\/u3\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0945_ ( .A(\u0\/u3\/_0124_ ), .X(\u0\/u3\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0946_ ( .A(\u0\/u3\/_0260_ ), .B(\u0\/u3\/_0325_ ), .X(\u0\/u3\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_0948_ ( .A(\u0\/u3\/_0128_ ), .B(\u0\/u3\/_0130_ ), .Y(\u0\/u3\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_0949_ ( .A(\u0\/u3\/_0127_ ), .B(\u0\/u3\/_0132_ ), .Y(\u0\/u3\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \u0/u3/_0950_ ( .A(\u0\/u3\/_0434_ ), .X(\u0\/u3\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_0951_ ( .A(\u0\/u3\/_0134_ ), .B(\u0\/u3\/_0128_ ), .Y(\u0\/u3\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u3/_0952_ ( .A(\u0\/u3\/_0126_ ), .B(\u0\/u3\/_0133_ ), .C_N(\u0\/u3\/_0135_ ), .Y(\u0\/u3\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_0953_ ( .A(\u0\/u3\/_0026_ ), .B(\u0\/u3\/_0123_ ), .X(\u0\/u3\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0955_ ( .A(\u0\/u3\/_0137_ ), .X(\u0\/u3\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_0956_ ( .A1(\u0\/u3\/_0110_ ), .A2(\u0\/u3\/_0293_ ), .A3(\u0\/u3\/_0084_ ), .B1(\u0\/u3\/_0139_ ), .Y(\u0\/u3\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0957_ ( .A(\u0\/u3\/_0096_ ), .B(\u0\/u3\/_0730_ ), .X(\u0\/u3\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0959_ ( .A(\u0\/u3\/_0142_ ), .X(\u0\/u3\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_0960_ ( .A1(\u0\/u3\/_0020_ ), .A2(\u0\/u3\/_0144_ ), .A3(\u0\/u3\/_0017_ ), .B1(\u0\/u3\/_0139_ ), .Y(\u0\/u3\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u3/_0961_ ( .A(\w3\[26\] ), .B(\u0\/u3\/_0050_ ), .C_N(\w3\[27\] ), .Y(\u0\/u3\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0962_ ( .A(\u0\/u3\/_0128_ ), .X(\u0\/u3\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_0963_ ( .A1(\u0\/u3\/_0146_ ), .A2(\u0\/u3\/_0032_ ), .A3(\u0\/u3\/_0640_ ), .B1(\u0\/u3\/_0147_ ), .Y(\u0\/u3\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_0964_ ( .A(\u0\/u3\/_0136_ ), .B(\u0\/u3\/_0141_ ), .C(\u0\/u3\/_0145_ ), .D(\u0\/u3\/_0148_ ), .X(\u0\/u3\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0965_ ( .A(\u0\/u3\/_0123_ ), .B(\u0\/u3\/_0151_ ), .X(\u0\/u3\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0967_ ( .A(\u0\/u3\/_0150_ ), .X(\u0\/u3\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_0968_ ( .A(\u0\/u3\/_0150_ ), .B(\u0\/u3\/_0062_ ), .X(\u0\/u3\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_0969_ ( .A(\u0\/u3\/_0079_ ), .B(\u0\/u3\/_0150_ ), .Y(\u0\/u3\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u3/_0970_ ( .A(\u0\/u3\/_0150_ ), .B(\u0\/u3\/_0412_ ), .C(\u0\/u3\/_0249_ ), .Y(\u0\/u3\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_0971_ ( .A(\u0\/u3\/_0155_ ), .B(\u0\/u3\/_0156_ ), .Y(\u0\/u3\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_0972_ ( .A1(\u0\/u3\/_0153_ ), .A2(\u0\/u3\/_0134_ ), .B1(\u0\/u3\/_0154_ ), .C1(\u0\/u3\/_0157_ ), .Y(\u0\/u3\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0973_ ( .A(\u0\/u3\/_0467_ ), .B(\u0\/u3\/_0123_ ), .X(\u0\/u3\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_0975_ ( .A(\u0\/u3\/_0159_ ), .X(\u0\/u3\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u3/_0976_ ( .A_N(\u0\/u3\/_0119_ ), .B(\u0\/u3\/_0161_ ), .X(\u0\/u3\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_0977_ ( .A(\u0\/u3\/_0163_ ), .Y(\u0\/u3\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_0978_ ( .A1(\u0\/u3\/_0146_ ), .A2(\u0\/u3\/_0575_ ), .A3(\u0\/u3\/_0608_ ), .B1(\u0\/u3\/_0153_ ), .Y(\u0\/u3\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_0979_ ( .A1(\u0\/u3\/_0062_ ), .A2(\u0\/u3\/_0084_ ), .A3(\u0\/u3\/_0134_ ), .B1(\u0\/u3\/_0161_ ), .Y(\u0\/u3\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_0980_ ( .A(\u0\/u3\/_0158_ ), .B(\u0\/u3\/_0164_ ), .C(\u0\/u3\/_0165_ ), .D(\u0\/u3\/_0166_ ), .X(\u0\/u3\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_0981_ ( .A(\u0\/u3\/_0097_ ), .B(\u0\/u3\/_0122_ ), .C(\u0\/u3\/_0149_ ), .D(\u0\/u3\/_0167_ ), .X(\u0\/u3\/_0168_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0982_ ( .A(\u0\/u3\/_0662_ ), .B(\u0\/u3\/_0150_ ), .X(\u0\/u3\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_0983_ ( .A(\u0\/u3\/_0154_ ), .B(\u0\/u3\/_0169_ ), .Y(\u0\/u3\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \u0/u3/_0984_ ( .A(\u0\/u3\/_0123_ ), .B(\u0\/u3\/_0151_ ), .C(\u0\/u3\/_0038_ ), .X(\u0\/u3\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0985_ ( .A(\u0\/u3\/_0170_ ), .B(\u0\/u3\/_0171_ ), .X(\u0\/u3\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_0986_ ( .A(\u0\/u3\/_0172_ ), .Y(\u0\/u3\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u3/_0987_ ( .A(\u0\/u3\/_0067_ ), .B(\u0\/u3\/_0168_ ), .C(\u0\/u3\/_0174_ ), .Y(\u0\/u3\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \u0/u3/_0988_ ( .A(\w3\[25\] ), .B(\w3\[24\] ), .Y(\u0\/u3\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_0989_ ( .A(\u0\/u3\/_0175_ ), .B(\u0\/u3\/_0358_ ), .X(\u0\/u3\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0990_ ( .A(\u0\/u3\/_0176_ ), .B(\u0\/u3\/_0478_ ), .X(\u0\/u3\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_0991_ ( .A(\u0\/u3\/_0084_ ), .B(\u0\/u3\/_0113_ ), .Y(\u0\/u3\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0992_ ( .A(\u0\/u3\/_0111_ ), .B(\u0\/u3\/_0062_ ), .X(\u0\/u3\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0993_ ( .A(\u0\/u3\/_0111_ ), .B(\u0\/u3\/_0662_ ), .X(\u0\/u3\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_0994_ ( .A(\u0\/u3\/_0179_ ), .B(\u0\/u3\/_0180_ ), .Y(\u0\/u3\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0995_ ( .A(\u0\/u3\/_0054_ ), .B(\u0\/u3\/_0058_ ), .X(\u0\/u3\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_0996_ ( .A(\u0\/u3\/_0182_ ), .Y(\u0\/u3\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u3/_0997_ ( .A_N(\u0\/u3\/_0177_ ), .B(\u0\/u3\/_0178_ ), .C(\u0\/u3\/_0181_ ), .D(\u0\/u3\/_0184_ ), .X(\u0\/u3\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0998_ ( .A(\u0\/u3\/_0098_ ), .B(\u0\/u3\/_0741_ ), .X(\u0\/u3\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_0999_ ( .A(\u0\/u3\/_0047_ ), .B(\u0\/u3\/_0098_ ), .X(\u0\/u3\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \u0/u3/_1000_ ( .A(\u0\/u3\/_0186_ ), .B(\u0\/u3\/_0187_ ), .X(\u0\/u3\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1001_ ( .A(\u0\/u3\/_0188_ ), .Y(\u0\/u3\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1002_ ( .A(\u0\/u3\/_0738_ ), .B(\u0\/u3\/_0735_ ), .X(\u0\/u3\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1003_ ( .A(\u0\/u3\/_0271_ ), .B(\u0\/u3\/_0736_ ), .X(\u0\/u3\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_1004_ ( .A(\u0\/u3\/_0190_ ), .B(\u0\/u3\/_0191_ ), .Y(\u0\/u3\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_1005_ ( .A(\u0\/u3\/_0096_ ), .B(\u0\/u3\/_0325_ ), .X(\u0\/u3\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1006_ ( .A1(\u0\/u3\/_0193_ ), .A2(\u0\/u3\/_0176_ ), .B1(\u0\/u3\/_0043_ ), .Y(\u0\/u3\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1007_ ( .A(\u0\/u3\/_0185_ ), .B(\u0\/u3\/_0189_ ), .C(\u0\/u3\/_0192_ ), .D(\u0\/u3\/_0195_ ), .X(\u0\/u3\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u3/_1008_ ( .A_N(\w3\[27\] ), .B(\u0\/u3\/_0734_ ), .C(\w3\[26\] ), .X(\u0\/u3\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1009_ ( .A(\u0\/u3\/_0137_ ), .B(\u0\/u3\/_0197_ ), .X(\u0\/u3\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_1010_ ( .A(\u0\/u3\/_0198_ ), .B(\u0\/u3\/_0040_ ), .Y(\u0\/u3\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1011_ ( .A(\u0\/u3\/_0293_ ), .B(\u0\/u3\/_0137_ ), .X(\u0\/u3\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1012_ ( .A(\u0\/u3\/_0200_ ), .Y(\u0\/u3\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1013_ ( .A(\u0\/u3\/_0137_ ), .B(\u0\/u3\/_0110_ ), .Y(\u0\/u3\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1014_ ( .A(\u0\/u3\/_0139_ ), .B(\u0\/u3\/_0020_ ), .Y(\u0\/u3\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1015_ ( .A(\u0\/u3\/_0199_ ), .B(\u0\/u3\/_0201_ ), .C(\u0\/u3\/_0202_ ), .D(\u0\/u3\/_0203_ ), .X(\u0\/u3\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u3/_1016_ ( .A1(\u0\/u3\/_0532_ ), .A2(\u0\/u3\/_0109_ ), .B1(\u0\/u3\/_0102_ ), .C1(\u0\/u3\/_0727_ ), .X(\u0\/u3\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1017_ ( .A(\u0\/u3\/_0022_ ), .B(\u0\/u3\/_0078_ ), .Y(\u0\/u3\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1018_ ( .A(\u0\/u3\/_0078_ ), .B(\u0\/u3\/_0142_ ), .Y(\u0\/u3\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1019_ ( .A(\u0\/u3\/_0207_ ), .B(\u0\/u3\/_0208_ ), .Y(\u0\/u3\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1020_ ( .A1(\u0\/u3\/_0094_ ), .A2(\u0\/u3\/_0176_ ), .B1(\u0\/u3\/_0206_ ), .C1(\u0\/u3\/_0209_ ), .Y(\u0\/u3\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1021_ ( .A(\u0\/u3\/_0662_ ), .B(\u0\/u3\/_0070_ ), .X(\u0\/u3\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u3/_1022_ ( .A(\u0\/u3\/_0731_ ), .B(\u0\/u3\/_0123_ ), .C(\u0\/u3\/_0749_ ), .Y(\u0\/u3\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u3/_1023_ ( .A(\u0\/u3\/_0731_ ), .B(\u0\/u3\/_0467_ ), .C(\u0\/u3\/_0069_ ), .Y(\u0\/u3\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u3/_1024_ ( .A_N(\u0\/u3\/_0211_ ), .B(\u0\/u3\/_0127_ ), .C(\u0\/u3\/_0212_ ), .D(\u0\/u3\/_0213_ ), .X(\u0\/u3\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1025_ ( .A(\u0\/u3\/_0137_ ), .Y(\u0\/u3\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1026_ ( .A(\u0\/u3\/_0128_ ), .B(\u0\/u3\/_0035_ ), .Y(\u0\/u3\/_0217_ ) );
sky130_fd_sc_hd__buf_2 \u0/u3/_1027_ ( .A(\u0\/u3\/_0478_ ), .X(\u0\/u3\/_0218_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1028_ ( .A1(\u0\/u3\/_0159_ ), .A2(\u0\/u3\/_0746_ ), .B1(\u0\/u3\/_0434_ ), .B2(\u0\/u3\/_0218_ ), .Y(\u0\/u3\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u3/_1029_ ( .A1(\u0\/u3\/_0116_ ), .A2(\u0\/u3\/_0215_ ), .B1(\u0\/u3\/_0217_ ), .C1(\u0\/u3\/_0219_ ), .X(\u0\/u3\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1030_ ( .A(\u0\/u3\/_0113_ ), .B(\u0\/u3\/_0746_ ), .X(\u0\/u3\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u3/_1031_ ( .A1(\u0\/u3\/_0098_ ), .A2(\u0\/u3\/_0746_ ), .B1(\u0\/u3\/_0434_ ), .B2(\u0\/u3\/_0750_ ), .X(\u0\/u3\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1032_ ( .A1(\u0\/u3\/_0047_ ), .A2(\u0\/u3\/_0113_ ), .B1(\u0\/u3\/_0221_ ), .C1(\u0\/u3\/_0222_ ), .Y(\u0\/u3\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u3/_1033_ ( .A1(\u0\/u3\/_0129_ ), .A2(\u0\/u3\/_0162_ ), .B1(\u0\/u3\/_0271_ ), .B2(\u0\/u3\/_0705_ ), .X(\u0\/u3\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1034_ ( .A1(\u0\/u3\/_0093_ ), .A2(\u0\/u3\/_0738_ ), .B1(\u0\/u3\/_0081_ ), .C1(\u0\/u3\/_0224_ ), .Y(\u0\/u3\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1035_ ( .A(\u0\/u3\/_0214_ ), .B(\u0\/u3\/_0220_ ), .C(\u0\/u3\/_0223_ ), .D(\u0\/u3\/_0225_ ), .X(\u0\/u3\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1036_ ( .A(\u0\/u3\/_0196_ ), .B(\u0\/u3\/_0204_ ), .C(\u0\/u3\/_0210_ ), .D(\u0\/u3\/_0226_ ), .X(\u0\/u3\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1037_ ( .A(\u0\/u3\/_0111_ ), .B(\u0\/u3\/_0554_ ), .X(\u0\/u3\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1038_ ( .A(\u0\/u3\/_0229_ ), .Y(\u0\/u3\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1039_ ( .A(\u0\/u3\/_0111_ ), .B(\u0\/u3\/_0129_ ), .Y(\u0\/u3\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1040_ ( .A(\u0\/u3\/_0017_ ), .B(\u0\/u3\/_0738_ ), .Y(\u0\/u3\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1041_ ( .A(\u0\/u3\/_0030_ ), .B(\u0\/u3\/_0304_ ), .Y(\u0\/u3\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1042_ ( .A(\u0\/u3\/_0230_ ), .B(\u0\/u3\/_0231_ ), .C(\u0\/u3\/_0232_ ), .D(\u0\/u3\/_0233_ ), .X(\u0\/u3\/_0234_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1043_ ( .A(\u0\/u3\/_0047_ ), .B(\u0\/u3\/_0478_ ), .X(\u0\/u3\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1044_ ( .A1(\u0\/u3\/_0129_ ), .A2(\u0\/u3\/_0554_ ), .B1(\u0\/u3\/_0137_ ), .Y(\u0\/u3\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u3/_1045_ ( .A(\u0\/u3\/_0235_ ), .B(\u0\/u3\/_0049_ ), .C_N(\u0\/u3\/_0236_ ), .Y(\u0\/u3\/_0237_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_1046_ ( .A(\u0\/u3\/_0047_ ), .B(\u0\/u3\/_0077_ ), .X(\u0\/u3\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1047_ ( .A(\u0\/u3\/_0070_ ), .B(\u0\/u3\/_0035_ ), .X(\u0\/u3\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u3/_1048_ ( .A1(\u0\/u3\/_0047_ ), .A2(\u0\/u3\/_0736_ ), .B1(\u0\/u3\/_0022_ ), .B2(\u0\/u3\/_0364_ ), .X(\u0\/u3\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u3/_1049_ ( .A(\u0\/u3\/_0239_ ), .B(\u0\/u3\/_0240_ ), .C(\u0\/u3\/_0241_ ), .Y(\u0\/u3\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1050_ ( .A(\u0\/u3\/_0554_ ), .B(\u0\/u3\/_0072_ ), .X(\u0\/u3\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u3/_1051_ ( .A1(\u0\/u3\/_0142_ ), .A2(\u0\/u3\/_0137_ ), .B1(\u0\/u3\/_0159_ ), .B2(\u0\/u3\/_0082_ ), .X(\u0\/u3\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1052_ ( .A1(\u0\/u3\/_0608_ ), .A2(\u0\/u3\/_0072_ ), .B1(\u0\/u3\/_0243_ ), .C1(\u0\/u3\/_0244_ ), .Y(\u0\/u3\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1053_ ( .A(\u0\/u3\/_0234_ ), .B(\u0\/u3\/_0237_ ), .C(\u0\/u3\/_0242_ ), .D(\u0\/u3\/_0245_ ), .X(\u0\/u3\/_0246_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u3/_1055_ ( .A1(\u0\/u3\/_0554_ ), .A2(\u0\/u3\/_0586_ ), .B1(\u0\/u3\/_0029_ ), .X(\u0\/u3\/_0248_ ) );
sky130_fd_sc_hd__and2_1 \u0/u3/_1056_ ( .A(\u0\/u3\/_0082_ ), .B(\u0\/u3\/_0478_ ), .X(\u0\/u3\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_1057_ ( .A(\u0\/u3\/_0079_ ), .X(\u0\/u3\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1058_ ( .A(\u0\/u3\/_0251_ ), .B(\u0\/u3\/_0478_ ), .X(\u0\/u3\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_1059_ ( .A(\u0\/u3\/_0250_ ), .B(\u0\/u3\/_0252_ ), .Y(\u0\/u3\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1060_ ( .A(\u0\/u3\/_0016_ ), .B(\u0\/u3\/_0064_ ), .Y(\u0\/u3\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_1061_ ( .A(\u0\/u3\/_0304_ ), .X(\u0\/u3\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1062_ ( .A(\u0\/u3\/_0255_ ), .B(\u0\/u3\/_0640_ ), .Y(\u0\/u3\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u3/_1063_ ( .A_N(\u0\/u3\/_0248_ ), .B(\u0\/u3\/_0253_ ), .C(\u0\/u3\/_0254_ ), .D(\u0\/u3\/_0256_ ), .X(\u0\/u3\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1064_ ( .A(\u0\/u3\/_0364_ ), .B(\u0\/u3\/_0110_ ), .X(\u0\/u3\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \u0/u3/_1065_ ( .A1(\u0\/u3\/_0161_ ), .A2(\u0\/u3\/_0130_ ), .B1(\u0\/u3\/_0258_ ), .Y(\u0\/u3\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1066_ ( .A(\u0\/u3\/_0194_ ), .B(\w3\[25\] ), .X(\u0\/u3\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1068_ ( .A(\u0\/u3\/_0261_ ), .B(\u0\/u3\/_0153_ ), .Y(\u0\/u3\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u3/_1069_ ( .A_N(\u0\/u3\/_0154_ ), .B(\u0\/u3\/_0259_ ), .C(\u0\/u3\/_0263_ ), .X(\u0\/u3\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1070_ ( .A(\u0\/u3\/_0246_ ), .B(\u0\/u3\/_0174_ ), .C(\u0\/u3\/_0257_ ), .D(\u0\/u3\/_0264_ ), .X(\u0\/u3\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u3/_1071_ ( .A1(\u0\/u3\/_0261_ ), .A2(\u0\/u3\/_0554_ ), .B1(\u0\/u3\/_0159_ ), .X(\u0\/u3\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1072_ ( .A(\u0\/u3\/_0746_ ), .B(\u0\/u3\/_0150_ ), .Y(\u0\/u3\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1073_ ( .A(\u0\/u3\/_0175_ ), .Y(\u0\/u3\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \u0/u3/_1074_ ( .A(\u0\/u3\/_0412_ ), .B(\u0\/u3\/_0123_ ), .C(\u0\/u3\/_0151_ ), .X(\u0\/u3\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1075_ ( .A(\u0\/u3\/_0268_ ), .B(\u0\/u3\/_0269_ ), .Y(\u0\/u3\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u3/_1076_ ( .A_N(\u0\/u3\/_0266_ ), .B(\u0\/u3\/_0267_ ), .C(\u0\/u3\/_0270_ ), .X(\u0\/u3\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1077_ ( .A(\u0\/u3\/_0554_ ), .B(\u0\/u3\/_0150_ ), .X(\u0\/u3\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1078_ ( .A(\u0\/u3\/_0273_ ), .Y(\u0\/u3\/_0274_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u3/_1079_ ( .A1(\u0\/u3\/_0734_ ), .A2(\u0\/u3\/_0325_ ), .B1(\u0\/u3\/_0380_ ), .Y(\u0\/u3\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1080_ ( .A(\u0\/u3\/_0275_ ), .Y(\u0\/u3\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1081_ ( .A(\u0\/u3\/_0276_ ), .B(\u0\/u3\/_0153_ ), .Y(\u0\/u3\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \u0/u3/_1082_ ( .A(\u0\/u3\/_0272_ ), .B(\u0\/u3\/_0274_ ), .C(\u0\/u3\/_0277_ ), .X(\u0\/u3\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_1083_ ( .A(\u0\/u3\/_0035_ ), .X(\u0\/u3\/_0279_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1085_ ( .A1(\u0\/u3\/_0218_ ), .A2(\u0\/u3\/_0279_ ), .B1(\u0\/u3\/_0084_ ), .B2(\u0\/u3\/_0060_ ), .Y(\u0\/u3\/_0281_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1086_ ( .A1(\u0\/u3\/_0251_ ), .A2(\u0\/u3\/_0434_ ), .B1(\u0\/u3\/_0304_ ), .Y(\u0\/u3\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1087_ ( .A(\u0\/u3\/_0091_ ), .B(\u0\/u3\/_0292_ ), .Y(\u0\/u3\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1088_ ( .A1(\u0\/u3\/_0118_ ), .A2(\u0\/u3\/_0050_ ), .B1(\u0\/u3\/_0038_ ), .C1(\u0\/u3\/_0255_ ), .Y(\u0\/u3\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1089_ ( .A(\u0\/u3\/_0281_ ), .B(\u0\/u3\/_0283_ ), .C(\u0\/u3\/_0284_ ), .D(\u0\/u3\/_0285_ ), .X(\u0\/u3\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1090_ ( .A(\u0\/u3\/_0082_ ), .B(\u0\/u3\/_0027_ ), .X(\u0\/u3\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1091_ ( .A(\u0\/u3\/_0129_ ), .B(\u0\/u3\/_0027_ ), .X(\u0\/u3\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_1092_ ( .A(\u0\/u3\/_0287_ ), .B(\u0\/u3\/_0288_ ), .Y(\u0\/u3\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1093_ ( .A1(\u0\/u3\/_0752_ ), .A2(\u0\/u3\/_0683_ ), .B1(\u0\/u3\/_0093_ ), .B2(\u0\/u3\/_0029_ ), .Y(\u0\/u3\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1094_ ( .A1(\u0\/u3\/_0092_ ), .A2(\u0\/u3\/_0575_ ), .B1(\u0\/u3\/_0292_ ), .Y(\u0\/u3\/_0291_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_1095_ ( .A(\u0\/u3\/_0054_ ), .X(\u0\/u3\/_0292_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1096_ ( .A1(\u0\/u3\/_0218_ ), .A2(\u0\/u3\/_0662_ ), .B1(\u0\/u3\/_0084_ ), .B2(\u0\/u3\/_0292_ ), .Y(\u0\/u3\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1097_ ( .A(\u0\/u3\/_0289_ ), .B(\u0\/u3\/_0290_ ), .C(\u0\/u3\/_0291_ ), .D(\u0\/u3\/_0294_ ), .X(\u0\/u3\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1098_ ( .A(\u0\/u3\/_0750_ ), .B(\u0\/u3\/_0193_ ), .X(\u0\/u3\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1099_ ( .A(\u0\/u3\/_0705_ ), .B(\u0\/u3\/_0380_ ), .X(\u0\/u3\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1100_ ( .A(\u0\/u3\/_0752_ ), .B(\u0\/u3\/_0129_ ), .Y(\u0\/u3\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u3/_1101_ ( .A(\u0\/u3\/_0296_ ), .B(\u0\/u3\/_0297_ ), .C_N(\u0\/u3\/_0298_ ), .Y(\u0\/u3\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1102_ ( .A(\u0\/u3\/_0089_ ), .B(\u0\/u3\/_0532_ ), .Y(\u0\/u3\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1103_ ( .A(\w3\[26\] ), .Y(\u0\/u3\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u3/_1104_ ( .A(\u0\/u3\/_0301_ ), .B(\w3\[27\] ), .C(\u0\/u3\/_0118_ ), .Y(\u0\/u3\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1105_ ( .A(\u0\/u3\/_0072_ ), .B(\u0\/u3\/_0302_ ), .X(\u0\/u3\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1106_ ( .A(\u0\/u3\/_0303_ ), .Y(\u0\/u3\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1107_ ( .A(\u0\/u3\/_0147_ ), .B(\u0\/u3\/_0302_ ), .Y(\u0\/u3\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1108_ ( .A(\u0\/u3\/_0299_ ), .B(\u0\/u3\/_0300_ ), .C(\u0\/u3\/_0305_ ), .D(\u0\/u3\/_0306_ ), .X(\u0\/u3\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1109_ ( .A(\u0\/u3\/_0278_ ), .B(\u0\/u3\/_0286_ ), .C(\u0\/u3\/_0295_ ), .D(\u0\/u3\/_0307_ ), .X(\u0\/u3\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u3/_1110_ ( .A(\u0\/u3\/_0228_ ), .B(\u0\/u3\/_0265_ ), .C(\u0\/u3\/_0308_ ), .Y(\u0\/u3\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1111_ ( .A(\u0\/u3\/_0235_ ), .Y(\u0\/u3\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1112_ ( .A(\u0\/u3\/_0478_ ), .B(\u0\/u3\/_0640_ ), .X(\u0\/u3\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1113_ ( .A(\u0\/u3\/_0310_ ), .Y(\u0\/u3\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1114_ ( .A(\u0\/u3\/_0022_ ), .B(\u0\/u3\/_0218_ ), .Y(\u0\/u3\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1115_ ( .A(\u0\/u3\/_0218_ ), .B(\u0\/u3\/_0032_ ), .Y(\u0\/u3\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1116_ ( .A(\u0\/u3\/_0309_ ), .B(\u0\/u3\/_0311_ ), .C(\u0\/u3\/_0312_ ), .D(\u0\/u3\/_0313_ ), .X(\u0\/u3\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1117_ ( .A(\u0\/u3\/_0218_ ), .B(\u0\/u3\/_0064_ ), .Y(\u0\/u3\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1118_ ( .A(\u0\/u3\/_0218_ ), .B(\u0\/u3\/_0683_ ), .Y(\u0\/u3\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1119_ ( .A(\u0\/u3\/_0315_ ), .B(\u0\/u3\/_0316_ ), .C(\u0\/u3\/_0317_ ), .D(\u0\/u3\/_0253_ ), .X(\u0\/u3\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1120_ ( .A(\u0\/u3\/_0047_ ), .B(\u0\/u3\/_0304_ ), .Y(\u0\/u3\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1121_ ( .A(\u0\/u3\/_0586_ ), .B(\u0\/u3\/_0162_ ), .Y(\u0\/u3\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1122_ ( .A(\u0\/u3\/_0319_ ), .B(\u0\/u3\/_0320_ ), .Y(\u0\/u3\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_1123_ ( .A(\u0\/u3\/_0321_ ), .B(\u0\/u3\/_0238_ ), .Y(\u0\/u3\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1124_ ( .A(\u0\/u3\/_0304_ ), .B(\u0\/u3\/_0062_ ), .Y(\u0\/u3\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_1125_ ( .A(\u0\/u3\/_0251_ ), .X(\u0\/u3\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1126_ ( .A1(\u0\/u3\/_0324_ ), .A2(\u0\/u3\/_0084_ ), .B1(\u0\/u3\/_0255_ ), .Y(\u0\/u3\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1127_ ( .A1(\u0\/u3\/_0050_ ), .A2(\u0\/u3\/_0216_ ), .B1(\u0\/u3\/_0109_ ), .C1(\u0\/u3\/_0255_ ), .Y(\u0\/u3\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1128_ ( .A(\u0\/u3\/_0322_ ), .B(\u0\/u3\/_0323_ ), .C(\u0\/u3\/_0326_ ), .D(\u0\/u3\/_0327_ ), .X(\u0\/u3\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1129_ ( .A1(\u0\/u3\/_0733_ ), .A2(\u0\/u3\/_0279_ ), .A3(\u0\/u3\/_0058_ ), .B1(\u0\/u3\/_0292_ ), .Y(\u0\/u3\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_1130_ ( .A(\u0\/u3\/_0047_ ), .X(\u0\/u3\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1131_ ( .A(\u0\/u3\/_0330_ ), .B(\u0\/u3\/_0292_ ), .Y(\u0\/u3\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1132_ ( .A(\u0\/u3\/_0054_ ), .B(\u0\/u3\/_0045_ ), .Y(\u0\/u3\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1133_ ( .A(\u0\/u3\/_0329_ ), .B(\u0\/u3\/_0331_ ), .C(\u0\/u3\/_0284_ ), .D(\u0\/u3\/_0332_ ), .X(\u0\/u3\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u3/_1134_ ( .A1(\u0\/u3\/_0249_ ), .A2(\u0\/u3\/_0216_ ), .B1(\u0\/u3\/_0532_ ), .C1(\u0\/u3\/_0060_ ), .X(\u0\/u3\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1135_ ( .A(\u0\/u3\/_0084_ ), .B(\u0\/u3\/_0060_ ), .Y(\u0\/u3\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1136_ ( .A(\u0\/u3\/_0324_ ), .B(\u0\/u3\/_0060_ ), .Y(\u0\/u3\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1137_ ( .A(\u0\/u3\/_0335_ ), .B(\u0\/u3\/_0337_ ), .Y(\u0\/u3\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1138_ ( .A1(\u0\/u3\/_0276_ ), .A2(\u0\/u3\/_0060_ ), .B1(\u0\/u3\/_0334_ ), .C1(\u0\/u3\/_0338_ ), .Y(\u0\/u3\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1139_ ( .A(\u0\/u3\/_0318_ ), .B(\u0\/u3\/_0328_ ), .C(\u0\/u3\/_0333_ ), .D(\u0\/u3\/_0339_ ), .X(\u0\/u3\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u3/_1140_ ( .A1(\u0\/u3\/_0746_ ), .A2(\u0\/u3\/_0134_ ), .B1(\u0\/u3\/_0128_ ), .X(\u0\/u3\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u3/_1141_ ( .A_N(\u0\/u3\/_0086_ ), .B(\u0\/u3\/_0128_ ), .X(\u0\/u3\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1142_ ( .A(\u0\/u3\/_0079_ ), .B(\u0\/u3\/_0124_ ), .X(\u0\/u3\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_1143_ ( .A(\u0\/u3\/_0126_ ), .B(\u0\/u3\/_0343_ ), .Y(\u0\/u3\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u3/_1144_ ( .A(\u0\/u3\/_0341_ ), .B(\u0\/u3\/_0342_ ), .C_N(\u0\/u3\/_0344_ ), .Y(\u0\/u3\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1146_ ( .A1(\u0\/u3\/_0193_ ), .A2(\u0\/u3\/_0092_ ), .A3(\u0\/u3\/_0330_ ), .B1(\u0\/u3\/_0147_ ), .Y(\u0\/u3\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1147_ ( .A1(\u0\/u3\/_0130_ ), .A2(\u0\/u3\/_0084_ ), .A3(\u0\/u3\/_0134_ ), .B1(\u0\/u3\/_0139_ ), .Y(\u0\/u3\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1148_ ( .A1(\u0\/u3\/_0144_ ), .A2(\u0\/u3\/_0608_ ), .A3(\u0\/u3\/_0092_ ), .B1(\u0\/u3\/_0139_ ), .Y(\u0\/u3\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1149_ ( .A(\u0\/u3\/_0345_ ), .B(\u0\/u3\/_0348_ ), .C(\u0\/u3\/_0349_ ), .D(\u0\/u3\/_0350_ ), .X(\u0\/u3\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \u0/u3/_1150_ ( .A(\u0\/u3\/_0150_ ), .B(\u0\/u3\/_0194_ ), .C(\u0\/u3\/_0249_ ), .X(\u0\/u3\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u3/_1151_ ( .A(\u0\/u3\/_0277_ ), .SLEEP(\u0\/u3\/_0352_ ), .X(\u0\/u3\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \u0/u3/_1152_ ( .A1(\u0\/u3\/_0268_ ), .A2(\u0\/u3\/_0171_ ), .B1(\u0\/u3\/_0157_ ), .Y(\u0\/u3\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_1153_ ( .A(\u0\/u3\/_0161_ ), .X(\u0\/u3\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1154_ ( .A1(\u0\/u3\/_0279_ ), .A2(\u0\/u3\/_0084_ ), .B1(\u0\/u3\/_0355_ ), .Y(\u0\/u3\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1155_ ( .A1(\u0\/u3\/_0020_ ), .A2(\u0\/u3\/_0193_ ), .A3(\u0\/u3\/_0091_ ), .B1(\u0\/u3\/_0355_ ), .Y(\u0\/u3\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1156_ ( .A(\u0\/u3\/_0353_ ), .B(\u0\/u3\/_0354_ ), .C(\u0\/u3\/_0356_ ), .D(\u0\/u3\/_0357_ ), .X(\u0\/u3\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1157_ ( .A(\u0\/u3\/_0111_ ), .B(\u0\/u3\/_0586_ ), .X(\u0\/u3\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1158_ ( .A(\u0\/u3\/_0360_ ), .Y(\u0\/u3\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u3/_1159_ ( .A1(\u0\/u3\/_0119_ ), .A2(\u0\/u3\/_0120_ ), .B1(\u0\/u3\/_0230_ ), .C1(\u0\/u3\/_0361_ ), .X(\u0\/u3\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1160_ ( .A1(\u0\/u3\/_0662_ ), .A2(\u0\/u3\/_0251_ ), .A3(\u0\/u3\/_0134_ ), .B1(\u0\/u3\/_0114_ ), .Y(\u0\/u3\/_0363_ ) );
sky130_fd_sc_hd__buf_2 \u0/u3/_1161_ ( .A(\u0\/u3\/_0098_ ), .X(\u0\/u3\/_0364_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1162_ ( .A1(\u0\/u3\/_0035_ ), .A2(\u0\/u3\/_0251_ ), .A3(\u0\/u3\/_0134_ ), .B1(\u0\/u3\/_0364_ ), .Y(\u0\/u3\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1163_ ( .A1(\u0\/u3\/_0193_ ), .A2(\u0\/u3\/_0608_ ), .B1(\u0\/u3\/_0364_ ), .Y(\u0\/u3\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1164_ ( .A(\u0\/u3\/_0362_ ), .B(\u0\/u3\/_0363_ ), .C(\u0\/u3\/_0365_ ), .D(\u0\/u3\/_0366_ ), .X(\u0\/u3\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1165_ ( .A1(\u0\/u3\/_0575_ ), .A2(\u0\/u3\/_0092_ ), .A3(\u0\/u3\/_0330_ ), .B1(\u0\/u3\/_0089_ ), .Y(\u0\/u3\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1166_ ( .A1(\u0\/u3\/_0586_ ), .A2(\u0\/u3\/_0017_ ), .A3(\u0\/u3\/_0330_ ), .B1(\u0\/u3\/_0094_ ), .Y(\u0\/u3\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u3/_1167_ ( .A1(\u0\/u3\/_0293_ ), .A2(\u0\/u3\/_0134_ ), .B1(\u0\/u3\/_0089_ ), .Y(\u0\/u3\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1168_ ( .A1(\u0\/u3\/_0279_ ), .A2(\u0\/u3\/_0134_ ), .B1(\u0\/u3\/_0094_ ), .Y(\u0\/u3\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1169_ ( .A(\u0\/u3\/_0368_ ), .B(\u0\/u3\/_0370_ ), .C(\u0\/u3\/_0371_ ), .D(\u0\/u3\/_0372_ ), .X(\u0\/u3\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1170_ ( .A(\u0\/u3\/_0351_ ), .B(\u0\/u3\/_0359_ ), .C(\u0\/u3\/_0367_ ), .D(\u0\/u3\/_0373_ ), .X(\u0\/u3\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1171_ ( .A1(\u0\/u3\/_0102_ ), .A2(\u0\/u3\/_0347_ ), .B1(\u0\/u3\/_0109_ ), .C1(\u0\/u3\/_0029_ ), .Y(\u0\/u3\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1172_ ( .A1(\u0\/u3\/_0102_ ), .A2(\u0\/u3\/_0347_ ), .B1(\u0\/u3\/_0532_ ), .C1(\u0\/u3\/_0029_ ), .Y(\u0\/u3\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1173_ ( .A1(\u0\/u3\/_0050_ ), .A2(\u0\/u3\/_0249_ ), .B1(\u0\/u3\/_0380_ ), .C1(\u0\/u3\/_0029_ ), .Y(\u0\/u3\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1174_ ( .A(\u0\/u3\/_0041_ ), .B(\u0\/u3\/_0375_ ), .C(\u0\/u3\/_0376_ ), .D(\u0\/u3\/_0377_ ), .X(\u0\/u3\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1175_ ( .A(\u0\/u3\/_0047_ ), .B(\u0\/u3\/_0750_ ), .X(\u0\/u3\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1176_ ( .A(\u0\/u3\/_0379_ ), .Y(\u0\/u3\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1177_ ( .A(\u0\/u3\/_0016_ ), .B(\u0\/u3\/_0608_ ), .Y(\u0\/u3\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1178_ ( .A(\u0\/u3\/_0752_ ), .B(\u0\/u3\/_0554_ ), .Y(\u0\/u3\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1179_ ( .A1(\w3\[25\] ), .A2(\u0\/u3\/_0734_ ), .B1(\u0\/u3\/_0109_ ), .C1(\u0\/u3\/_0016_ ), .Y(\u0\/u3\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1180_ ( .A(\u0\/u3\/_0381_ ), .B(\u0\/u3\/_0382_ ), .C(\u0\/u3\/_0383_ ), .D(\u0\/u3\/_0384_ ), .X(\u0\/u3\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \u0/u3/_1181_ ( .A(\u0\/u3\/_0086_ ), .B_N(\u0\/u3\/_0736_ ), .X(\u0\/u3\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1182_ ( .A1(\u0\/u3\/_0748_ ), .A2(\u0\/u3\/_0134_ ), .B1(\u0\/u3\/_0739_ ), .Y(\u0\/u3\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1183_ ( .A1(\u0\/u3\/_0118_ ), .A2(\u0\/u3\/_0249_ ), .B1(\u0\/u3\/_0109_ ), .C1(\u0\/u3\/_0739_ ), .Y(\u0\/u3\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1184_ ( .A1(\u0\/u3\/_0102_ ), .A2(\u0\/u3\/_0301_ ), .B1(\w3\[27\] ), .C1(\u0\/u3\/_0739_ ), .Y(\u0\/u3\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1185_ ( .A(\u0\/u3\/_0386_ ), .B(\u0\/u3\/_0387_ ), .C(\u0\/u3\/_0388_ ), .D(\u0\/u3\/_0389_ ), .X(\u0\/u3\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1186_ ( .A(\u0\/u3\/_0020_ ), .Y(\u0\/u3\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1187_ ( .A(\u0\/u3\/_0727_ ), .Y(\u0\/u3\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1188_ ( .A(\u0\/u3\/_0727_ ), .B(\u0\/u3\/_0064_ ), .Y(\u0\/u3\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1189_ ( .A1(\u0\/u3\/_0102_ ), .A2(\u0\/u3\/_0734_ ), .B1(\u0\/u3\/_0532_ ), .C1(\u0\/u3\/_0727_ ), .Y(\u0\/u3\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u3/_1190_ ( .A1(\u0\/u3\/_0392_ ), .A2(\u0\/u3\/_0393_ ), .B1(\u0\/u3\/_0394_ ), .C1(\u0\/u3\/_0395_ ), .X(\u0\/u3\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1191_ ( .A(\u0\/u3\/_0378_ ), .B(\u0\/u3\/_0385_ ), .C(\u0\/u3\/_0390_ ), .D(\u0\/u3\/_0396_ ), .X(\u0\/u3\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u3/_1192_ ( .A(\u0\/u3\/_0340_ ), .B(\u0\/u3\/_0374_ ), .C(\u0\/u3\/_0397_ ), .Y(\u0\/u3\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1193_ ( .A(\u0\/u3\/_0077_ ), .B(\u0\/u3\/_0129_ ), .X(\u0\/u3\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_1194_ ( .A(\u0\/u3\/_0398_ ), .B(\u0\/u3\/_0239_ ), .Y(\u0\/u3\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1195_ ( .A(\u0\/u3\/_0022_ ), .B(\u0\/u3\/_0111_ ), .X(\u0\/u3\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u3/_1196_ ( .A_N(\u0\/u3\/_0400_ ), .B(\u0\/u3\/_0231_ ), .Y(\u0\/u3\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u3/_1197_ ( .A(\u0\/u3\/_0399_ ), .SLEEP(\u0\/u3\/_0402_ ), .X(\u0\/u3\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_1198_ ( .A(\u0\/u3\/_0746_ ), .B(\u0\/u3\/_0251_ ), .Y(\u0\/u3\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u3/_1199_ ( .A_N(\u0\/u3\/_0404_ ), .B(\u0\/u3\/_0752_ ), .Y(\u0\/u3\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \u0/u3/_1200_ ( .A(\u0\/u3\/_0467_ ), .B(\u0\/u3\/_0194_ ), .C(\u0\/u3\/_0694_ ), .X(\u0\/u3\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u3/_1201_ ( .A_N(\u0\/u3\/_0175_ ), .B(\u0\/u3\/_0406_ ), .X(\u0\/u3\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1202_ ( .A(\u0\/u3\/_0407_ ), .Y(\u0\/u3\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1203_ ( .A1(\u0\/u3\/_0094_ ), .A2(\u0\/u3\/_0197_ ), .B1(\u0\/u3\/_0114_ ), .B2(\u0\/u3\/_0640_ ), .Y(\u0\/u3\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1204_ ( .A(\u0\/u3\/_0403_ ), .B(\u0\/u3\/_0405_ ), .C(\u0\/u3\/_0408_ ), .D(\u0\/u3\/_0409_ ), .X(\u0\/u3\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1205_ ( .A(\u0\/u3\/_0030_ ), .B(\u0\/u3\/_0150_ ), .Y(\u0\/u3\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u3/_1206_ ( .A_N(\u0\/u3\/_0169_ ), .B(\u0\/u3\/_0289_ ), .C(\u0\/u3\/_0411_ ), .X(\u0\/u3\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u3/_1207_ ( .A1(\u0\/u3\/_0467_ ), .A2(\u0\/u3\/_0151_ ), .B1(\u0\/u3\/_0140_ ), .C1(\u0\/u3\/_0129_ ), .X(\u0\/u3\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1208_ ( .A1(\u0\/u3\/_0608_ ), .A2(\u0\/u3\/_0364_ ), .B1(\u0\/u3\/_0037_ ), .C1(\u0\/u3\/_0414_ ), .Y(\u0\/u3\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1209_ ( .A(\u0\/u3\/_0738_ ), .Y(\u0\/u3\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1210_ ( .A(\u0\/u3\/_0586_ ), .B(\u0\/u3\/_0736_ ), .Y(\u0\/u3\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1211_ ( .A1(\u0\/u3\/_0194_ ), .A2(\u0\/u3\/_0038_ ), .B1(\u0\/u3\/_0118_ ), .C1(\u0\/u3\/_0153_ ), .Y(\u0\/u3\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u3/_1212_ ( .A1(\u0\/u3\/_0416_ ), .A2(\u0\/u3\/_0117_ ), .B1(\u0\/u3\/_0417_ ), .C1(\u0\/u3\/_0418_ ), .X(\u0\/u3\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1213_ ( .A(\u0\/u3\/_0077_ ), .B(\u0\/u3\/_0035_ ), .X(\u0\/u3\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1214_ ( .A(\u0\/u3\/_0662_ ), .B(\u0\/u3\/_0124_ ), .Y(\u0\/u3\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1215_ ( .A(\u0\/u3\/_0030_ ), .B(\u0\/u3\/_0137_ ), .Y(\u0\/u3\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1216_ ( .A(\u0\/u3\/_0072_ ), .B(\u0\/u3\/_0731_ ), .Y(\u0\/u3\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u3/_1217_ ( .A_N(\u0\/u3\/_0420_ ), .B(\u0\/u3\/_0421_ ), .C(\u0\/u3\/_0422_ ), .D(\u0\/u3\/_0424_ ), .X(\u0\/u3\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1218_ ( .A(\u0\/u3\/_0413_ ), .B(\u0\/u3\/_0415_ ), .C(\u0\/u3\/_0419_ ), .D(\u0\/u3\/_0425_ ), .X(\u0\/u3\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u3/_1219_ ( .A(\u0\/u3\/_0355_ ), .B(\u0\/u3\/_0102_ ), .C(\u0\/u3\/_0109_ ), .Y(\u0\/u3\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1220_ ( .A(\u0\/u3\/_0077_ ), .B(\u0\/u3\/_0017_ ), .X(\u0\/u3\/_0428_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1221_ ( .A(\u0\/u3\/_0077_ ), .B(\u0\/u3\/_0554_ ), .X(\u0\/u3\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u3/_1222_ ( .A1(\u0\/u3\/_0050_ ), .A2(\u0\/u3\/_0216_ ), .B1(\u0\/u3\/_0380_ ), .C1(\u0\/u3\/_0078_ ), .X(\u0\/u3\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u3/_1223_ ( .A(\u0\/u3\/_0428_ ), .B(\u0\/u3\/_0429_ ), .C(\u0\/u3\/_0430_ ), .Y(\u0\/u3\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u3/_1224_ ( .A_N(\u0\/u3\/_0209_ ), .B(\u0\/u3\/_0431_ ), .X(\u0\/u3\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u3/_1225_ ( .A1(\u0\/u3\/_0215_ ), .A2(\u0\/u3\/_0404_ ), .B1(\u0\/u3\/_0427_ ), .C1(\u0\/u3\/_0432_ ), .X(\u0\/u3\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1226_ ( .A(\u0\/u3\/_0043_ ), .B(\u0\/u3\/_0058_ ), .Y(\u0\/u3\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1227_ ( .A(\u0\/u3\/_0195_ ), .B(\u0\/u3\/_0233_ ), .C(\u0\/u3\/_0320_ ), .D(\u0\/u3\/_0435_ ), .X(\u0\/u3\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1228_ ( .A(\u0\/u3\/_0261_ ), .B(\u0\/u3\/_0738_ ), .Y(\u0\/u3\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1229_ ( .A1(\u0\/u3\/_0218_ ), .A2(\u0\/u3\/_0640_ ), .B1(\u0\/u3\/_0261_ ), .B2(\u0\/u3\/_0292_ ), .Y(\u0\/u3\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1230_ ( .A(\u0\/u3\/_0436_ ), .B(\u0\/u3\/_0394_ ), .C(\u0\/u3\/_0437_ ), .D(\u0\/u3\/_0438_ ), .X(\u0\/u3\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1231_ ( .A(\u0\/u3\/_0410_ ), .B(\u0\/u3\/_0426_ ), .C(\u0\/u3\/_0433_ ), .D(\u0\/u3\/_0439_ ), .X(\u0\/u3\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \u0/u3/_1232_ ( .A(\u0\/u3\/_0135_ ), .SLEEP(\u0\/u3\/_0273_ ), .X(\u0\/u3\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1233_ ( .A1(\u0\/u3\/_0279_ ), .A2(\u0\/u3\/_0134_ ), .B1(\u0\/u3\/_0364_ ), .Y(\u0\/u3\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1234_ ( .A(\u0\/u3\/_0441_ ), .B(\u0\/u3\/_0164_ ), .C(\u0\/u3\/_0270_ ), .D(\u0\/u3\/_0442_ ), .X(\u0\/u3\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1235_ ( .A(\u0\/u3\/_0051_ ), .B(\u0\/u3\/_0662_ ), .Y(\u0\/u3\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1236_ ( .A(\u0\/u3\/_0051_ ), .B(\u0\/u3\/_0271_ ), .Y(\u0\/u3\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1237_ ( .A(\u0\/u3\/_0444_ ), .B(\u0\/u3\/_0446_ ), .X(\u0\/u3\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1238_ ( .A(\u0\/u3\/_0193_ ), .B(\u0\/u3\/_0304_ ), .X(\u0\/u3\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1239_ ( .A(\u0\/u3\/_0448_ ), .Y(\u0\/u3\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1240_ ( .A(\u0\/u3\/_0162_ ), .B(\u0\/u3\/_0130_ ), .X(\u0\/u3\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1241_ ( .A(\u0\/u3\/_0450_ ), .Y(\u0\/u3\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1242_ ( .A1(\u0\/u3\/_0129_ ), .A2(\u0\/u3\/_0554_ ), .B1(\u0\/u3\/_0043_ ), .Y(\u0\/u3\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1243_ ( .A(\u0\/u3\/_0447_ ), .B(\u0\/u3\/_0449_ ), .C(\u0\/u3\/_0451_ ), .D(\u0\/u3\/_0452_ ), .X(\u0\/u3\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1244_ ( .A(\u0\/u3\/_0292_ ), .B(\u0\/u3\/_0064_ ), .Y(\u0\/u3\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u3/_1245_ ( .A_N(\u0\/u3\/_0248_ ), .B(\u0\/u3\/_0454_ ), .C(\u0\/u3\/_0254_ ), .D(\u0\/u3\/_0256_ ), .X(\u0\/u3\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1246_ ( .A1(\u0\/u3\/_0330_ ), .A2(\u0\/u3\/_0364_ ), .B1(\u0\/u3\/_0134_ ), .B2(\u0\/u3\/_0705_ ), .Y(\u0\/u3\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1247_ ( .A1(\u0\/u3\/_0748_ ), .A2(\u0\/u3\/_0738_ ), .B1(\u0\/u3\/_0092_ ), .B2(\u0\/u3\/_0752_ ), .Y(\u0\/u3\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1248_ ( .A1(\u0\/u3\/_0072_ ), .A2(\u0\/u3\/_0035_ ), .B1(\u0\/u3\/_0748_ ), .B2(\u0\/u3\/_0292_ ), .Y(\u0\/u3\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1249_ ( .A1(\u0\/u3\/_0748_ ), .A2(\u0\/u3\/_0251_ ), .B1(\u0\/u3\/_0029_ ), .Y(\u0\/u3\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1250_ ( .A(\u0\/u3\/_0457_ ), .B(\u0\/u3\/_0458_ ), .C(\u0\/u3\/_0459_ ), .D(\u0\/u3\/_0460_ ), .X(\u0\/u3\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1251_ ( .A(\u0\/u3\/_0443_ ), .B(\u0\/u3\/_0453_ ), .C(\u0\/u3\/_0455_ ), .D(\u0\/u3\/_0461_ ), .X(\u0\/u3\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1252_ ( .A(\u0\/u3\/_0705_ ), .B(\u0\/u3\/_0079_ ), .X(\u0\/u3\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1253_ ( .A(\u0\/u3\/_0586_ ), .B(\u0\/u3\/_0124_ ), .Y(\u0\/u3\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1254_ ( .A(\u0\/u3\/_0218_ ), .B(\u0\/u3\/_0746_ ), .Y(\u0\/u3\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u3/_1255_ ( .A_N(\u0\/u3\/_0463_ ), .B(\u0\/u3\/_0464_ ), .C(\u0\/u3\/_0465_ ), .X(\u0\/u3\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u3/_1256_ ( .A1(\u0\/u3\/_0271_ ), .A2(\u0\/u3\/_0072_ ), .B1(\u0\/u3\/_0142_ ), .B2(\u0\/u3\/_0027_ ), .X(\u0\/u3\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1257_ ( .A1(\u0\/u3\/_0144_ ), .A2(\u0\/u3\/_0364_ ), .B1(\u0\/u3\/_0360_ ), .C1(\u0\/u3\/_0468_ ), .Y(\u0\/u3\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u3/_1258_ ( .A1(\u0\/u3\/_0662_ ), .A2(\u0\/u3\/_0251_ ), .B1(\u0\/u3\/_0218_ ), .X(\u0\/u3\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1259_ ( .A1(\u0\/u3\/_0575_ ), .A2(\u0\/u3\/_0292_ ), .B1(\u0\/u3\/_0379_ ), .C1(\u0\/u3\/_0470_ ), .Y(\u0\/u3\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1260_ ( .A(\u0\/u3\/_0466_ ), .B(\u0\/u3\/_0469_ ), .C(\u0\/u3\/_0471_ ), .D(\u0\/u3\/_0305_ ), .X(\u0\/u3\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u3/_1261_ ( .A1(\u0\/u3\/_0029_ ), .A2(\u0\/u3\/_0683_ ), .B1(\u0\/u3\/_0324_ ), .B2(\u0\/u3\/_0292_ ), .X(\u0\/u3\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1262_ ( .A(\u0\/u3\/_0084_ ), .B(\u0\/u3\/_0364_ ), .X(\u0\/u3\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \u0/u3/_1263_ ( .A1(\u0\/u3\/_0092_ ), .A2(\u0\/u3\/_0029_ ), .B1(\u0\/u3\/_0474_ ), .X(\u0\/u3\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u3/_1264_ ( .A(\u0\/u3\/_0075_ ), .B(\u0\/u3\/_0473_ ), .C(\u0\/u3\/_0475_ ), .Y(\u0\/u3\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1265_ ( .A1(\u0\/u3\/_0279_ ), .A2(\u0\/u3\/_0255_ ), .B1(\u0\/u3\/_0084_ ), .B2(\u0\/u3\/_0060_ ), .Y(\u0\/u3\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1266_ ( .A1(\u0\/u3\/_0093_ ), .A2(\u0\/u3\/_0292_ ), .B1(\u0\/u3\/_0134_ ), .B2(\u0\/u3\/_0114_ ), .Y(\u0\/u3\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1267_ ( .A1(\u0\/u3\/_0161_ ), .A2(\u0\/u3\/_0032_ ), .B1(\u0\/u3\/_0324_ ), .B2(\u0\/u3\/_0147_ ), .Y(\u0\/u3\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1268_ ( .A1(\u0\/u3\/_0054_ ), .A2(\u0\/u3\/_0731_ ), .B1(\u0\/u3\/_0748_ ), .B2(\u0\/u3\/_0304_ ), .Y(\u0\/u3\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1269_ ( .A(\u0\/u3\/_0477_ ), .B(\u0\/u3\/_0479_ ), .C(\u0\/u3\/_0480_ ), .D(\u0\/u3\/_0481_ ), .X(\u0\/u3\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1270_ ( .A(\u0\/u3\/_0161_ ), .B(\u0\/u3\/_0064_ ), .Y(\u0\/u3\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u3/_1271_ ( .A(\u0\/u3\/_0731_ ), .B(\u0\/u3\/_0123_ ), .C(\u0\/u3\/_0467_ ), .Y(\u0\/u3\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1272_ ( .A(\u0\/u3\/_0483_ ), .B(\u0\/u3\/_0484_ ), .Y(\u0\/u3\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1273_ ( .A(\u0\/u3\/_0297_ ), .Y(\u0\/u3\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u3/_1274_ ( .A_N(\u0\/u3\/_0485_ ), .B(\u0\/u3\/_0181_ ), .C(\u0\/u3\/_0486_ ), .D(\u0\/u3\/_0386_ ), .X(\u0\/u3\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1275_ ( .A(\u0\/u3\/_0472_ ), .B(\u0\/u3\/_0476_ ), .C(\u0\/u3\/_0482_ ), .D(\u0\/u3\/_0487_ ), .X(\u0\/u3\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u3/_1276_ ( .A(\u0\/u3\/_0440_ ), .B(\u0\/u3\/_0462_ ), .C(\u0\/u3\/_0488_ ), .Y(\u0\/u3\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1277_ ( .A(\u0\/u3\/_0403_ ), .B(\u0\/u3\/_0230_ ), .C(\u0\/u3\/_0451_ ), .D(\u0\/u3\/_0361_ ), .X(\u0\/u3\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1278_ ( .A1(\u0\/u3\/_0118_ ), .A2(\u0\/u3\/_0050_ ), .B1(\u0\/u3\/_0109_ ), .C1(\u0\/u3\/_0139_ ), .Y(\u0\/u3\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1279_ ( .A(\u0\/u3\/_0447_ ), .B(\u0\/u3\/_0437_ ), .C(\u0\/u3\/_0491_ ), .D(\u0\/u3\/_0427_ ), .X(\u0\/u3\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1280_ ( .A1(\u0\/u3\/_0084_ ), .A2(\u0\/u3\/_0255_ ), .B1(\u0\/u3\/_0608_ ), .B2(\u0\/u3\/_0029_ ), .Y(\u0\/u3\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1281_ ( .A1(\u0\/u3\/_0144_ ), .A2(\u0\/u3\/_0147_ ), .B1(\u0\/u3\/_0355_ ), .B2(\u0\/u3\/_0093_ ), .Y(\u0\/u3\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1282_ ( .A1(\u0\/u3\/_0705_ ), .A2(\u0\/u3\/_0279_ ), .B1(\u0\/u3\/_0330_ ), .B2(\u0\/u3\/_0029_ ), .Y(\u0\/u3\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1283_ ( .A1(\u0\/u3\/_0279_ ), .A2(\u0\/u3\/_0084_ ), .B1(\u0\/u3\/_0114_ ), .Y(\u0\/u3\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1284_ ( .A(\u0\/u3\/_0493_ ), .B(\u0\/u3\/_0494_ ), .C(\u0\/u3\/_0495_ ), .D(\u0\/u3\/_0496_ ), .X(\u0\/u3\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1285_ ( .A1(\u0\/u3\/_0134_ ), .A2(\u0\/u3\/_0137_ ), .B1(\u0\/u3\/_0355_ ), .B2(\u0\/u3\/_0575_ ), .Y(\u0\/u3\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1286_ ( .A1(\u0\/u3\/_0364_ ), .A2(\u0\/u3\/_0733_ ), .B1(\u0\/u3\/_0093_ ), .B2(\u0\/u3\/_0218_ ), .Y(\u0\/u3\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1287_ ( .A(\u0\/u3\/_0147_ ), .B(\u0\/u3\/_0640_ ), .Y(\u0\/u3\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1288_ ( .A1(\u0\/u3\/_0153_ ), .A2(\u0\/u3\/_0292_ ), .B1(\u0\/u3\/_0748_ ), .Y(\u0\/u3\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1289_ ( .A(\u0\/u3\/_0498_ ), .B(\u0\/u3\/_0500_ ), .C(\u0\/u3\/_0501_ ), .D(\u0\/u3\/_0502_ ), .X(\u0\/u3\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1290_ ( .A(\u0\/u3\/_0490_ ), .B(\u0\/u3\/_0492_ ), .C(\u0\/u3\/_0497_ ), .D(\u0\/u3\/_0503_ ), .X(\u0\/u3\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u3/_1291_ ( .A_N(\u0\/u3\/_0275_ ), .B(\u0\/u3\/_0705_ ), .X(\u0\/u3\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1292_ ( .A(\u0\/u3\/_0505_ ), .Y(\u0\/u3\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1293_ ( .A(\u0\/u3\/_0380_ ), .B(\u0\/u3\/_0347_ ), .X(\u0\/u3\/_0507_ ) );
sky130_fd_sc_hd__o21ai_1 \u0/u3/_1294_ ( .A1(\u0\/u3\/_0507_ ), .A2(\u0\/u3\/_0093_ ), .B1(\u0\/u3\/_0292_ ), .Y(\u0\/u3\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1295_ ( .A(\u0\/u3\/_0322_ ), .B(\u0\/u3\/_0277_ ), .C(\u0\/u3\/_0506_ ), .D(\u0\/u3\/_0508_ ), .X(\u0\/u3\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1296_ ( .A(\u0\/u3\/_0084_ ), .B(\u0\/u3\/_0705_ ), .X(\u0\/u3\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1297_ ( .A1(\u0\/u3\/_0733_ ), .A2(\u0\/u3\/_0114_ ), .B1(\u0\/u3\/_0429_ ), .C1(\u0\/u3\/_0511_ ), .Y(\u0\/u3\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_1298_ ( .A(\u0\/u3\/_0019_ ), .B(\u0\/u3\/_0024_ ), .Y(\u0\/u3\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1299_ ( .A(\u0\/u3\/_0512_ ), .B(\u0\/u3\/_0513_ ), .C(\u0\/u3\/_0742_ ), .D(\u0\/u3\/_0306_ ), .X(\u0\/u3\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1300_ ( .A1(\u0\/u3\/_0532_ ), .A2(\u0\/u3\/_0089_ ), .B1(\u0\/u3\/_0154_ ), .C1(\u0\/u3\/_0169_ ), .Y(\u0\/u3\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u3/_1301_ ( .A1(\u0\/u3\/_0749_ ), .A2(\u0\/u3\/_0026_ ), .B1(\u0\/u3\/_0069_ ), .C1(\u0\/u3\/_0032_ ), .X(\u0\/u3\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u3/_1302_ ( .A1(\u0\/u3\/_0324_ ), .A2(\u0\/u3\/_0355_ ), .B1(\u0\/u3\/_0330_ ), .B2(\u0\/u3\/_0727_ ), .X(\u0\/u3\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u3/_1303_ ( .A(\u0\/u3\/_0133_ ), .B(\u0\/u3\/_0516_ ), .C(\u0\/u3\/_0517_ ), .Y(\u0\/u3\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1304_ ( .A(\u0\/u3\/_0509_ ), .B(\u0\/u3\/_0514_ ), .C(\u0\/u3\/_0515_ ), .D(\u0\/u3\/_0518_ ), .X(\u0\/u3\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1305_ ( .A(\u0\/u3\/_0746_ ), .B(\u0\/u3\/_0072_ ), .Y(\u0\/u3\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1306_ ( .A1(\u0\/u3\/_0082_ ), .A2(\u0\/u3\/_0070_ ), .B1(\u0\/u3\/_0043_ ), .B2(\u0\/u3\/_0193_ ), .Y(\u0\/u3\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1307_ ( .A(\u0\/u3\/_0311_ ), .B(\u0\/u3\/_0520_ ), .C(\u0\/u3\/_0332_ ), .D(\u0\/u3\/_0522_ ), .X(\u0\/u3\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1308_ ( .A(\u0\/u3\/_0129_ ), .B(\u0\/u3\/_0218_ ), .X(\u0\/u3\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_1309_ ( .A(\u0\/u3\/_0235_ ), .B(\u0\/u3\/_0524_ ), .Y(\u0\/u3\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \u0/u3/_1310_ ( .A(\u0\/u3\/_0081_ ), .B(\u0\/u3\/_0085_ ), .Y(\u0\/u3\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1311_ ( .A1(\u0\/u3\/_0051_ ), .A2(\u0\/u3\/_0045_ ), .B1(\u0\/u3\/_0130_ ), .B2(\u0\/u3\/_0094_ ), .Y(\u0\/u3\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1312_ ( .A(\u0\/u3\/_0523_ ), .B(\u0\/u3\/_0525_ ), .C(\u0\/u3\/_0526_ ), .D(\u0\/u3\/_0527_ ), .X(\u0\/u3\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u3/_1313_ ( .A_N(\u0\/u3\/_0250_ ), .B(\u0\/u3\/_0521_ ), .Y(\u0\/u3\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1314_ ( .A(\u0\/u3\/_0128_ ), .B(\u0\/u3\/_0020_ ), .X(\u0\/u3\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1315_ ( .A(\u0\/u3\/_0530_ ), .Y(\u0\/u3\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1316_ ( .A(\u0\/u3\/_0364_ ), .B(\u0\/u3\/_0058_ ), .X(\u0\/u3\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1317_ ( .A(\u0\/u3\/_0533_ ), .Y(\u0\/u3\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u3/_1318_ ( .A_N(\u0\/u3\/_0529_ ), .B(\u0\/u3\/_0531_ ), .C(\u0\/u3\/_0534_ ), .D(\u0\/u3\/_0192_ ), .X(\u0\/u3\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1319_ ( .A(\u0\/u3\/_0434_ ), .B(\u0\/u3\/_0078_ ), .X(\u0\/u3\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u3/_1320_ ( .A1(\u0\/u3\/_0750_ ), .A2(\u0\/u3\/_0079_ ), .B1(\u0\/u3\/_0129_ ), .B2(\u0\/u3\/_0705_ ), .X(\u0\/u3\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1321_ ( .A1(\u0\/u3\/_0161_ ), .A2(\u0\/u3\/_0032_ ), .B1(\u0\/u3\/_0536_ ), .C1(\u0\/u3\/_0537_ ), .Y(\u0\/u3\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u3/_1322_ ( .A1(\u0\/u3\/_0746_ ), .A2(\u0\/u3\/_0162_ ), .B1(\u0\/u3\/_0079_ ), .B2(\u0\/u3\/_0043_ ), .X(\u0\/u3\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1323_ ( .A1(\u0\/u3\/_0093_ ), .A2(\u0\/u3\/_0029_ ), .B1(\u0\/u3\/_0240_ ), .C1(\u0\/u3\/_0539_ ), .Y(\u0\/u3\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1324_ ( .A(\u0\/u3\/_0434_ ), .B(\u0\/u3\/_0043_ ), .X(\u0\/u3\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u3/_1325_ ( .A1(\u0\/u3\/_0142_ ), .A2(\u0\/u3\/_0150_ ), .B1(\u0\/u3\/_0022_ ), .B2(\u0\/u3\/_0137_ ), .X(\u0\/u3\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1326_ ( .A1(\u0\/u3\/_0279_ ), .A2(\u0\/u3\/_0051_ ), .B1(\u0\/u3\/_0541_ ), .C1(\u0\/u3\/_0542_ ), .Y(\u0\/u3\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1327_ ( .A(\u0\/u3\/_0159_ ), .B(\u0\/u3\/_0035_ ), .X(\u0\/u3\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u3/_1328_ ( .A1(\u0\/u3\/_0271_ ), .A2(\u0\/u3\/_0434_ ), .B1(\u0\/u3\/_0027_ ), .X(\u0\/u3\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1329_ ( .A1(\u0\/u3\/_0091_ ), .A2(\u0\/u3\/_0128_ ), .B1(\u0\/u3\/_0545_ ), .C1(\u0\/u3\/_0546_ ), .Y(\u0\/u3\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1330_ ( .A(\u0\/u3\/_0538_ ), .B(\u0\/u3\/_0540_ ), .C(\u0\/u3\/_0544_ ), .D(\u0\/u3\/_0547_ ), .X(\u0\/u3\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1331_ ( .A(\u0\/u3\/_0364_ ), .B(\u0\/u3\/_0193_ ), .X(\u0\/u3\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u3/_1332_ ( .A(\u0\/u3\/_0549_ ), .B(\u0\/u3\/_0186_ ), .C(\u0\/u3\/_0187_ ), .Y(\u0\/u3\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1333_ ( .A(\u0\/u3\/_0062_ ), .B(\u0\/u3\/_0347_ ), .C(\u0\/u3\/_0749_ ), .D(\u0\/u3\/_0694_ ), .X(\u0\/u3\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1334_ ( .A1(\u0\/u3\/_0130_ ), .A2(\u0\/u3\/_0218_ ), .B1(\u0\/u3\/_0551_ ), .C1(\u0\/u3\/_0101_ ), .Y(\u0\/u3\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1335_ ( .A(\u0\/u3\/_0139_ ), .B(\u0\/u3\/_0640_ ), .Y(\u0\/u3\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1336_ ( .A1(\u0\/u3\/_0752_ ), .A2(\u0\/u3\/_0662_ ), .B1(\u0\/u3\/_0084_ ), .B2(\u0\/u3\/_0364_ ), .Y(\u0\/u3\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1337_ ( .A(\u0\/u3\/_0550_ ), .B(\u0\/u3\/_0552_ ), .C(\u0\/u3\/_0553_ ), .D(\u0\/u3\/_0555_ ), .X(\u0\/u3\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1338_ ( .A(\u0\/u3\/_0528_ ), .B(\u0\/u3\/_0535_ ), .C(\u0\/u3\/_0548_ ), .D(\u0\/u3\/_0556_ ), .X(\u0\/u3\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u3/_1339_ ( .A(\u0\/u3\/_0504_ ), .B(\u0\/u3\/_0519_ ), .C(\u0\/u3\/_0557_ ), .Y(\u0\/u3\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1340_ ( .A(\u0\/u3\/_0054_ ), .B(\u0\/u3\/_0507_ ), .X(\u0\/u3\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u3/_1341_ ( .A_N(\u0\/u3\/_0558_ ), .B(\u0\/u3\/_0408_ ), .C(\u0\/u3\/_0451_ ), .D(\u0\/u3\/_0452_ ), .X(\u0\/u3\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1342_ ( .A(\u0\/u3\/_0549_ ), .Y(\u0\/u3\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1343_ ( .A(\u0\/u3\/_0559_ ), .B(\u0\/u3\/_0403_ ), .C(\u0\/u3\/_0560_ ), .D(\u0\/u3\/_0371_ ), .X(\u0\/u3\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1344_ ( .A(\u0\/u3\/_0181_ ), .B(\u0\/u3\/_0178_ ), .X(\u0\/u3\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1345_ ( .A(\u0\/u3\/_0562_ ), .B(\u0\/u3\/_0552_ ), .C(\u0\/u3\/_0553_ ), .D(\u0\/u3\/_0555_ ), .X(\u0\/u3\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1346_ ( .A(\u0\/u3\/_0029_ ), .B(\u0\/u3\/_0020_ ), .Y(\u0\/u3\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1347_ ( .A(\u0\/u3\/_0051_ ), .B(\u0\/u3\/_0130_ ), .X(\u0\/u3\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1348_ ( .A(\u0\/u3\/_0566_ ), .Y(\u0\/u3\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1349_ ( .A(\u0\/u3\/_0159_ ), .B(\u0\/u3\/_0412_ ), .X(\u0\/u3\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1350_ ( .A1(\u0\/u3\/_0752_ ), .A2(\u0\/u3\/_0640_ ), .B1(\u0\/u3\/_0568_ ), .B2(\u0\/u3\/_0175_ ), .Y(\u0\/u3\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1351_ ( .A(\u0\/u3\/_0076_ ), .B(\u0\/u3\/_0565_ ), .C(\u0\/u3\/_0567_ ), .D(\u0\/u3\/_0569_ ), .X(\u0\/u3\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u3/_1352_ ( .A1(\u0\/u3\/_0035_ ), .A2(\u0\/u3\/_0142_ ), .B1(\u0\/u3\/_0161_ ), .X(\u0\/u3\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1353_ ( .A(\u0\/u3\/_0364_ ), .B(\u0\/u3\/_0662_ ), .Y(\u0\/u3\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u3/_1354_ ( .A(\u0\/u3\/_0420_ ), .B(\u0\/u3\/_0571_ ), .C_N(\u0\/u3\/_0572_ ), .Y(\u0\/u3\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1355_ ( .A(\u0\/u3\/_0051_ ), .B(\u0\/u3\/_0746_ ), .Y(\u0\/u3\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1356_ ( .A(\u0\/u3\/_0574_ ), .B(\u0\/u3\/_0319_ ), .C(\u0\/u3\/_0320_ ), .D(\u0\/u3\/_0411_ ), .X(\u0\/u3\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1357_ ( .A(\u0\/u3\/_0736_ ), .B(\u0\/u3\/_0035_ ), .Y(\u0\/u3\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1358_ ( .A(\u0\/u3\/_0736_ ), .B(\u0\/u3\/_0030_ ), .Y(\u0\/u3\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1359_ ( .A(\u0\/u3\/_0298_ ), .B(\u0\/u3\/_0208_ ), .C(\u0\/u3\/_0577_ ), .D(\u0\/u3\/_0578_ ), .X(\u0\/u3\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1360_ ( .A1(\u0\/u3\/_0020_ ), .A2(\u0\/u3\/_0137_ ), .B1(\u0\/u3\/_0261_ ), .B2(\u0\/u3\/_0128_ ), .Y(\u0\/u3\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1361_ ( .A(\u0\/u3\/_0573_ ), .B(\u0\/u3\/_0576_ ), .C(\u0\/u3\/_0579_ ), .D(\u0\/u3\/_0580_ ), .X(\u0\/u3\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1362_ ( .A(\u0\/u3\/_0561_ ), .B(\u0\/u3\/_0563_ ), .C(\u0\/u3\/_0570_ ), .D(\u0\/u3\/_0581_ ), .X(\u0\/u3\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1363_ ( .A(\u0\/u3\/_0128_ ), .B(\u0\/u3\/_0193_ ), .X(\u0\/u3\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1364_ ( .A(\u0\/u3\/_0082_ ), .B(\u0\/u3\/_0162_ ), .X(\u0\/u3\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u3/_1365_ ( .A(\u0\/u3\/_0583_ ), .B(\u0\/u3\/_0584_ ), .C_N(\u0\/u3\/_0437_ ), .Y(\u0\/u3\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u3/_1366_ ( .A(\u0\/u3\/_0150_ ), .B(\u0\/u3\/_0118_ ), .C(\u0\/u3\/_0380_ ), .Y(\u0\/u3\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u3/_1367_ ( .A_N(\u0\/u3\/_0182_ ), .B(\u0\/u3\/_0587_ ), .C(\u0\/u3\/_0323_ ), .X(\u0\/u3\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1368_ ( .A1(\u0\/u3\/_0575_ ), .A2(\u0\/u3\/_0153_ ), .B1(\u0\/u3\/_0727_ ), .B2(\u0\/u3\/_0058_ ), .Y(\u0\/u3\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1369_ ( .A1(\u0\/u3\/_0218_ ), .A2(\u0\/u3\/_0064_ ), .B1(\u0\/u3\/_0134_ ), .B2(\u0\/u3\/_0255_ ), .Y(\u0\/u3\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1370_ ( .A(\u0\/u3\/_0585_ ), .B(\u0\/u3\/_0588_ ), .C(\u0\/u3\/_0589_ ), .D(\u0\/u3\/_0590_ ), .X(\u0\/u3\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \u0/u3/_1371_ ( .A1(\u0\/u3\/_0091_ ), .A2(\u0\/u3\/_0139_ ), .B1(\u0\/u3\/_0250_ ), .Y(\u0\/u3\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1372_ ( .A1(\u0\/u3\/_0092_ ), .A2(\u0\/u3\/_0739_ ), .B1(\u0\/u3\/_0324_ ), .B2(\u0\/u3\/_0029_ ), .Y(\u0\/u3\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1373_ ( .A1(\u0\/u3\/_0144_ ), .A2(\u0\/u3\/_0153_ ), .B1(\u0\/u3\/_0683_ ), .B2(\u0\/u3\/_0292_ ), .Y(\u0\/u3\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1374_ ( .A1(\u0\/u3\/_0091_ ), .A2(\u0\/u3\/_0218_ ), .B1(\u0\/u3\/_0330_ ), .B2(\u0\/u3\/_0292_ ), .Y(\u0\/u3\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1375_ ( .A(\u0\/u3\/_0592_ ), .B(\u0\/u3\/_0593_ ), .C(\u0\/u3\/_0594_ ), .D(\u0\/u3\/_0595_ ), .X(\u0\/u3\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1376_ ( .A(\u0\/u3\/_0218_ ), .B(\u0\/u3\/_0144_ ), .Y(\u0\/u3\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1377_ ( .A(\u0\/u3\/_0312_ ), .B(\u0\/u3\/_0598_ ), .Y(\u0\/u3\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1378_ ( .A(\u0\/u3\/_0575_ ), .B(\u0\/u3\/_0147_ ), .Y(\u0\/u3\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1379_ ( .A1(\u0\/u3\/_0293_ ), .A2(\u0\/u3\/_0137_ ), .B1(\u0\/u3\/_0093_ ), .B2(\u0\/u3\/_0739_ ), .Y(\u0\/u3\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1380_ ( .A1(\u0\/u3\/_0734_ ), .A2(\u0\/u3\/_0531_ ), .B1(\u0\/u3\/_0600_ ), .C1(\u0\/u3\/_0601_ ), .Y(\u0\/u3\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1381_ ( .A1(\u0\/u3\/_0153_ ), .A2(\u0\/u3\/_0261_ ), .B1(\u0\/u3\/_0599_ ), .C1(\u0\/u3\/_0602_ ), .Y(\u0\/u3\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1382_ ( .A(\u0\/u3\/_0591_ ), .B(\u0\/u3\/_0596_ ), .C(\u0\/u3\/_0174_ ), .D(\u0\/u3\/_0603_ ), .X(\u0\/u3\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1383_ ( .A(\u0\/u3\/_0029_ ), .B(\u0\/u3\/_0144_ ), .Y(\u0\/u3\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1384_ ( .A(\u0\/u3\/_0113_ ), .B(\u0\/u3\/_0017_ ), .Y(\u0\/u3\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1385_ ( .A(\u0\/u3\/_0381_ ), .B(\u0\/u3\/_0605_ ), .C(\u0\/u3\/_0361_ ), .D(\u0\/u3\/_0606_ ), .X(\u0\/u3\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1386_ ( .A1(\u0\/u3\/_0016_ ), .A2(\u0\/u3\/_0727_ ), .B1(\u0\/u3\/_0733_ ), .Y(\u0\/u3\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1387_ ( .A1(\u0\/u3\/_0586_ ), .A2(\u0\/u3\/_0159_ ), .B1(\u0\/u3\/_0082_ ), .B2(\u0\/u3\/_0750_ ), .Y(\u0\/u3\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1388_ ( .A1(\u0\/u3\/_0142_ ), .A2(\u0\/u3\/_0162_ ), .B1(\u0\/u3\/_0079_ ), .B2(\u0\/u3\/_0054_ ), .Y(\u0\/u3\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1389_ ( .A(\u0\/u3\/_0610_ ), .B(\u0\/u3\/_0611_ ), .C(\u0\/u3\/_0105_ ), .D(\u0\/u3\/_0106_ ), .X(\u0\/u3\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1390_ ( .A1(\u0\/u3\/_0094_ ), .A2(\u0\/u3\/_0302_ ), .B1(\u0\/u3\/_0324_ ), .B2(\u0\/u3\/_0089_ ), .Y(\u0\/u3\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1391_ ( .A(\u0\/u3\/_0607_ ), .B(\u0\/u3\/_0609_ ), .C(\u0\/u3\/_0612_ ), .D(\u0\/u3\/_0613_ ), .X(\u0\/u3\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1392_ ( .A(\u0\/u3\/_0041_ ), .B(\u0\/u3\/_0170_ ), .X(\u0\/u3\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1393_ ( .A(\u0\/u3\/_0554_ ), .B(\u0\/u3\/_0027_ ), .X(\u0\/u3\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1394_ ( .A(\u0\/u3\/_0027_ ), .B(\u0\/u3\/_0261_ ), .Y(\u0\/u3\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u3/_1395_ ( .A_N(\u0\/u3\/_0616_ ), .B(\u0\/u3\/_0617_ ), .Y(\u0\/u3\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1396_ ( .A1(\u0\/u3\/_0147_ ), .A2(\u0\/u3\/_0302_ ), .B1(\u0\/u3\/_0342_ ), .C1(\u0\/u3\/_0618_ ), .Y(\u0\/u3\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1397_ ( .A(\u0\/u3\/_0614_ ), .B(\u0\/u3\/_0272_ ), .C(\u0\/u3\/_0615_ ), .D(\u0\/u3\/_0620_ ), .X(\u0\/u3\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u3/_1398_ ( .A(\u0\/u3\/_0582_ ), .B(\u0\/u3\/_0604_ ), .C(\u0\/u3\/_0621_ ), .Y(\u0\/u3\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1399_ ( .A1(\u0\/u3\/_0084_ ), .A2(\u0\/u3\/_0134_ ), .B1(\u0\/u3\/_0089_ ), .Y(\u0\/u3\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1400_ ( .A1(\u0\/u3\/_0144_ ), .A2(\u0\/u3\/_0608_ ), .A3(\u0\/u3\/_0330_ ), .B1(\u0\/u3\/_0089_ ), .Y(\u0\/u3\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1401_ ( .A1(\u0\/u3\/_0197_ ), .A2(\u0\/u3\/_0130_ ), .A3(\u0\/u3\/_0110_ ), .B1(\u0\/u3\/_0094_ ), .Y(\u0\/u3\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1402_ ( .A(\u0\/u3\/_0432_ ), .B(\u0\/u3\/_0622_ ), .C(\u0\/u3\/_0623_ ), .D(\u0\/u3\/_0624_ ), .X(\u0\/u3\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \u0/u3/_1403_ ( .A1(\u0\/u3\/_0554_ ), .A2(\u0\/u3\/_0017_ ), .A3(\u0\/u3\/_0022_ ), .B1(\u0\/u3\/_0161_ ), .X(\u0\/u3\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u3/_1404_ ( .A_N(\u0\/u3\/_0269_ ), .B(\u0\/u3\/_0170_ ), .X(\u0\/u3\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1405_ ( .A1(\u0\/u3\/_0109_ ), .A2(\u0\/u3\/_0064_ ), .A3(\u0\/u3\/_0733_ ), .B1(\u0\/u3\/_0355_ ), .Y(\u0\/u3\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u3/_1406_ ( .A_N(\u0\/u3\/_0626_ ), .B(\u0\/u3\/_0627_ ), .C(\u0\/u3\/_0353_ ), .D(\u0\/u3\/_0628_ ), .X(\u0\/u3\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1407_ ( .A1(\u0\/u3\/_0091_ ), .A2(\u0\/u3\/_0110_ ), .A3(\u0\/u3\/_0176_ ), .B1(\u0\/u3\/_0139_ ), .Y(\u0\/u3\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1408_ ( .A1(\u0\/u3\/_0020_ ), .A2(\u0\/u3\/_0261_ ), .B1(\u0\/u3\/_0147_ ), .Y(\u0\/u3\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1409_ ( .A(\u0\/u3\/_0631_ ), .B(\u0\/u3\/_0344_ ), .C(\u0\/u3\/_0421_ ), .D(\u0\/u3\/_0632_ ), .X(\u0\/u3\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u3/_1410_ ( .A1(\u0\/u3\/_0325_ ), .A2(\u0\/u3\/_0734_ ), .B1(\u0\/u3\/_0038_ ), .C1(\u0\/u3\/_0113_ ), .X(\u0\/u3\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1411_ ( .A1(\u0\/u3\/_0134_ ), .A2(\u0\/u3\/_0114_ ), .B1(\u0\/u3\/_0221_ ), .C1(\u0\/u3\/_0634_ ), .Y(\u0\/u3\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \u0/u3/_1412_ ( .A(\u0\/u3\/_0119_ ), .B_N(\u0\/u3\/_0111_ ), .Y(\u0\/u3\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1413_ ( .A1(\u0\/u3\/_0032_ ), .A2(\u0\/u3\/_0113_ ), .B1(\u0\/u3\/_0636_ ), .C1(\u0\/u3\/_0400_ ), .Y(\u0\/u3\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1414_ ( .A1(\u0\/u3\/_0731_ ), .A2(\u0\/u3\/_0293_ ), .A3(\u0\/u3\/_0251_ ), .B1(\u0\/u3\/_0364_ ), .Y(\u0\/u3\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1415_ ( .A(\u0\/u3\/_0189_ ), .B(\u0\/u3\/_0635_ ), .C(\u0\/u3\/_0637_ ), .D(\u0\/u3\/_0638_ ), .X(\u0\/u3\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1416_ ( .A(\u0\/u3\/_0625_ ), .B(\u0\/u3\/_0630_ ), .C(\u0\/u3\/_0633_ ), .D(\u0\/u3\/_0639_ ), .X(\u0\/u3\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1417_ ( .A(\u0\/u3\/_0746_ ), .B(\u0\/u3\/_0738_ ), .X(\u0\/u3\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1418_ ( .A(\u0\/u3\/_0736_ ), .B(\u0\/u3\/_0731_ ), .X(\u0\/u3\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \u0/u3/_1419_ ( .A_N(\u0\/u3\/_0643_ ), .B(\u0\/u3\/_0577_ ), .Y(\u0\/u3\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1420_ ( .A1(\u0\/u3\/_0084_ ), .A2(\u0\/u3\/_0739_ ), .B1(\u0\/u3\/_0642_ ), .C1(\u0\/u3\/_0644_ ), .Y(\u0\/u3\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1421_ ( .A1(\u0\/u3\/_0050_ ), .A2(\u0\/u3\/_0249_ ), .B1(\u0\/u3\/_0194_ ), .C1(\u0\/u3\/_0738_ ), .Y(\u0\/u3\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1422_ ( .A(\u0\/u3\/_0646_ ), .B(\u0\/u3\/_0232_ ), .C(\u0\/u3\/_0417_ ), .D(\u0\/u3\/_0578_ ), .X(\u0\/u3\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1423_ ( .A1(\u0\/u3\/_0064_ ), .A2(\u0\/u3\/_0733_ ), .B1(\u0\/u3\/_0727_ ), .Y(\u0\/u3\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1424_ ( .A1(\u0\/u3\/_0193_ ), .A2(\u0\/u3\/_0276_ ), .B1(\u0\/u3\/_0727_ ), .Y(\u0\/u3\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1425_ ( .A(\u0\/u3\/_0645_ ), .B(\u0\/u3\/_0647_ ), .C(\u0\/u3\/_0648_ ), .D(\u0\/u3\/_0649_ ), .X(\u0\/u3\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1426_ ( .A1(\u0\/u3\/_0325_ ), .A2(\u0\/u3\/_0734_ ), .B1(\u0\/u3\/_0038_ ), .C1(\u0\/u3\/_0029_ ), .Y(\u0\/u3\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1427_ ( .A1(\u0\/u3\/_0249_ ), .A2(\u0\/u3\/_0216_ ), .B1(\u0\/u3\/_0412_ ), .C1(\u0\/u3\/_0029_ ), .Y(\u0\/u3\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1428_ ( .A(\u0\/u3\/_0652_ ), .B(\u0\/u3\/_0653_ ), .X(\u0\/u3\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1429_ ( .A1(\u0\/u3\/_0733_ ), .A2(\u0\/u3\/_0748_ ), .A3(\u0\/u3\/_0324_ ), .B1(\u0\/u3\/_0016_ ), .Y(\u0\/u3\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1430_ ( .A1(\u0\/u3\/_0640_ ), .A2(\u0\/u3\/_0193_ ), .A3(\u0\/u3\/_0091_ ), .B1(\u0\/u3\/_0016_ ), .Y(\u0\/u3\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1431_ ( .A1(\u0\/u3\/_0102_ ), .A2(\u0\/u3\/_0301_ ), .B1(\w3\[27\] ), .C1(\u0\/u3\/_0029_ ), .Y(\u0\/u3\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1432_ ( .A(\u0\/u3\/_0654_ ), .B(\u0\/u3\/_0655_ ), .C(\u0\/u3\/_0656_ ), .D(\u0\/u3\/_0657_ ), .X(\u0\/u3\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1433_ ( .A1(\u0\/u3\/_0118_ ), .A2(\u0\/u3\/_0050_ ), .B1(\u0\/u3\/_0038_ ), .C1(\u0\/u3\/_0478_ ), .Y(\u0\/u3\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \u0/u3/_1434_ ( .A_N(\u0\/u3\/_0250_ ), .B(\u0\/u3\/_0465_ ), .C(\u0\/u3\/_0659_ ), .X(\u0\/u3\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1435_ ( .A1(\u0\/u3\/_0683_ ), .A2(\u0\/u3\/_0324_ ), .B1(\u0\/u3\/_0255_ ), .Y(\u0\/u3\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1436_ ( .A1(\u0\/u3\/_0032_ ), .A2(\u0\/u3\/_0193_ ), .A3(\u0\/u3\/_0047_ ), .B1(\u0\/u3\/_0255_ ), .Y(\u0\/u3\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1437_ ( .A1(\u0\/u3\/_0144_ ), .A2(\u0\/u3\/_0586_ ), .A3(\u0\/u3\/_0047_ ), .B1(\u0\/u3\/_0218_ ), .Y(\u0\/u3\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1438_ ( .A(\u0\/u3\/_0660_ ), .B(\u0\/u3\/_0661_ ), .C(\u0\/u3\/_0663_ ), .D(\u0\/u3\/_0664_ ), .X(\u0\/u3\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1439_ ( .A1(\u0\/u3\/_0091_ ), .A2(\u0\/u3\/_0276_ ), .B1(\u0\/u3\/_0060_ ), .Y(\u0\/u3\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1440_ ( .A1(\u0\/u3\/_0144_ ), .A2(\u0\/u3\/_0608_ ), .B1(\u0\/u3\/_0292_ ), .Y(\u0\/u3\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1441_ ( .A1(\u0\/u3\/_0412_ ), .A2(\u0\/u3\/_0038_ ), .B1(\u0\/u3\/_0102_ ), .C1(\u0\/u3\/_0060_ ), .Y(\u0\/u3\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1442_ ( .A1(\w3\[25\] ), .A2(\u0\/u3\/_0734_ ), .B1(\u0\/u3\/_0109_ ), .C1(\u0\/u3\/_0292_ ), .Y(\u0\/u3\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1443_ ( .A(\u0\/u3\/_0666_ ), .B(\u0\/u3\/_0667_ ), .C(\u0\/u3\/_0668_ ), .D(\u0\/u3\/_0669_ ), .X(\u0\/u3\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1444_ ( .A(\u0\/u3\/_0650_ ), .B(\u0\/u3\/_0658_ ), .C(\u0\/u3\/_0665_ ), .D(\u0\/u3\/_0670_ ), .X(\u0\/u3\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u3/_1445_ ( .A(\u0\/u3\/_0641_ ), .B(\u0\/u3\/_0174_ ), .C(\u0\/u3\/_0671_ ), .Y(\u0\/u3\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \u0/u3/_1446_ ( .A(\u0\/u3\/_0049_ ), .B(\u0\/u3\/_0618_ ), .C_N(\u0\/u3\/_0052_ ), .Y(\u0\/u3\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \u0/u3/_1447_ ( .A(\u0\/u3\/_0239_ ), .Y(\u0\/u3\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1448_ ( .A(\u0\/u3\/_0705_ ), .B(\u0\/u3\/_0032_ ), .Y(\u0\/u3\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1449_ ( .A1(\u0\/u3\/_0054_ ), .A2(\u0\/u3\/_0731_ ), .B1(\u0\/u3\/_0035_ ), .B2(\u0\/u3\/_0705_ ), .Y(\u0\/u3\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1450_ ( .A1(\u0\/u3\/_0304_ ), .A2(\u0\/u3\/_0731_ ), .B1(\u0\/u3\/_0047_ ), .B2(\u0\/u3\/_0750_ ), .Y(\u0\/u3\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1451_ ( .A(\u0\/u3\/_0674_ ), .B(\u0\/u3\/_0675_ ), .C(\u0\/u3\/_0676_ ), .D(\u0\/u3\/_0677_ ), .X(\u0\/u3\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \u0/u3/_1452_ ( .A_N(\u0\/u3\/_0584_ ), .B(\u0\/u3\/_0283_ ), .X(\u0\/u3\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1453_ ( .A(\u0\/u3\/_0673_ ), .B(\u0\/u3\/_0678_ ), .C(\u0\/u3\/_0679_ ), .D(\u0\/u3\/_0508_ ), .X(\u0\/u3\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1454_ ( .A1(\u0\/u3\/_0016_ ), .A2(\u0\/u3\/_0733_ ), .B1(\u0\/u3\/_0355_ ), .B2(\u0\/u3\/_0092_ ), .Y(\u0\/u3\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1455_ ( .A(\u0\/u3\/_0681_ ), .B(\u0\/u3\/_0034_ ), .X(\u0\/u3\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u3/_1456_ ( .A1(\u0\/u3\/_0330_ ), .A2(\u0\/u3\/_0139_ ), .B1(\u0\/u3\/_0324_ ), .B2(\u0\/u3\/_0089_ ), .X(\u0\/u3\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1457_ ( .A1(\u0\/u3\/_0146_ ), .A2(\u0\/u3\/_0147_ ), .B1(\u0\/u3\/_0133_ ), .C1(\u0\/u3\/_0684_ ), .Y(\u0\/u3\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1458_ ( .A(\u0\/u3\/_0113_ ), .B(\u0\/u3\/_0251_ ), .Y(\u0\/u3\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u3/_1459_ ( .A_N(\u0\/u3\/_0463_ ), .B(\u0\/u3\/_0686_ ), .C(\u0\/u3\/_0383_ ), .D(\u0\/u3\/_0464_ ), .X(\u0\/u3\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1460_ ( .A1(\u0\/u3\/_0051_ ), .A2(\u0\/u3\/_0293_ ), .B1(\u0\/u3\/_0084_ ), .B2(\u0\/u3\/_0705_ ), .Y(\u0\/u3\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1461_ ( .A1(\u0\/u3\/_0017_ ), .A2(\u0\/u3\/_0072_ ), .B1(\u0\/u3\/_0134_ ), .B2(\u0\/u3\/_0078_ ), .Y(\u0\/u3\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1462_ ( .A(\u0\/u3\/_0687_ ), .B(\u0\/u3\/_0236_ ), .C(\u0\/u3\/_0688_ ), .D(\u0\/u3\/_0689_ ), .X(\u0\/u3\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1463_ ( .A(\u0\/u3\/_0680_ ), .B(\u0\/u3\/_0682_ ), .C(\u0\/u3\/_0685_ ), .D(\u0\/u3\/_0690_ ), .X(\u0\/u3\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \u0/u3/_1464_ ( .A1(\u0\/u3\/_0532_ ), .A2(\u0\/u3\/_0380_ ), .B1(\u0\/u3\/_0102_ ), .C1(\u0\/u3\/_0355_ ), .X(\u0\/u3\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u3/_1465_ ( .A(\u0\/u3\/_0692_ ), .B(\u0\/u3\/_0338_ ), .C(\u0\/u3\/_0644_ ), .Y(\u0\/u3\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1466_ ( .A(\u0\/u3\/_0016_ ), .B(\u0\/u3\/_0020_ ), .Y(\u0\/u3\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1467_ ( .A1(\u0\/u3\/_0032_ ), .A2(\u0\/u3\/_0137_ ), .B1(\u0\/u3\/_0279_ ), .B2(\u0\/u3\/_0094_ ), .Y(\u0\/u3\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1468_ ( .A1(\u0\/u3\/_0575_ ), .A2(\u0\/u3\/_0153_ ), .B1(\u0\/u3\/_0161_ ), .B2(\u0\/u3\/_0293_ ), .Y(\u0\/u3\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1469_ ( .A(\u0\/u3\/_0259_ ), .B(\u0\/u3\/_0695_ ), .C(\u0\/u3\/_0696_ ), .D(\u0\/u3\/_0697_ ), .X(\u0\/u3\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u3/_1470_ ( .A1(\u0\/u3\/_0255_ ), .A2(\u0\/u3\/_0640_ ), .B1(\u0\/u3\/_0016_ ), .B2(\u0\/u3\/_0193_ ), .X(\u0\/u3\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1471_ ( .A1(\u0\/u3\/_0060_ ), .A2(\u0\/u3\/_0176_ ), .B1(\u0\/u3\/_0699_ ), .C1(\u0\/u3\/_0177_ ), .Y(\u0\/u3\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1472_ ( .A1(\u0\/u3\/_0091_ ), .A2(\u0\/u3\/_0218_ ), .B1(\u0\/u3\/_0092_ ), .B2(\u0\/u3\/_0705_ ), .Y(\u0\/u3\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \u0/u3/_1473_ ( .A1(\u0\/u3\/_0705_ ), .A2(\u0\/u3\/_0683_ ), .B1(\u0\/u3\/_0093_ ), .B2(\u0\/u3\/_0114_ ), .Y(\u0\/u3\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \u0/u3/_1474_ ( .A1(\u0\/u3\/_0683_ ), .A2(\u0\/u3\/_0084_ ), .B1(\u0\/u3\/_0094_ ), .Y(\u0\/u3\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \u0/u3/_1475_ ( .A1(\u0\/u3\/_0249_ ), .A2(\u0\/u3\/_0216_ ), .B1(\u0\/u3\/_0038_ ), .C1(\u0\/u3\/_0292_ ), .Y(\u0\/u3\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1476_ ( .A(\u0\/u3\/_0701_ ), .B(\u0\/u3\/_0702_ ), .C(\u0\/u3\/_0703_ ), .D(\u0\/u3\/_0704_ ), .X(\u0\/u3\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1477_ ( .A(\u0\/u3\/_0693_ ), .B(\u0\/u3\/_0698_ ), .C(\u0\/u3\/_0700_ ), .D(\u0\/u3\/_0706_ ), .X(\u0\/u3\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u3/_1478_ ( .A1(\u0\/u3\/_0113_ ), .A2(\u0\/u3\/_0640_ ), .B1(\u0\/u3\/_0364_ ), .B2(\u0\/u3\/_0058_ ), .X(\u0\/u3\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \u0/u3/_1479_ ( .A(\u0\/u3\/_0407_ ), .B(\u0\/u3\/_0708_ ), .C(\u0\/u3\/_0529_ ), .Y(\u0\/u3\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1480_ ( .A(\u0\/u3\/_0568_ ), .B(\u0\/u3\/_0175_ ), .Y(\u0\/u3\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \u0/u3/_1481_ ( .A1(\u0\/u3\/_0029_ ), .A2(\u0\/u3\/_0114_ ), .A3(\u0\/u3\/_0051_ ), .B1(\u0\/u3\/_0130_ ), .Y(\u0\/u3\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1482_ ( .A(\u0\/u3\/_0709_ ), .B(\u0\/u3\/_0550_ ), .C(\u0\/u3\/_0710_ ), .D(\u0\/u3\/_0711_ ), .X(\u0\/u3\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \u0/u3/_1483_ ( .A1(\u0\/u3\/_0114_ ), .A2(\u0\/u3\/_0064_ ), .B1(\u0\/u3\/_0261_ ), .B2(\u0\/u3\/_0089_ ), .X(\u0\/u3\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1484_ ( .A1(\u0\/u3\/_0355_ ), .A2(\u0\/u3\/_0261_ ), .B1(\u0\/u3\/_0198_ ), .C1(\u0\/u3\/_0713_ ), .Y(\u0\/u3\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1485_ ( .A(\u0\/u3\/_0586_ ), .B(\u0\/u3\/_0478_ ), .Y(\u0\/u3\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u3/_1486_ ( .A_N(\u0\/u3\/_0541_ ), .B(\u0\/u3\/_0267_ ), .C(\u0\/u3\/_0715_ ), .D(\u0\/u3\/_0320_ ), .X(\u0\/u3\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1487_ ( .A(\u0\/u3\/_0586_ ), .B(\u0\/u3\/_0070_ ), .Y(\u0\/u3\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \u0/u3/_1488_ ( .A_N(\u0\/u3\/_0211_ ), .B(\u0\/u3\/_0155_ ), .C(\u0\/u3\/_0202_ ), .D(\u0\/u3\/_0718_ ), .X(\u0\/u3\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u3/_1489_ ( .A(\u0\/u3\/_0150_ ), .B(\u0\/u3\/_0216_ ), .C(\u0\/u3\/_0380_ ), .Y(\u0\/u3\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \u0/u3/_1490_ ( .A(\u0\/u3\/_0411_ ), .B(\u0\/u3\/_0720_ ), .X(\u0\/u3\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \u0/u3/_1491_ ( .A1(\u0\/u3\/_0017_ ), .A2(\u0\/u3\/_0022_ ), .B1(\u0\/u3\/_0078_ ), .X(\u0\/u3\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \u0/u3/_1492_ ( .A1(\u0\/u3\/_0134_ ), .A2(\u0\/u3\/_0738_ ), .B1(\u0\/u3\/_0101_ ), .C1(\u0\/u3\/_0722_ ), .Y(\u0\/u3\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1493_ ( .A(\u0\/u3\/_0717_ ), .B(\u0\/u3\/_0719_ ), .C(\u0\/u3\/_0721_ ), .D(\u0\/u3\/_0723_ ), .X(\u0\/u3\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \u0/u3/_1494_ ( .A(\u0\/u3\/_0739_ ), .B(\u0\/u3\/_0193_ ), .Y(\u0\/u3\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1495_ ( .A(\u0\/u3\/_0344_ ), .B(\u0\/u3\/_0184_ ), .C(\u0\/u3\/_0449_ ), .D(\u0\/u3\/_0725_ ), .X(\u0\/u3\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \u0/u3/_1496_ ( .A(\u0\/u3\/_0712_ ), .B(\u0\/u3\/_0714_ ), .C(\u0\/u3\/_0724_ ), .D(\u0\/u3\/_0726_ ), .X(\u0\/u3\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \u0/u3/_1497_ ( .A(\u0\/u3\/_0691_ ), .B(\u0\/u3\/_0707_ ), .C(\u0\/u3\/_0728_ ), .Y(\u0\/u3\/_0015_ ) );
sky130_fd_sc_hd__clkbuf_1 \u0/u3/_1500_ ( .A(\w3\[31\] ), .X(\u0\/u3\/_0007_ ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__1 ( .HI( ), .LO(net1 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__10 ( .HI( ), .LO(net10 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__11 ( .HI( ), .LO(net11 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__12 ( .HI( ), .LO(net12 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__13 ( .HI( ), .LO(net13 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__14 ( .HI( ), .LO(net14 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__15 ( .HI( ), .LO(net15 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__16 ( .HI( ), .LO(net16 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__17 ( .HI( ), .LO(net17 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__18 ( .HI( ), .LO(net18 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__19 ( .HI( ), .LO(net19 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__2 ( .HI( ), .LO(net2 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__20 ( .HI( ), .LO(net20 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__21 ( .HI( ), .LO(net21 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__22 ( .HI( ), .LO(net22 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__23 ( .HI( ), .LO(net23 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__24 ( .HI( ), .LO(net24 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__25 ( .HI( ), .LO(net25 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__26 ( .HI( ), .LO(net26 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__27 ( .HI( ), .LO(net27 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__28 ( .HI( ), .LO(net28 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__29 ( .HI( ), .LO(net29 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__3 ( .HI( ), .LO(net3 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__30 ( .HI( ), .LO(net30 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__31 ( .HI( ), .LO(net31 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__32 ( .HI( ), .LO(net32 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__33 ( .HI( ), .LO(net33 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__4 ( .HI( ), .LO(net4 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__5 ( .HI( ), .LO(net5 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__6 ( .HI( ), .LO(net6 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__7 ( .HI( ), .LO(net7 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__8 ( .HI( ), .LO(net8 ) );
sky130_fd_sc_hd__conb_1 \u0/r0/_102__9 ( .HI( ), .LO(net9 ) );
sky130_fd_sc_hd__nor2b_1 \us00/_0753_ ( .A(\sa00\[2\] ), .B_N(\sa00\[3\] ), .Y(\us00\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0755_ ( .A(\sa00\[1\] ), .B(\sa00\[0\] ), .X(\us00\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0756_ ( .A(\us00\/_0096_ ), .B(\us00\/_0118_ ), .X(\us00\/_0129_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0757_ ( .A(\sa00\[7\] ), .B(\sa00\[6\] ), .X(\us00\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_0758_ ( .A(\sa00\[4\] ), .B(\sa00\[5\] ), .Y(\us00\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0759_ ( .A(\us00\/_0140_ ), .B(\us00\/_0151_ ), .X(\us00\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0761_ ( .A(\us00\/_0129_ ), .B(\us00\/_0162_ ), .X(\us00\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0762_ ( .A(\us00\/_0096_ ), .X(\us00\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \us00/_0763_ ( .A(\sa00\[1\] ), .B_N(\sa00\[0\] ), .Y(\us00\/_0205_ ) );
sky130_fd_sc_hd__and3_1 \us00/_0765_ ( .A(\us00\/_0162_ ), .B(\us00\/_0194_ ), .C(\us00\/_0205_ ), .X(\us00\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us00/_0766_ ( .A(\us00\/_0183_ ), .SLEEP(\us00\/_0227_ ), .X(\us00\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \us00/_0767_ ( .A(\sa00\[0\] ), .B_N(\sa00\[1\] ), .Y(\us00\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_0768_ ( .A(\sa00\[2\] ), .B(\sa00\[3\] ), .Y(\us00\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0769_ ( .A(\us00\/_0249_ ), .B(\us00\/_0260_ ), .X(\us00\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0771_ ( .A(\us00\/_0271_ ), .X(\us00\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0772_ ( .A(\us00\/_0162_ ), .X(\us00\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_0773_ ( .A(\us00\/_0293_ ), .B(\us00\/_0304_ ), .Y(\us00\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us00/_0774_ ( .A(\sa00\[1\] ), .Y(\us00\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us00/_0776_ ( .A(\sa00\[0\] ), .Y(\us00\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0777_ ( .A(\sa00\[2\] ), .B(\sa00\[3\] ), .X(\us00\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0779_ ( .A(\us00\/_0358_ ), .X(\us00\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_0780_ ( .A1(\us00\/_0325_ ), .A2(\us00\/_0347_ ), .B1(\us00\/_0380_ ), .C1(\us00\/_0304_ ), .Y(\us00\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us00/_0781_ ( .A_N(\us00\/_0238_ ), .B(\us00\/_0314_ ), .C(\us00\/_0391_ ), .X(\us00\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us00/_0782_ ( .A(\sa00\[3\] ), .B_N(\sa00\[2\] ), .Y(\us00\/_0412_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0784_ ( .A(\us00\/_0412_ ), .B(\us00\/_0205_ ), .X(\us00\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \us00/_0787_ ( .A(\sa00\[5\] ), .B_N(\sa00\[4\] ), .Y(\us00\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0788_ ( .A(\us00\/_0467_ ), .B(\us00\/_0140_ ), .X(\us00\/_0478_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_0791_ ( .A(\us00\/_0134_ ), .B(\us00\/_0218_ ), .Y(\us00\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_0792_ ( .A(\us00\/_0478_ ), .B(\us00\/_0271_ ), .Y(\us00\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0793_ ( .A(\us00\/_0194_ ), .X(\us00\/_0532_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0795_ ( .A(\us00\/_0249_ ), .B(\us00\/_0358_ ), .X(\us00\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0797_ ( .A(\us00\/_0554_ ), .X(\us00\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0798_ ( .A(\us00\/_0205_ ), .B(\us00\/_0358_ ), .X(\us00\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0800_ ( .A(\us00\/_0586_ ), .X(\us00\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_0801_ ( .A1(\us00\/_0532_ ), .A2(\us00\/_0575_ ), .A3(\us00\/_0608_ ), .B1(\us00\/_0218_ ), .Y(\us00\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us00/_0802_ ( .A(\us00\/_0401_ ), .B(\us00\/_0510_ ), .C(\us00\/_0521_ ), .D(\us00\/_0619_ ), .X(\us00\/_0629_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0803_ ( .A(\us00\/_0358_ ), .B(\sa00\[1\] ), .X(\us00\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0805_ ( .A(\us00\/_0205_ ), .B(\us00\/_0260_ ), .X(\us00\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0807_ ( .A(\us00\/_0662_ ), .X(\us00\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us00/_0808_ ( .A(\sa00\[6\] ), .B_N(\sa00\[7\] ), .Y(\us00\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0809_ ( .A(\us00\/_0467_ ), .B(\us00\/_0694_ ), .X(\us00\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0811_ ( .A(\us00\/_0705_ ), .X(\us00\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_0812_ ( .A1(\us00\/_0640_ ), .A2(\us00\/_0293_ ), .A3(\us00\/_0683_ ), .B1(\us00\/_0727_ ), .Y(\us00\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_0813_ ( .A(\sa00\[1\] ), .B(\sa00\[0\] ), .Y(\us00\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0814_ ( .A(\us00\/_0730_ ), .B(\us00\/_0260_ ), .X(\us00\/_0731_ ) );
sky130_fd_sc_hd__buf_1 \us00/_0815_ ( .A(\us00\/_0731_ ), .X(\us00\/_0732_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0816_ ( .A(\us00\/_0732_ ), .X(\us00\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0817_ ( .A(\sa00\[0\] ), .X(\us00\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us00/_0818_ ( .A1(\us00\/_0325_ ), .A2(\us00\/_0734_ ), .B1(\us00\/_0412_ ), .X(\us00\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0819_ ( .A(\us00\/_0694_ ), .B(\us00\/_0151_ ), .X(\us00\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0821_ ( .A(\us00\/_0736_ ), .X(\us00\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0822_ ( .A(\us00\/_0738_ ), .X(\us00\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_0823_ ( .A1(\us00\/_0733_ ), .A2(\us00\/_0735_ ), .A3(\us00\/_0293_ ), .B1(\us00\/_0739_ ), .Y(\us00\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us00/_0824_ ( .A(\us00\/_0730_ ), .B_N(\us00\/_0358_ ), .Y(\us00\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_0825_ ( .A(\us00\/_0741_ ), .B(\us00\/_0739_ ), .Y(\us00\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_0827_ ( .A1(\us00\/_0118_ ), .A2(\us00\/_0205_ ), .B1(\us00\/_0532_ ), .C1(\us00\/_0739_ ), .Y(\us00\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us00/_0828_ ( .A(\us00\/_0729_ ), .B(\us00\/_0740_ ), .C(\us00\/_0742_ ), .D(\us00\/_0744_ ), .X(\us00\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0829_ ( .A(\us00\/_0412_ ), .B(\us00\/_0730_ ), .X(\us00\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0830_ ( .A(\us00\/_0746_ ), .X(\us00\/_0747_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0831_ ( .A(\us00\/_0747_ ), .X(\us00\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us00/_0832_ ( .A(\sa00\[4\] ), .B_N(\sa00\[5\] ), .Y(\us00\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0833_ ( .A(\us00\/_0749_ ), .B(\us00\/_0694_ ), .X(\us00\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0835_ ( .A(\us00\/_0750_ ), .X(\us00\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0836_ ( .A(\us00\/_0752_ ), .X(\us00\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0837_ ( .A(\us00\/_0118_ ), .B(\us00\/_0358_ ), .X(\us00\/_0017_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0839_ ( .A(\us00\/_0752_ ), .B(\us00\/_0017_ ), .X(\us00\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0840_ ( .A(\us00\/_0358_ ), .B(\us00\/_0325_ ), .X(\us00\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0842_ ( .A(\us00\/_0096_ ), .B(\us00\/_0205_ ), .X(\us00\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \us00/_0844_ ( .A1(\us00\/_0020_ ), .A2(\us00\/_0022_ ), .B1(\us00\/_0752_ ), .X(\us00\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_0845_ ( .A1(\us00\/_0748_ ), .A2(\us00\/_0016_ ), .B1(\us00\/_0019_ ), .C1(\us00\/_0024_ ), .Y(\us00\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0846_ ( .A(\sa00\[4\] ), .B(\sa00\[5\] ), .X(\us00\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0847_ ( .A(\us00\/_0694_ ), .B(\us00\/_0026_ ), .X(\us00\/_0027_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0850_ ( .A(\us00\/_0358_ ), .B(\us00\/_0730_ ), .X(\us00\/_0030_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0852_ ( .A(\us00\/_0030_ ), .X(\us00\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_0853_ ( .A(\us00\/_0247_ ), .B(\us00\/_0032_ ), .Y(\us00\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_0854_ ( .A(\us00\/_0247_ ), .B(\us00\/_0735_ ), .Y(\us00\/_0034_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0855_ ( .A(\us00\/_0118_ ), .B(\us00\/_0260_ ), .X(\us00\/_0035_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0857_ ( .A(\us00\/_0027_ ), .B(\us00\/_0035_ ), .X(\us00\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0858_ ( .A(\us00\/_0260_ ), .X(\us00\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_0859_ ( .A(\us00\/_0038_ ), .B(\us00\/_0347_ ), .Y(\us00\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us00/_0860_ ( .A_N(\us00\/_0039_ ), .B(\us00\/_0027_ ), .X(\us00\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_0861_ ( .A(\us00\/_0037_ ), .B(\us00\/_0040_ ), .Y(\us00\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us00/_0862_ ( .A(\us00\/_0025_ ), .B(\us00\/_0033_ ), .C(\us00\/_0034_ ), .D(\us00\/_0041_ ), .X(\us00\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0863_ ( .A(\us00\/_0749_ ), .B(\us00\/_0140_ ), .X(\us00\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us00/_0865_ ( .A(\sa00\[0\] ), .B(\sa00\[2\] ), .C(\sa00\[3\] ), .X(\us00\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0866_ ( .A(\us00\/_0043_ ), .B(\us00\/_0045_ ), .X(\us00\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0867_ ( .A(\us00\/_0096_ ), .B(\us00\/_0249_ ), .X(\us00\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0869_ ( .A(\us00\/_0047_ ), .B(\us00\/_0043_ ), .X(\us00\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0870_ ( .A(\us00\/_0730_ ), .X(\us00\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0871_ ( .A(\us00\/_0043_ ), .X(\us00\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_0872_ ( .A1(\us00\/_0118_ ), .A2(\us00\/_0050_ ), .B1(\us00\/_0194_ ), .C1(\us00\/_0051_ ), .Y(\us00\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us00/_0873_ ( .A(\us00\/_0046_ ), .B(\us00\/_0049_ ), .C_N(\us00\/_0052_ ), .Y(\us00\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0874_ ( .A(\us00\/_0026_ ), .B(\us00\/_0140_ ), .X(\us00\/_0054_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_0877_ ( .A1(\us00\/_0532_ ), .A2(\us00\/_0575_ ), .B1(\us00\/_0292_ ), .Y(\us00\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0878_ ( .A(\us00\/_0412_ ), .B(\us00\/_0325_ ), .X(\us00\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0880_ ( .A(\us00\/_0051_ ), .X(\us00\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_0881_ ( .A1(\us00\/_0732_ ), .A2(\us00\/_0035_ ), .A3(\us00\/_0058_ ), .B1(\us00\/_0060_ ), .Y(\us00\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0882_ ( .A(\us00\/_0260_ ), .B(\sa00\[1\] ), .X(\us00\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0884_ ( .A(\us00\/_0062_ ), .X(\us00\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_0885_ ( .A1(\us00\/_0064_ ), .A2(\us00\/_0748_ ), .A3(\us00\/_0683_ ), .B1(\us00\/_0292_ ), .Y(\us00\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us00/_0886_ ( .A(\us00\/_0053_ ), .B(\us00\/_0057_ ), .C(\us00\/_0061_ ), .D(\us00\/_0065_ ), .X(\us00\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us00/_0887_ ( .A(\us00\/_0629_ ), .B(\us00\/_0745_ ), .C(\us00\/_0042_ ), .D(\us00\/_0066_ ), .X(\us00\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us00/_0889_ ( .A(\sa00\[7\] ), .B_N(\sa00\[6\] ), .Y(\us00\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0890_ ( .A(\us00\/_0069_ ), .B(\us00\/_0151_ ), .X(\us00\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0892_ ( .A(\us00\/_0070_ ), .X(\us00\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_0893_ ( .A1(\us00\/_0129_ ), .A2(\us00\/_0586_ ), .B1(\us00\/_0072_ ), .Y(\us00\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_0894_ ( .A1(\us00\/_0380_ ), .A2(\us00\/_0347_ ), .B1(\us00\/_0194_ ), .B2(\us00\/_0205_ ), .Y(\us00\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us00/_0895_ ( .A(\us00\/_0074_ ), .B_N(\us00\/_0070_ ), .Y(\us00\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us00/_0896_ ( .A(\us00\/_0073_ ), .SLEEP(\us00\/_0075_ ), .X(\us00\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0897_ ( .A(\us00\/_0467_ ), .B(\us00\/_0069_ ), .X(\us00\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0898_ ( .A(\us00\/_0077_ ), .X(\us00\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0899_ ( .A(\us00\/_0412_ ), .B(\us00\/_0118_ ), .X(\us00\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0901_ ( .A(\us00\/_0078_ ), .B(\us00\/_0079_ ), .X(\us00\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0902_ ( .A(\us00\/_0412_ ), .B(\us00\/_0249_ ), .X(\us00\/_0082_ ) );
sky130_fd_sc_hd__buf_2 \us00/_0904_ ( .A(\us00\/_0082_ ), .X(\us00\/_0084_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0905_ ( .A(\us00\/_0084_ ), .B(\us00\/_0078_ ), .X(\us00\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us00/_0906_ ( .A1(\sa00\[0\] ), .A2(\us00\/_0325_ ), .B1(\us00\/_0260_ ), .Y(\us00\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us00/_0907_ ( .A_N(\us00\/_0086_ ), .B(\us00\/_0078_ ), .X(\us00\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us00/_0908_ ( .A(\us00\/_0081_ ), .B(\us00\/_0085_ ), .C(\us00\/_0087_ ), .Y(\us00\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0909_ ( .A(\us00\/_0072_ ), .X(\us00\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_0910_ ( .A1(\us00\/_0733_ ), .A2(\us00\/_0748_ ), .A3(\us00\/_0683_ ), .B1(\us00\/_0089_ ), .Y(\us00\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0911_ ( .A(\us00\/_0129_ ), .X(\us00\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0912_ ( .A(\us00\/_0017_ ), .X(\us00\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0913_ ( .A(\us00\/_0022_ ), .X(\us00\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0914_ ( .A(\us00\/_0078_ ), .X(\us00\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_0915_ ( .A1(\us00\/_0091_ ), .A2(\us00\/_0092_ ), .A3(\us00\/_0093_ ), .B1(\us00\/_0094_ ), .Y(\us00\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us00/_0916_ ( .A(\us00\/_0076_ ), .B(\us00\/_0088_ ), .C(\us00\/_0090_ ), .D(\us00\/_0095_ ), .X(\us00\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0917_ ( .A(\us00\/_0069_ ), .B(\us00\/_0026_ ), .X(\us00\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \us00/_0918_ ( .A(\us00\/_0098_ ), .X(\us00\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0919_ ( .A(\us00\/_0434_ ), .B(\us00\/_0099_ ), .X(\us00\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0920_ ( .A(\us00\/_0079_ ), .B(\us00\/_0098_ ), .X(\us00\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0921_ ( .A(\us00\/_0325_ ), .X(\us00\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_0922_ ( .A1(\us00\/_0102_ ), .A2(\us00\/_0734_ ), .B1(\us00\/_0038_ ), .C1(\us00\/_0099_ ), .Y(\us00\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us00/_0923_ ( .A(\us00\/_0100_ ), .B(\us00\/_0101_ ), .C_N(\us00\/_0103_ ), .Y(\us00\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_0924_ ( .A1(\us00\/_0554_ ), .A2(\us00\/_0586_ ), .B1(\us00\/_0099_ ), .Y(\us00\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_0925_ ( .A(\us00\/_0129_ ), .B(\us00\/_0099_ ), .Y(\us00\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0926_ ( .A(\us00\/_0105_ ), .B(\us00\/_0106_ ), .X(\us00\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0927_ ( .A(\us00\/_0412_ ), .X(\us00\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0928_ ( .A(\us00\/_0260_ ), .B(\sa00\[0\] ), .X(\us00\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0929_ ( .A(\us00\/_0069_ ), .B(\us00\/_0749_ ), .X(\us00\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0931_ ( .A(\us00\/_0111_ ), .X(\us00\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0932_ ( .A(\us00\/_0113_ ), .X(\us00\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_0933_ ( .A1(\us00\/_0109_ ), .A2(\us00\/_0110_ ), .B1(\us00\/_0114_ ), .Y(\us00\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us00/_0934_ ( .A(\us00\/_0022_ ), .Y(\us00\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us00/_0935_ ( .A(\us00\/_0554_ ), .Y(\us00\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us00/_0936_ ( .A1(\us00\/_0050_ ), .A2(\us00\/_0118_ ), .B1(\us00\/_0194_ ), .Y(\us00\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us00/_0937_ ( .A(\us00\/_0113_ ), .Y(\us00\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us00/_0938_ ( .A1(\us00\/_0116_ ), .A2(\us00\/_0117_ ), .A3(\us00\/_0119_ ), .B1(\us00\/_0120_ ), .X(\us00\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us00/_0939_ ( .A(\us00\/_0104_ ), .B(\us00\/_0108_ ), .C(\us00\/_0115_ ), .D(\us00\/_0121_ ), .X(\us00\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_0940_ ( .A(\sa00\[7\] ), .B(\sa00\[6\] ), .Y(\us00\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0941_ ( .A(\us00\/_0749_ ), .B(\us00\/_0123_ ), .X(\us00\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0943_ ( .A(\us00\/_0082_ ), .B(\us00\/_0124_ ), .X(\us00\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_0944_ ( .A(\us00\/_0271_ ), .B(\us00\/_0124_ ), .Y(\us00\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0945_ ( .A(\us00\/_0124_ ), .X(\us00\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0946_ ( .A(\us00\/_0260_ ), .B(\us00\/_0325_ ), .X(\us00\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_0948_ ( .A(\us00\/_0128_ ), .B(\us00\/_0130_ ), .Y(\us00\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_0949_ ( .A(\us00\/_0127_ ), .B(\us00\/_0132_ ), .Y(\us00\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us00/_0950_ ( .A(\us00\/_0434_ ), .X(\us00\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_0951_ ( .A(\us00\/_0134_ ), .B(\us00\/_0128_ ), .Y(\us00\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us00/_0952_ ( .A(\us00\/_0126_ ), .B(\us00\/_0133_ ), .C_N(\us00\/_0135_ ), .Y(\us00\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0953_ ( .A(\us00\/_0026_ ), .B(\us00\/_0123_ ), .X(\us00\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0955_ ( .A(\us00\/_0137_ ), .X(\us00\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_0956_ ( .A1(\us00\/_0110_ ), .A2(\us00\/_0293_ ), .A3(\us00\/_0084_ ), .B1(\us00\/_0139_ ), .Y(\us00\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0957_ ( .A(\us00\/_0096_ ), .B(\us00\/_0730_ ), .X(\us00\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0959_ ( .A(\us00\/_0142_ ), .X(\us00\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_0960_ ( .A1(\us00\/_0020_ ), .A2(\us00\/_0144_ ), .A3(\us00\/_0017_ ), .B1(\us00\/_0139_ ), .Y(\us00\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \us00/_0961_ ( .A(\sa00\[2\] ), .B(\us00\/_0050_ ), .C_N(\sa00\[3\] ), .Y(\us00\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0962_ ( .A(\us00\/_0128_ ), .X(\us00\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_0963_ ( .A1(\us00\/_0146_ ), .A2(\us00\/_0032_ ), .A3(\us00\/_0640_ ), .B1(\us00\/_0147_ ), .Y(\us00\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us00/_0964_ ( .A(\us00\/_0136_ ), .B(\us00\/_0141_ ), .C(\us00\/_0145_ ), .D(\us00\/_0148_ ), .X(\us00\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0965_ ( .A(\us00\/_0123_ ), .B(\us00\/_0151_ ), .X(\us00\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0967_ ( .A(\us00\/_0150_ ), .X(\us00\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0968_ ( .A(\us00\/_0150_ ), .B(\us00\/_0062_ ), .X(\us00\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_0969_ ( .A(\us00\/_0079_ ), .B(\us00\/_0150_ ), .Y(\us00\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us00/_0970_ ( .A(\us00\/_0150_ ), .B(\us00\/_0412_ ), .C(\us00\/_0249_ ), .Y(\us00\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_0971_ ( .A(\us00\/_0155_ ), .B(\us00\/_0156_ ), .Y(\us00\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_0972_ ( .A1(\us00\/_0153_ ), .A2(\us00\/_0134_ ), .B1(\us00\/_0154_ ), .C1(\us00\/_0157_ ), .Y(\us00\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0973_ ( .A(\us00\/_0467_ ), .B(\us00\/_0123_ ), .X(\us00\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_0975_ ( .A(\us00\/_0159_ ), .X(\us00\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us00/_0976_ ( .A_N(\us00\/_0119_ ), .B(\us00\/_0161_ ), .X(\us00\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us00/_0977_ ( .A(\us00\/_0163_ ), .Y(\us00\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_0978_ ( .A1(\us00\/_0146_ ), .A2(\us00\/_0575_ ), .A3(\us00\/_0608_ ), .B1(\us00\/_0153_ ), .Y(\us00\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_0979_ ( .A1(\us00\/_0062_ ), .A2(\us00\/_0084_ ), .A3(\us00\/_0134_ ), .B1(\us00\/_0161_ ), .Y(\us00\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us00/_0980_ ( .A(\us00\/_0158_ ), .B(\us00\/_0164_ ), .C(\us00\/_0165_ ), .D(\us00\/_0166_ ), .X(\us00\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us00/_0981_ ( .A(\us00\/_0097_ ), .B(\us00\/_0122_ ), .C(\us00\/_0149_ ), .D(\us00\/_0167_ ), .X(\us00\/_0168_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0982_ ( .A(\us00\/_0662_ ), .B(\us00\/_0150_ ), .X(\us00\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_0983_ ( .A(\us00\/_0154_ ), .B(\us00\/_0169_ ), .Y(\us00\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us00/_0984_ ( .A(\us00\/_0123_ ), .B(\us00\/_0151_ ), .C(\us00\/_0038_ ), .X(\us00\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0985_ ( .A(\us00\/_0170_ ), .B(\us00\/_0171_ ), .X(\us00\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \us00/_0986_ ( .A(\us00\/_0172_ ), .Y(\us00\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \us00/_0987_ ( .A(\us00\/_0067_ ), .B(\us00\/_0168_ ), .C(\us00\/_0174_ ), .Y(\us00\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us00/_0988_ ( .A(\sa00\[1\] ), .B(\sa00\[0\] ), .Y(\us00\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us00/_0989_ ( .A(\us00\/_0175_ ), .B(\us00\/_0358_ ), .X(\us00\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0990_ ( .A(\us00\/_0176_ ), .B(\us00\/_0478_ ), .X(\us00\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_0991_ ( .A(\us00\/_0084_ ), .B(\us00\/_0113_ ), .Y(\us00\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0992_ ( .A(\us00\/_0111_ ), .B(\us00\/_0062_ ), .X(\us00\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0993_ ( .A(\us00\/_0111_ ), .B(\us00\/_0662_ ), .X(\us00\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_0994_ ( .A(\us00\/_0179_ ), .B(\us00\/_0180_ ), .Y(\us00\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0995_ ( .A(\us00\/_0054_ ), .B(\us00\/_0058_ ), .X(\us00\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us00/_0996_ ( .A(\us00\/_0182_ ), .Y(\us00\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us00/_0997_ ( .A_N(\us00\/_0177_ ), .B(\us00\/_0178_ ), .C(\us00\/_0181_ ), .D(\us00\/_0184_ ), .X(\us00\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0998_ ( .A(\us00\/_0098_ ), .B(\us00\/_0741_ ), .X(\us00\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us00/_0999_ ( .A(\us00\/_0047_ ), .B(\us00\/_0098_ ), .X(\us00\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us00/_1000_ ( .A(\us00\/_0186_ ), .B(\us00\/_0187_ ), .X(\us00\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1001_ ( .A(\us00\/_0188_ ), .Y(\us00\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1002_ ( .A(\us00\/_0738_ ), .B(\us00\/_0735_ ), .X(\us00\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1003_ ( .A(\us00\/_0271_ ), .B(\us00\/_0736_ ), .X(\us00\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_1004_ ( .A(\us00\/_0190_ ), .B(\us00\/_0191_ ), .Y(\us00\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us00/_1005_ ( .A(\us00\/_0096_ ), .B(\us00\/_0325_ ), .X(\us00\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1006_ ( .A1(\us00\/_0193_ ), .A2(\us00\/_0176_ ), .B1(\us00\/_0043_ ), .Y(\us00\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1007_ ( .A(\us00\/_0185_ ), .B(\us00\/_0189_ ), .C(\us00\/_0192_ ), .D(\us00\/_0195_ ), .X(\us00\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us00/_1008_ ( .A_N(\sa00\[3\] ), .B(\us00\/_0734_ ), .C(\sa00\[2\] ), .X(\us00\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1009_ ( .A(\us00\/_0137_ ), .B(\us00\/_0197_ ), .X(\us00\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_1010_ ( .A(\us00\/_0198_ ), .B(\us00\/_0040_ ), .Y(\us00\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1011_ ( .A(\us00\/_0293_ ), .B(\us00\/_0137_ ), .X(\us00\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1012_ ( .A(\us00\/_0200_ ), .Y(\us00\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1013_ ( .A(\us00\/_0137_ ), .B(\us00\/_0110_ ), .Y(\us00\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1014_ ( .A(\us00\/_0139_ ), .B(\us00\/_0020_ ), .Y(\us00\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1015_ ( .A(\us00\/_0199_ ), .B(\us00\/_0201_ ), .C(\us00\/_0202_ ), .D(\us00\/_0203_ ), .X(\us00\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us00/_1016_ ( .A1(\us00\/_0532_ ), .A2(\us00\/_0109_ ), .B1(\us00\/_0102_ ), .C1(\us00\/_0727_ ), .X(\us00\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1017_ ( .A(\us00\/_0022_ ), .B(\us00\/_0078_ ), .Y(\us00\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1018_ ( .A(\us00\/_0078_ ), .B(\us00\/_0142_ ), .Y(\us00\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1019_ ( .A(\us00\/_0207_ ), .B(\us00\/_0208_ ), .Y(\us00\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1020_ ( .A1(\us00\/_0094_ ), .A2(\us00\/_0176_ ), .B1(\us00\/_0206_ ), .C1(\us00\/_0209_ ), .Y(\us00\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1021_ ( .A(\us00\/_0662_ ), .B(\us00\/_0070_ ), .X(\us00\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us00/_1022_ ( .A(\us00\/_0732_ ), .B(\us00\/_0123_ ), .C(\us00\/_0749_ ), .Y(\us00\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us00/_1023_ ( .A(\us00\/_0732_ ), .B(\us00\/_0467_ ), .C(\us00\/_0069_ ), .Y(\us00\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us00/_1024_ ( .A_N(\us00\/_0211_ ), .B(\us00\/_0127_ ), .C(\us00\/_0212_ ), .D(\us00\/_0213_ ), .X(\us00\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1025_ ( .A(\us00\/_0137_ ), .Y(\us00\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1026_ ( .A(\us00\/_0128_ ), .B(\us00\/_0035_ ), .Y(\us00\/_0217_ ) );
sky130_fd_sc_hd__buf_2 \us00/_1027_ ( .A(\us00\/_0478_ ), .X(\us00\/_0218_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1028_ ( .A1(\us00\/_0159_ ), .A2(\us00\/_0747_ ), .B1(\us00\/_0434_ ), .B2(\us00\/_0218_ ), .Y(\us00\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us00/_1029_ ( .A1(\us00\/_0116_ ), .A2(\us00\/_0215_ ), .B1(\us00\/_0217_ ), .C1(\us00\/_0219_ ), .X(\us00\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1030_ ( .A(\us00\/_0113_ ), .B(\us00\/_0746_ ), .X(\us00\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us00/_1031_ ( .A1(\us00\/_0098_ ), .A2(\us00\/_0746_ ), .B1(\us00\/_0434_ ), .B2(\us00\/_0750_ ), .X(\us00\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1032_ ( .A1(\us00\/_0047_ ), .A2(\us00\/_0113_ ), .B1(\us00\/_0221_ ), .C1(\us00\/_0222_ ), .Y(\us00\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us00/_1033_ ( .A1(\us00\/_0129_ ), .A2(\us00\/_0162_ ), .B1(\us00\/_0271_ ), .B2(\us00\/_0705_ ), .X(\us00\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1034_ ( .A1(\us00\/_0093_ ), .A2(\us00\/_0738_ ), .B1(\us00\/_0081_ ), .C1(\us00\/_0224_ ), .Y(\us00\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1035_ ( .A(\us00\/_0214_ ), .B(\us00\/_0220_ ), .C(\us00\/_0223_ ), .D(\us00\/_0225_ ), .X(\us00\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1036_ ( .A(\us00\/_0196_ ), .B(\us00\/_0204_ ), .C(\us00\/_0210_ ), .D(\us00\/_0226_ ), .X(\us00\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1037_ ( .A(\us00\/_0111_ ), .B(\us00\/_0554_ ), .X(\us00\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1038_ ( .A(\us00\/_0229_ ), .Y(\us00\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1039_ ( .A(\us00\/_0111_ ), .B(\us00\/_0129_ ), .Y(\us00\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1040_ ( .A(\us00\/_0017_ ), .B(\us00\/_0738_ ), .Y(\us00\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1041_ ( .A(\us00\/_0030_ ), .B(\us00\/_0304_ ), .Y(\us00\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1042_ ( .A(\us00\/_0230_ ), .B(\us00\/_0231_ ), .C(\us00\/_0232_ ), .D(\us00\/_0233_ ), .X(\us00\/_0234_ ) );
sky130_fd_sc_hd__and2_1 \us00/_1043_ ( .A(\us00\/_0047_ ), .B(\us00\/_0478_ ), .X(\us00\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1044_ ( .A1(\us00\/_0129_ ), .A2(\us00\/_0554_ ), .B1(\us00\/_0137_ ), .Y(\us00\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us00/_1045_ ( .A(\us00\/_0235_ ), .B(\us00\/_0049_ ), .C_N(\us00\/_0236_ ), .Y(\us00\/_0237_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1046_ ( .A(\us00\/_0047_ ), .B(\us00\/_0077_ ), .X(\us00\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1047_ ( .A(\us00\/_0070_ ), .B(\us00\/_0035_ ), .X(\us00\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us00/_1048_ ( .A1(\us00\/_0047_ ), .A2(\us00\/_0736_ ), .B1(\us00\/_0022_ ), .B2(\us00\/_0099_ ), .X(\us00\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us00/_1049_ ( .A(\us00\/_0239_ ), .B(\us00\/_0240_ ), .C(\us00\/_0241_ ), .Y(\us00\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1050_ ( .A(\us00\/_0554_ ), .B(\us00\/_0072_ ), .X(\us00\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us00/_1051_ ( .A1(\us00\/_0142_ ), .A2(\us00\/_0137_ ), .B1(\us00\/_0159_ ), .B2(\us00\/_0082_ ), .X(\us00\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1052_ ( .A1(\us00\/_0608_ ), .A2(\us00\/_0072_ ), .B1(\us00\/_0243_ ), .C1(\us00\/_0244_ ), .Y(\us00\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1053_ ( .A(\us00\/_0234_ ), .B(\us00\/_0237_ ), .C(\us00\/_0242_ ), .D(\us00\/_0245_ ), .X(\us00\/_0246_ ) );
sky130_fd_sc_hd__buf_2 \us00/_1054_ ( .A(\us00\/_0027_ ), .X(\us00\/_0247_ ) );
sky130_fd_sc_hd__o21a_1 \us00/_1055_ ( .A1(\us00\/_0554_ ), .A2(\us00\/_0586_ ), .B1(\us00\/_0247_ ), .X(\us00\/_0248_ ) );
sky130_fd_sc_hd__and2_1 \us00/_1056_ ( .A(\us00\/_0082_ ), .B(\us00\/_0478_ ), .X(\us00\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_1057_ ( .A(\us00\/_0079_ ), .X(\us00\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1058_ ( .A(\us00\/_0251_ ), .B(\us00\/_0478_ ), .X(\us00\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_1059_ ( .A(\us00\/_0250_ ), .B(\us00\/_0252_ ), .Y(\us00\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1060_ ( .A(\us00\/_0016_ ), .B(\us00\/_0064_ ), .Y(\us00\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_1061_ ( .A(\us00\/_0304_ ), .X(\us00\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1062_ ( .A(\us00\/_0255_ ), .B(\us00\/_0640_ ), .Y(\us00\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us00/_1063_ ( .A_N(\us00\/_0248_ ), .B(\us00\/_0253_ ), .C(\us00\/_0254_ ), .D(\us00\/_0256_ ), .X(\us00\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1064_ ( .A(\us00\/_0099_ ), .B(\us00\/_0110_ ), .X(\us00\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us00/_1065_ ( .A1(\us00\/_0161_ ), .A2(\us00\/_0130_ ), .B1(\us00\/_0258_ ), .Y(\us00\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1066_ ( .A(\us00\/_0194_ ), .B(\sa00\[1\] ), .X(\us00\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1068_ ( .A(\us00\/_0261_ ), .B(\us00\/_0153_ ), .Y(\us00\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us00/_1069_ ( .A_N(\us00\/_0154_ ), .B(\us00\/_0259_ ), .C(\us00\/_0263_ ), .X(\us00\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1070_ ( .A(\us00\/_0246_ ), .B(\us00\/_0174_ ), .C(\us00\/_0257_ ), .D(\us00\/_0264_ ), .X(\us00\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us00/_1071_ ( .A1(\us00\/_0261_ ), .A2(\us00\/_0554_ ), .B1(\us00\/_0159_ ), .X(\us00\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1072_ ( .A(\us00\/_0747_ ), .B(\us00\/_0150_ ), .Y(\us00\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1073_ ( .A(\us00\/_0175_ ), .Y(\us00\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us00/_1074_ ( .A(\us00\/_0412_ ), .B(\us00\/_0123_ ), .C(\us00\/_0151_ ), .X(\us00\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1075_ ( .A(\us00\/_0268_ ), .B(\us00\/_0269_ ), .Y(\us00\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us00/_1076_ ( .A_N(\us00\/_0266_ ), .B(\us00\/_0267_ ), .C(\us00\/_0270_ ), .X(\us00\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1077_ ( .A(\us00\/_0554_ ), .B(\us00\/_0150_ ), .X(\us00\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1078_ ( .A(\us00\/_0273_ ), .Y(\us00\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1079_ ( .A1(\us00\/_0734_ ), .A2(\us00\/_0325_ ), .B1(\us00\/_0380_ ), .Y(\us00\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1080_ ( .A(\us00\/_0275_ ), .Y(\us00\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1081_ ( .A(\us00\/_0276_ ), .B(\us00\/_0153_ ), .Y(\us00\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us00/_1082_ ( .A(\us00\/_0272_ ), .B(\us00\/_0274_ ), .C(\us00\/_0277_ ), .X(\us00\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_1083_ ( .A(\us00\/_0035_ ), .X(\us00\/_0279_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1085_ ( .A1(\us00\/_0218_ ), .A2(\us00\/_0279_ ), .B1(\us00\/_0084_ ), .B2(\us00\/_0060_ ), .Y(\us00\/_0281_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1086_ ( .A1(\us00\/_0251_ ), .A2(\us00\/_0434_ ), .B1(\us00\/_0304_ ), .Y(\us00\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1087_ ( .A(\us00\/_0091_ ), .B(\us00\/_0292_ ), .Y(\us00\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1088_ ( .A1(\us00\/_0118_ ), .A2(\us00\/_0050_ ), .B1(\us00\/_0038_ ), .C1(\us00\/_0255_ ), .Y(\us00\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1089_ ( .A(\us00\/_0281_ ), .B(\us00\/_0283_ ), .C(\us00\/_0284_ ), .D(\us00\/_0285_ ), .X(\us00\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1090_ ( .A(\us00\/_0082_ ), .B(\us00\/_0027_ ), .X(\us00\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1091_ ( .A(\us00\/_0129_ ), .B(\us00\/_0027_ ), .X(\us00\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_1092_ ( .A(\us00\/_0287_ ), .B(\us00\/_0288_ ), .Y(\us00\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1093_ ( .A1(\us00\/_0752_ ), .A2(\us00\/_0683_ ), .B1(\us00\/_0093_ ), .B2(\us00\/_0247_ ), .Y(\us00\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1094_ ( .A1(\us00\/_0092_ ), .A2(\us00\/_0575_ ), .B1(\us00\/_0292_ ), .Y(\us00\/_0291_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_1095_ ( .A(\us00\/_0054_ ), .X(\us00\/_0292_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1096_ ( .A1(\us00\/_0218_ ), .A2(\us00\/_0662_ ), .B1(\us00\/_0084_ ), .B2(\us00\/_0292_ ), .Y(\us00\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1097_ ( .A(\us00\/_0289_ ), .B(\us00\/_0290_ ), .C(\us00\/_0291_ ), .D(\us00\/_0294_ ), .X(\us00\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1098_ ( .A(\us00\/_0750_ ), .B(\us00\/_0193_ ), .X(\us00\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1099_ ( .A(\us00\/_0705_ ), .B(\us00\/_0380_ ), .X(\us00\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1100_ ( .A(\us00\/_0752_ ), .B(\us00\/_0129_ ), .Y(\us00\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us00/_1101_ ( .A(\us00\/_0296_ ), .B(\us00\/_0297_ ), .C_N(\us00\/_0298_ ), .Y(\us00\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1102_ ( .A(\us00\/_0089_ ), .B(\us00\/_0532_ ), .Y(\us00\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1103_ ( .A(\sa00\[2\] ), .Y(\us00\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \us00/_1104_ ( .A(\us00\/_0301_ ), .B(\sa00\[3\] ), .C(\us00\/_0118_ ), .Y(\us00\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1105_ ( .A(\us00\/_0072_ ), .B(\us00\/_0302_ ), .X(\us00\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1106_ ( .A(\us00\/_0303_ ), .Y(\us00\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1107_ ( .A(\us00\/_0147_ ), .B(\us00\/_0302_ ), .Y(\us00\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1108_ ( .A(\us00\/_0299_ ), .B(\us00\/_0300_ ), .C(\us00\/_0305_ ), .D(\us00\/_0306_ ), .X(\us00\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1109_ ( .A(\us00\/_0278_ ), .B(\us00\/_0286_ ), .C(\us00\/_0295_ ), .D(\us00\/_0307_ ), .X(\us00\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us00/_1110_ ( .A(\us00\/_0228_ ), .B(\us00\/_0265_ ), .C(\us00\/_0308_ ), .Y(\us00\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1111_ ( .A(\us00\/_0235_ ), .Y(\us00\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1112_ ( .A(\us00\/_0478_ ), .B(\us00\/_0640_ ), .X(\us00\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1113_ ( .A(\us00\/_0310_ ), .Y(\us00\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1114_ ( .A(\us00\/_0022_ ), .B(\us00\/_0218_ ), .Y(\us00\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1115_ ( .A(\us00\/_0218_ ), .B(\us00\/_0032_ ), .Y(\us00\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1116_ ( .A(\us00\/_0309_ ), .B(\us00\/_0311_ ), .C(\us00\/_0312_ ), .D(\us00\/_0313_ ), .X(\us00\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1117_ ( .A(\us00\/_0218_ ), .B(\us00\/_0064_ ), .Y(\us00\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1118_ ( .A(\us00\/_0218_ ), .B(\us00\/_0683_ ), .Y(\us00\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1119_ ( .A(\us00\/_0315_ ), .B(\us00\/_0316_ ), .C(\us00\/_0317_ ), .D(\us00\/_0253_ ), .X(\us00\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1120_ ( .A(\us00\/_0047_ ), .B(\us00\/_0304_ ), .Y(\us00\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1121_ ( .A(\us00\/_0586_ ), .B(\us00\/_0162_ ), .Y(\us00\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1122_ ( .A(\us00\/_0319_ ), .B(\us00\/_0320_ ), .Y(\us00\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_1123_ ( .A(\us00\/_0321_ ), .B(\us00\/_0238_ ), .Y(\us00\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1124_ ( .A(\us00\/_0304_ ), .B(\us00\/_0062_ ), .Y(\us00\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_1125_ ( .A(\us00\/_0251_ ), .X(\us00\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1126_ ( .A1(\us00\/_0324_ ), .A2(\us00\/_0084_ ), .B1(\us00\/_0255_ ), .Y(\us00\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1127_ ( .A1(\us00\/_0050_ ), .A2(\us00\/_0205_ ), .B1(\us00\/_0109_ ), .C1(\us00\/_0255_ ), .Y(\us00\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1128_ ( .A(\us00\/_0322_ ), .B(\us00\/_0323_ ), .C(\us00\/_0326_ ), .D(\us00\/_0327_ ), .X(\us00\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1129_ ( .A1(\us00\/_0733_ ), .A2(\us00\/_0279_ ), .A3(\us00\/_0058_ ), .B1(\us00\/_0292_ ), .Y(\us00\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_1130_ ( .A(\us00\/_0047_ ), .X(\us00\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1131_ ( .A(\us00\/_0330_ ), .B(\us00\/_0292_ ), .Y(\us00\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1132_ ( .A(\us00\/_0054_ ), .B(\us00\/_0045_ ), .Y(\us00\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1133_ ( .A(\us00\/_0329_ ), .B(\us00\/_0331_ ), .C(\us00\/_0284_ ), .D(\us00\/_0332_ ), .X(\us00\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us00/_1134_ ( .A1(\us00\/_0249_ ), .A2(\us00\/_0205_ ), .B1(\us00\/_0532_ ), .C1(\us00\/_0060_ ), .X(\us00\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1135_ ( .A(\us00\/_0084_ ), .B(\us00\/_0060_ ), .Y(\us00\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1136_ ( .A(\us00\/_0324_ ), .B(\us00\/_0060_ ), .Y(\us00\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1137_ ( .A(\us00\/_0335_ ), .B(\us00\/_0337_ ), .Y(\us00\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1138_ ( .A1(\us00\/_0276_ ), .A2(\us00\/_0060_ ), .B1(\us00\/_0334_ ), .C1(\us00\/_0338_ ), .Y(\us00\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1139_ ( .A(\us00\/_0318_ ), .B(\us00\/_0328_ ), .C(\us00\/_0333_ ), .D(\us00\/_0339_ ), .X(\us00\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us00/_1140_ ( .A1(\us00\/_0747_ ), .A2(\us00\/_0134_ ), .B1(\us00\/_0128_ ), .X(\us00\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us00/_1141_ ( .A_N(\us00\/_0086_ ), .B(\us00\/_0128_ ), .X(\us00\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1142_ ( .A(\us00\/_0079_ ), .B(\us00\/_0124_ ), .X(\us00\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_1143_ ( .A(\us00\/_0126_ ), .B(\us00\/_0343_ ), .Y(\us00\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us00/_1144_ ( .A(\us00\/_0341_ ), .B(\us00\/_0342_ ), .C_N(\us00\/_0344_ ), .Y(\us00\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1146_ ( .A1(\us00\/_0193_ ), .A2(\us00\/_0092_ ), .A3(\us00\/_0330_ ), .B1(\us00\/_0147_ ), .Y(\us00\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1147_ ( .A1(\us00\/_0130_ ), .A2(\us00\/_0084_ ), .A3(\us00\/_0134_ ), .B1(\us00\/_0139_ ), .Y(\us00\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1148_ ( .A1(\us00\/_0144_ ), .A2(\us00\/_0608_ ), .A3(\us00\/_0092_ ), .B1(\us00\/_0139_ ), .Y(\us00\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1149_ ( .A(\us00\/_0345_ ), .B(\us00\/_0348_ ), .C(\us00\/_0349_ ), .D(\us00\/_0350_ ), .X(\us00\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us00/_1150_ ( .A(\us00\/_0150_ ), .B(\us00\/_0194_ ), .C(\us00\/_0249_ ), .X(\us00\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us00/_1151_ ( .A(\us00\/_0277_ ), .SLEEP(\us00\/_0352_ ), .X(\us00\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us00/_1152_ ( .A1(\us00\/_0268_ ), .A2(\us00\/_0171_ ), .B1(\us00\/_0157_ ), .Y(\us00\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us00/_1153_ ( .A(\us00\/_0161_ ), .X(\us00\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1154_ ( .A1(\us00\/_0279_ ), .A2(\us00\/_0084_ ), .B1(\us00\/_0355_ ), .Y(\us00\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1155_ ( .A1(\us00\/_0020_ ), .A2(\us00\/_0193_ ), .A3(\us00\/_0091_ ), .B1(\us00\/_0355_ ), .Y(\us00\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1156_ ( .A(\us00\/_0353_ ), .B(\us00\/_0354_ ), .C(\us00\/_0356_ ), .D(\us00\/_0357_ ), .X(\us00\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1157_ ( .A(\us00\/_0111_ ), .B(\us00\/_0586_ ), .X(\us00\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1158_ ( .A(\us00\/_0360_ ), .Y(\us00\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us00/_1159_ ( .A1(\us00\/_0119_ ), .A2(\us00\/_0120_ ), .B1(\us00\/_0230_ ), .C1(\us00\/_0361_ ), .X(\us00\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1160_ ( .A1(\us00\/_0662_ ), .A2(\us00\/_0251_ ), .A3(\us00\/_0134_ ), .B1(\us00\/_0114_ ), .Y(\us00\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1162_ ( .A1(\us00\/_0035_ ), .A2(\us00\/_0251_ ), .A3(\us00\/_0134_ ), .B1(\us00\/_0099_ ), .Y(\us00\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1163_ ( .A1(\us00\/_0193_ ), .A2(\us00\/_0608_ ), .B1(\us00\/_0099_ ), .Y(\us00\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1164_ ( .A(\us00\/_0362_ ), .B(\us00\/_0363_ ), .C(\us00\/_0365_ ), .D(\us00\/_0366_ ), .X(\us00\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1165_ ( .A1(\us00\/_0575_ ), .A2(\us00\/_0092_ ), .A3(\us00\/_0330_ ), .B1(\us00\/_0089_ ), .Y(\us00\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1166_ ( .A1(\us00\/_0586_ ), .A2(\us00\/_0017_ ), .A3(\us00\/_0330_ ), .B1(\us00\/_0094_ ), .Y(\us00\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \us00/_1167_ ( .A1(\us00\/_0293_ ), .A2(\us00\/_0134_ ), .B1(\us00\/_0089_ ), .Y(\us00\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1168_ ( .A1(\us00\/_0279_ ), .A2(\us00\/_0134_ ), .B1(\us00\/_0094_ ), .Y(\us00\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1169_ ( .A(\us00\/_0368_ ), .B(\us00\/_0370_ ), .C(\us00\/_0371_ ), .D(\us00\/_0372_ ), .X(\us00\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1170_ ( .A(\us00\/_0351_ ), .B(\us00\/_0359_ ), .C(\us00\/_0367_ ), .D(\us00\/_0373_ ), .X(\us00\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1171_ ( .A1(\us00\/_0102_ ), .A2(\us00\/_0347_ ), .B1(\us00\/_0109_ ), .C1(\us00\/_0247_ ), .Y(\us00\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1172_ ( .A1(\us00\/_0102_ ), .A2(\us00\/_0347_ ), .B1(\us00\/_0532_ ), .C1(\us00\/_0247_ ), .Y(\us00\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1173_ ( .A1(\us00\/_0050_ ), .A2(\us00\/_0249_ ), .B1(\us00\/_0380_ ), .C1(\us00\/_0247_ ), .Y(\us00\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1174_ ( .A(\us00\/_0041_ ), .B(\us00\/_0375_ ), .C(\us00\/_0376_ ), .D(\us00\/_0377_ ), .X(\us00\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1175_ ( .A(\us00\/_0047_ ), .B(\us00\/_0750_ ), .X(\us00\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1176_ ( .A(\us00\/_0379_ ), .Y(\us00\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1177_ ( .A(\us00\/_0016_ ), .B(\us00\/_0608_ ), .Y(\us00\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1178_ ( .A(\us00\/_0752_ ), .B(\us00\/_0554_ ), .Y(\us00\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1179_ ( .A1(\sa00\[1\] ), .A2(\us00\/_0734_ ), .B1(\us00\/_0109_ ), .C1(\us00\/_0016_ ), .Y(\us00\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1180_ ( .A(\us00\/_0381_ ), .B(\us00\/_0382_ ), .C(\us00\/_0383_ ), .D(\us00\/_0384_ ), .X(\us00\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us00/_1181_ ( .A(\us00\/_0086_ ), .B_N(\us00\/_0736_ ), .X(\us00\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1182_ ( .A1(\us00\/_0748_ ), .A2(\us00\/_0134_ ), .B1(\us00\/_0739_ ), .Y(\us00\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1183_ ( .A1(\us00\/_0118_ ), .A2(\us00\/_0249_ ), .B1(\us00\/_0109_ ), .C1(\us00\/_0739_ ), .Y(\us00\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1184_ ( .A1(\us00\/_0102_ ), .A2(\us00\/_0301_ ), .B1(\sa00\[3\] ), .C1(\us00\/_0739_ ), .Y(\us00\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1185_ ( .A(\us00\/_0386_ ), .B(\us00\/_0387_ ), .C(\us00\/_0388_ ), .D(\us00\/_0389_ ), .X(\us00\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1186_ ( .A(\us00\/_0020_ ), .Y(\us00\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1187_ ( .A(\us00\/_0727_ ), .Y(\us00\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1188_ ( .A(\us00\/_0727_ ), .B(\us00\/_0064_ ), .Y(\us00\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1189_ ( .A1(\us00\/_0102_ ), .A2(\us00\/_0734_ ), .B1(\us00\/_0532_ ), .C1(\us00\/_0727_ ), .Y(\us00\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us00/_1190_ ( .A1(\us00\/_0392_ ), .A2(\us00\/_0393_ ), .B1(\us00\/_0394_ ), .C1(\us00\/_0395_ ), .X(\us00\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1191_ ( .A(\us00\/_0378_ ), .B(\us00\/_0385_ ), .C(\us00\/_0390_ ), .D(\us00\/_0396_ ), .X(\us00\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us00/_1192_ ( .A(\us00\/_0340_ ), .B(\us00\/_0374_ ), .C(\us00\/_0397_ ), .Y(\us00\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1193_ ( .A(\us00\/_0077_ ), .B(\us00\/_0129_ ), .X(\us00\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_1194_ ( .A(\us00\/_0398_ ), .B(\us00\/_0239_ ), .Y(\us00\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1195_ ( .A(\us00\/_0022_ ), .B(\us00\/_0111_ ), .X(\us00\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us00/_1196_ ( .A_N(\us00\/_0400_ ), .B(\us00\/_0231_ ), .Y(\us00\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us00/_1197_ ( .A(\us00\/_0399_ ), .SLEEP(\us00\/_0402_ ), .X(\us00\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_1198_ ( .A(\us00\/_0747_ ), .B(\us00\/_0251_ ), .Y(\us00\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us00/_1199_ ( .A_N(\us00\/_0404_ ), .B(\us00\/_0752_ ), .Y(\us00\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us00/_1200_ ( .A(\us00\/_0467_ ), .B(\us00\/_0194_ ), .C(\us00\/_0694_ ), .X(\us00\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us00/_1201_ ( .A_N(\us00\/_0175_ ), .B(\us00\/_0406_ ), .X(\us00\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1202_ ( .A(\us00\/_0407_ ), .Y(\us00\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1203_ ( .A1(\us00\/_0094_ ), .A2(\us00\/_0197_ ), .B1(\us00\/_0114_ ), .B2(\us00\/_0640_ ), .Y(\us00\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1204_ ( .A(\us00\/_0403_ ), .B(\us00\/_0405_ ), .C(\us00\/_0408_ ), .D(\us00\/_0409_ ), .X(\us00\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1205_ ( .A(\us00\/_0030_ ), .B(\us00\/_0150_ ), .Y(\us00\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us00/_1206_ ( .A_N(\us00\/_0169_ ), .B(\us00\/_0289_ ), .C(\us00\/_0411_ ), .X(\us00\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us00/_1207_ ( .A1(\us00\/_0467_ ), .A2(\us00\/_0151_ ), .B1(\us00\/_0140_ ), .C1(\us00\/_0129_ ), .X(\us00\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1208_ ( .A1(\us00\/_0608_ ), .A2(\us00\/_0099_ ), .B1(\us00\/_0037_ ), .C1(\us00\/_0414_ ), .Y(\us00\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1209_ ( .A(\us00\/_0738_ ), .Y(\us00\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1210_ ( .A(\us00\/_0586_ ), .B(\us00\/_0736_ ), .Y(\us00\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1211_ ( .A1(\us00\/_0194_ ), .A2(\us00\/_0038_ ), .B1(\us00\/_0118_ ), .C1(\us00\/_0153_ ), .Y(\us00\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us00/_1212_ ( .A1(\us00\/_0416_ ), .A2(\us00\/_0117_ ), .B1(\us00\/_0417_ ), .C1(\us00\/_0418_ ), .X(\us00\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1213_ ( .A(\us00\/_0077_ ), .B(\us00\/_0035_ ), .X(\us00\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1214_ ( .A(\us00\/_0662_ ), .B(\us00\/_0124_ ), .Y(\us00\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1215_ ( .A(\us00\/_0030_ ), .B(\us00\/_0137_ ), .Y(\us00\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1216_ ( .A(\us00\/_0072_ ), .B(\us00\/_0732_ ), .Y(\us00\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us00/_1217_ ( .A_N(\us00\/_0420_ ), .B(\us00\/_0421_ ), .C(\us00\/_0422_ ), .D(\us00\/_0424_ ), .X(\us00\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1218_ ( .A(\us00\/_0413_ ), .B(\us00\/_0415_ ), .C(\us00\/_0419_ ), .D(\us00\/_0425_ ), .X(\us00\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us00/_1219_ ( .A(\us00\/_0355_ ), .B(\us00\/_0102_ ), .C(\us00\/_0109_ ), .Y(\us00\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1220_ ( .A(\us00\/_0077_ ), .B(\us00\/_0017_ ), .X(\us00\/_0428_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1221_ ( .A(\us00\/_0077_ ), .B(\us00\/_0554_ ), .X(\us00\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us00/_1222_ ( .A1(\us00\/_0050_ ), .A2(\us00\/_0205_ ), .B1(\us00\/_0380_ ), .C1(\us00\/_0078_ ), .X(\us00\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us00/_1223_ ( .A(\us00\/_0428_ ), .B(\us00\/_0429_ ), .C(\us00\/_0430_ ), .Y(\us00\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us00/_1224_ ( .A_N(\us00\/_0209_ ), .B(\us00\/_0431_ ), .X(\us00\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us00/_1225_ ( .A1(\us00\/_0215_ ), .A2(\us00\/_0404_ ), .B1(\us00\/_0427_ ), .C1(\us00\/_0432_ ), .X(\us00\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1226_ ( .A(\us00\/_0043_ ), .B(\us00\/_0058_ ), .Y(\us00\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1227_ ( .A(\us00\/_0195_ ), .B(\us00\/_0233_ ), .C(\us00\/_0320_ ), .D(\us00\/_0435_ ), .X(\us00\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1228_ ( .A(\us00\/_0261_ ), .B(\us00\/_0738_ ), .Y(\us00\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1229_ ( .A1(\us00\/_0218_ ), .A2(\us00\/_0640_ ), .B1(\us00\/_0261_ ), .B2(\us00\/_0292_ ), .Y(\us00\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1230_ ( .A(\us00\/_0436_ ), .B(\us00\/_0394_ ), .C(\us00\/_0437_ ), .D(\us00\/_0438_ ), .X(\us00\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1231_ ( .A(\us00\/_0410_ ), .B(\us00\/_0426_ ), .C(\us00\/_0433_ ), .D(\us00\/_0439_ ), .X(\us00\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us00/_1232_ ( .A(\us00\/_0135_ ), .SLEEP(\us00\/_0273_ ), .X(\us00\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1233_ ( .A1(\us00\/_0279_ ), .A2(\us00\/_0134_ ), .B1(\us00\/_0099_ ), .Y(\us00\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1234_ ( .A(\us00\/_0441_ ), .B(\us00\/_0164_ ), .C(\us00\/_0270_ ), .D(\us00\/_0442_ ), .X(\us00\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1235_ ( .A(\us00\/_0051_ ), .B(\us00\/_0662_ ), .Y(\us00\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1236_ ( .A(\us00\/_0051_ ), .B(\us00\/_0271_ ), .Y(\us00\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1237_ ( .A(\us00\/_0444_ ), .B(\us00\/_0446_ ), .X(\us00\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1238_ ( .A(\us00\/_0193_ ), .B(\us00\/_0304_ ), .X(\us00\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1239_ ( .A(\us00\/_0448_ ), .Y(\us00\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1240_ ( .A(\us00\/_0162_ ), .B(\us00\/_0130_ ), .X(\us00\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1241_ ( .A(\us00\/_0450_ ), .Y(\us00\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1242_ ( .A1(\us00\/_0129_ ), .A2(\us00\/_0554_ ), .B1(\us00\/_0043_ ), .Y(\us00\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1243_ ( .A(\us00\/_0447_ ), .B(\us00\/_0449_ ), .C(\us00\/_0451_ ), .D(\us00\/_0452_ ), .X(\us00\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1244_ ( .A(\us00\/_0292_ ), .B(\us00\/_0064_ ), .Y(\us00\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us00/_1245_ ( .A_N(\us00\/_0248_ ), .B(\us00\/_0454_ ), .C(\us00\/_0254_ ), .D(\us00\/_0256_ ), .X(\us00\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1246_ ( .A1(\us00\/_0330_ ), .A2(\us00\/_0099_ ), .B1(\us00\/_0134_ ), .B2(\us00\/_0705_ ), .Y(\us00\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1247_ ( .A1(\us00\/_0748_ ), .A2(\us00\/_0738_ ), .B1(\us00\/_0092_ ), .B2(\us00\/_0752_ ), .Y(\us00\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1248_ ( .A1(\us00\/_0072_ ), .A2(\us00\/_0035_ ), .B1(\us00\/_0748_ ), .B2(\us00\/_0292_ ), .Y(\us00\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1249_ ( .A1(\us00\/_0748_ ), .A2(\us00\/_0251_ ), .B1(\us00\/_0247_ ), .Y(\us00\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1250_ ( .A(\us00\/_0457_ ), .B(\us00\/_0458_ ), .C(\us00\/_0459_ ), .D(\us00\/_0460_ ), .X(\us00\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1251_ ( .A(\us00\/_0443_ ), .B(\us00\/_0453_ ), .C(\us00\/_0455_ ), .D(\us00\/_0461_ ), .X(\us00\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1252_ ( .A(\us00\/_0705_ ), .B(\us00\/_0079_ ), .X(\us00\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1253_ ( .A(\us00\/_0586_ ), .B(\us00\/_0124_ ), .Y(\us00\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1254_ ( .A(\us00\/_0218_ ), .B(\us00\/_0747_ ), .Y(\us00\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us00/_1255_ ( .A_N(\us00\/_0463_ ), .B(\us00\/_0464_ ), .C(\us00\/_0465_ ), .X(\us00\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us00/_1256_ ( .A1(\us00\/_0271_ ), .A2(\us00\/_0072_ ), .B1(\us00\/_0142_ ), .B2(\us00\/_0027_ ), .X(\us00\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1257_ ( .A1(\us00\/_0144_ ), .A2(\us00\/_0099_ ), .B1(\us00\/_0360_ ), .C1(\us00\/_0468_ ), .Y(\us00\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us00/_1258_ ( .A1(\us00\/_0662_ ), .A2(\us00\/_0251_ ), .B1(\us00\/_0218_ ), .X(\us00\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1259_ ( .A1(\us00\/_0575_ ), .A2(\us00\/_0292_ ), .B1(\us00\/_0379_ ), .C1(\us00\/_0470_ ), .Y(\us00\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1260_ ( .A(\us00\/_0466_ ), .B(\us00\/_0469_ ), .C(\us00\/_0471_ ), .D(\us00\/_0305_ ), .X(\us00\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us00/_1261_ ( .A1(\us00\/_0247_ ), .A2(\us00\/_0683_ ), .B1(\us00\/_0324_ ), .B2(\us00\/_0292_ ), .X(\us00\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1262_ ( .A(\us00\/_0084_ ), .B(\us00\/_0099_ ), .X(\us00\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us00/_1263_ ( .A1(\us00\/_0092_ ), .A2(\us00\/_0247_ ), .B1(\us00\/_0474_ ), .X(\us00\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us00/_1264_ ( .A(\us00\/_0075_ ), .B(\us00\/_0473_ ), .C(\us00\/_0475_ ), .Y(\us00\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1265_ ( .A1(\us00\/_0279_ ), .A2(\us00\/_0255_ ), .B1(\us00\/_0084_ ), .B2(\us00\/_0060_ ), .Y(\us00\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1266_ ( .A1(\us00\/_0093_ ), .A2(\us00\/_0292_ ), .B1(\us00\/_0134_ ), .B2(\us00\/_0114_ ), .Y(\us00\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1267_ ( .A1(\us00\/_0161_ ), .A2(\us00\/_0032_ ), .B1(\us00\/_0324_ ), .B2(\us00\/_0147_ ), .Y(\us00\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1268_ ( .A1(\us00\/_0054_ ), .A2(\us00\/_0732_ ), .B1(\us00\/_0748_ ), .B2(\us00\/_0304_ ), .Y(\us00\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1269_ ( .A(\us00\/_0477_ ), .B(\us00\/_0479_ ), .C(\us00\/_0480_ ), .D(\us00\/_0481_ ), .X(\us00\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1270_ ( .A(\us00\/_0161_ ), .B(\us00\/_0064_ ), .Y(\us00\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us00/_1271_ ( .A(\us00\/_0732_ ), .B(\us00\/_0123_ ), .C(\us00\/_0467_ ), .Y(\us00\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1272_ ( .A(\us00\/_0483_ ), .B(\us00\/_0484_ ), .Y(\us00\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1273_ ( .A(\us00\/_0297_ ), .Y(\us00\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us00/_1274_ ( .A_N(\us00\/_0485_ ), .B(\us00\/_0181_ ), .C(\us00\/_0486_ ), .D(\us00\/_0386_ ), .X(\us00\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1275_ ( .A(\us00\/_0472_ ), .B(\us00\/_0476_ ), .C(\us00\/_0482_ ), .D(\us00\/_0487_ ), .X(\us00\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \us00/_1276_ ( .A(\us00\/_0440_ ), .B(\us00\/_0462_ ), .C(\us00\/_0488_ ), .Y(\us00\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1277_ ( .A(\us00\/_0403_ ), .B(\us00\/_0230_ ), .C(\us00\/_0451_ ), .D(\us00\/_0361_ ), .X(\us00\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1278_ ( .A1(\us00\/_0118_ ), .A2(\us00\/_0050_ ), .B1(\us00\/_0109_ ), .C1(\us00\/_0139_ ), .Y(\us00\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1279_ ( .A(\us00\/_0447_ ), .B(\us00\/_0437_ ), .C(\us00\/_0491_ ), .D(\us00\/_0427_ ), .X(\us00\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1280_ ( .A1(\us00\/_0084_ ), .A2(\us00\/_0255_ ), .B1(\us00\/_0608_ ), .B2(\us00\/_0247_ ), .Y(\us00\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1281_ ( .A1(\us00\/_0144_ ), .A2(\us00\/_0147_ ), .B1(\us00\/_0355_ ), .B2(\us00\/_0093_ ), .Y(\us00\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1282_ ( .A1(\us00\/_0705_ ), .A2(\us00\/_0279_ ), .B1(\us00\/_0330_ ), .B2(\us00\/_0247_ ), .Y(\us00\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1283_ ( .A1(\us00\/_0279_ ), .A2(\us00\/_0084_ ), .B1(\us00\/_0114_ ), .Y(\us00\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1284_ ( .A(\us00\/_0493_ ), .B(\us00\/_0494_ ), .C(\us00\/_0495_ ), .D(\us00\/_0496_ ), .X(\us00\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1285_ ( .A1(\us00\/_0134_ ), .A2(\us00\/_0137_ ), .B1(\us00\/_0355_ ), .B2(\us00\/_0575_ ), .Y(\us00\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1286_ ( .A1(\us00\/_0099_ ), .A2(\us00\/_0733_ ), .B1(\us00\/_0093_ ), .B2(\us00\/_0218_ ), .Y(\us00\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1287_ ( .A(\us00\/_0147_ ), .B(\us00\/_0640_ ), .Y(\us00\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1288_ ( .A1(\us00\/_0153_ ), .A2(\us00\/_0292_ ), .B1(\us00\/_0748_ ), .Y(\us00\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1289_ ( .A(\us00\/_0498_ ), .B(\us00\/_0500_ ), .C(\us00\/_0501_ ), .D(\us00\/_0502_ ), .X(\us00\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1290_ ( .A(\us00\/_0490_ ), .B(\us00\/_0492_ ), .C(\us00\/_0497_ ), .D(\us00\/_0503_ ), .X(\us00\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us00/_1291_ ( .A_N(\us00\/_0275_ ), .B(\us00\/_0705_ ), .X(\us00\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1292_ ( .A(\us00\/_0505_ ), .Y(\us00\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1293_ ( .A(\us00\/_0380_ ), .B(\us00\/_0347_ ), .X(\us00\/_0507_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1294_ ( .A1(\us00\/_0507_ ), .A2(\us00\/_0093_ ), .B1(\us00\/_0292_ ), .Y(\us00\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1295_ ( .A(\us00\/_0322_ ), .B(\us00\/_0277_ ), .C(\us00\/_0506_ ), .D(\us00\/_0508_ ), .X(\us00\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1296_ ( .A(\us00\/_0084_ ), .B(\us00\/_0705_ ), .X(\us00\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1297_ ( .A1(\us00\/_0733_ ), .A2(\us00\/_0114_ ), .B1(\us00\/_0429_ ), .C1(\us00\/_0511_ ), .Y(\us00\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_1298_ ( .A(\us00\/_0019_ ), .B(\us00\/_0024_ ), .Y(\us00\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1299_ ( .A(\us00\/_0512_ ), .B(\us00\/_0513_ ), .C(\us00\/_0742_ ), .D(\us00\/_0306_ ), .X(\us00\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1300_ ( .A1(\us00\/_0532_ ), .A2(\us00\/_0089_ ), .B1(\us00\/_0154_ ), .C1(\us00\/_0169_ ), .Y(\us00\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us00/_1301_ ( .A1(\us00\/_0749_ ), .A2(\us00\/_0026_ ), .B1(\us00\/_0069_ ), .C1(\us00\/_0032_ ), .X(\us00\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us00/_1302_ ( .A1(\us00\/_0324_ ), .A2(\us00\/_0355_ ), .B1(\us00\/_0330_ ), .B2(\us00\/_0727_ ), .X(\us00\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us00/_1303_ ( .A(\us00\/_0133_ ), .B(\us00\/_0516_ ), .C(\us00\/_0517_ ), .Y(\us00\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1304_ ( .A(\us00\/_0509_ ), .B(\us00\/_0514_ ), .C(\us00\/_0515_ ), .D(\us00\/_0518_ ), .X(\us00\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1305_ ( .A(\us00\/_0747_ ), .B(\us00\/_0072_ ), .Y(\us00\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1306_ ( .A1(\us00\/_0082_ ), .A2(\us00\/_0070_ ), .B1(\us00\/_0043_ ), .B2(\us00\/_0193_ ), .Y(\us00\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1307_ ( .A(\us00\/_0311_ ), .B(\us00\/_0520_ ), .C(\us00\/_0332_ ), .D(\us00\/_0522_ ), .X(\us00\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1308_ ( .A(\us00\/_0129_ ), .B(\us00\/_0218_ ), .X(\us00\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_1309_ ( .A(\us00\/_0235_ ), .B(\us00\/_0524_ ), .Y(\us00\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us00/_1310_ ( .A(\us00\/_0081_ ), .B(\us00\/_0085_ ), .Y(\us00\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1311_ ( .A1(\us00\/_0051_ ), .A2(\us00\/_0045_ ), .B1(\us00\/_0130_ ), .B2(\us00\/_0094_ ), .Y(\us00\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1312_ ( .A(\us00\/_0523_ ), .B(\us00\/_0525_ ), .C(\us00\/_0526_ ), .D(\us00\/_0527_ ), .X(\us00\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us00/_1313_ ( .A_N(\us00\/_0250_ ), .B(\us00\/_0521_ ), .Y(\us00\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1314_ ( .A(\us00\/_0128_ ), .B(\us00\/_0020_ ), .X(\us00\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1315_ ( .A(\us00\/_0530_ ), .Y(\us00\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1316_ ( .A(\us00\/_0099_ ), .B(\us00\/_0058_ ), .X(\us00\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1317_ ( .A(\us00\/_0533_ ), .Y(\us00\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us00/_1318_ ( .A_N(\us00\/_0529_ ), .B(\us00\/_0531_ ), .C(\us00\/_0534_ ), .D(\us00\/_0192_ ), .X(\us00\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1319_ ( .A(\us00\/_0434_ ), .B(\us00\/_0078_ ), .X(\us00\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us00/_1320_ ( .A1(\us00\/_0750_ ), .A2(\us00\/_0079_ ), .B1(\us00\/_0129_ ), .B2(\us00\/_0705_ ), .X(\us00\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1321_ ( .A1(\us00\/_0161_ ), .A2(\us00\/_0032_ ), .B1(\us00\/_0536_ ), .C1(\us00\/_0537_ ), .Y(\us00\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us00/_1322_ ( .A1(\us00\/_0747_ ), .A2(\us00\/_0162_ ), .B1(\us00\/_0079_ ), .B2(\us00\/_0043_ ), .X(\us00\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1323_ ( .A1(\us00\/_0093_ ), .A2(\us00\/_0247_ ), .B1(\us00\/_0240_ ), .C1(\us00\/_0539_ ), .Y(\us00\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1324_ ( .A(\us00\/_0434_ ), .B(\us00\/_0043_ ), .X(\us00\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us00/_1325_ ( .A1(\us00\/_0142_ ), .A2(\us00\/_0150_ ), .B1(\us00\/_0022_ ), .B2(\us00\/_0137_ ), .X(\us00\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1326_ ( .A1(\us00\/_0279_ ), .A2(\us00\/_0051_ ), .B1(\us00\/_0541_ ), .C1(\us00\/_0542_ ), .Y(\us00\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1327_ ( .A(\us00\/_0159_ ), .B(\us00\/_0035_ ), .X(\us00\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us00/_1328_ ( .A1(\us00\/_0271_ ), .A2(\us00\/_0434_ ), .B1(\us00\/_0027_ ), .X(\us00\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1329_ ( .A1(\us00\/_0091_ ), .A2(\us00\/_0128_ ), .B1(\us00\/_0545_ ), .C1(\us00\/_0546_ ), .Y(\us00\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1330_ ( .A(\us00\/_0538_ ), .B(\us00\/_0540_ ), .C(\us00\/_0544_ ), .D(\us00\/_0547_ ), .X(\us00\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1331_ ( .A(\us00\/_0099_ ), .B(\us00\/_0193_ ), .X(\us00\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us00/_1332_ ( .A(\us00\/_0549_ ), .B(\us00\/_0186_ ), .C(\us00\/_0187_ ), .Y(\us00\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1333_ ( .A(\us00\/_0062_ ), .B(\us00\/_0347_ ), .C(\us00\/_0749_ ), .D(\us00\/_0694_ ), .X(\us00\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1334_ ( .A1(\us00\/_0130_ ), .A2(\us00\/_0218_ ), .B1(\us00\/_0551_ ), .C1(\us00\/_0101_ ), .Y(\us00\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1335_ ( .A(\us00\/_0139_ ), .B(\us00\/_0640_ ), .Y(\us00\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1336_ ( .A1(\us00\/_0752_ ), .A2(\us00\/_0662_ ), .B1(\us00\/_0084_ ), .B2(\us00\/_0099_ ), .Y(\us00\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1337_ ( .A(\us00\/_0550_ ), .B(\us00\/_0552_ ), .C(\us00\/_0553_ ), .D(\us00\/_0555_ ), .X(\us00\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1338_ ( .A(\us00\/_0528_ ), .B(\us00\/_0535_ ), .C(\us00\/_0548_ ), .D(\us00\/_0556_ ), .X(\us00\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us00/_1339_ ( .A(\us00\/_0504_ ), .B(\us00\/_0519_ ), .C(\us00\/_0557_ ), .Y(\us00\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1340_ ( .A(\us00\/_0054_ ), .B(\us00\/_0507_ ), .X(\us00\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us00/_1341_ ( .A_N(\us00\/_0558_ ), .B(\us00\/_0408_ ), .C(\us00\/_0451_ ), .D(\us00\/_0452_ ), .X(\us00\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1342_ ( .A(\us00\/_0549_ ), .Y(\us00\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1343_ ( .A(\us00\/_0559_ ), .B(\us00\/_0403_ ), .C(\us00\/_0560_ ), .D(\us00\/_0371_ ), .X(\us00\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1344_ ( .A(\us00\/_0181_ ), .B(\us00\/_0178_ ), .X(\us00\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1345_ ( .A(\us00\/_0562_ ), .B(\us00\/_0552_ ), .C(\us00\/_0553_ ), .D(\us00\/_0555_ ), .X(\us00\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1346_ ( .A(\us00\/_0247_ ), .B(\us00\/_0020_ ), .Y(\us00\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1347_ ( .A(\us00\/_0051_ ), .B(\us00\/_0130_ ), .X(\us00\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1348_ ( .A(\us00\/_0566_ ), .Y(\us00\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1349_ ( .A(\us00\/_0159_ ), .B(\us00\/_0412_ ), .X(\us00\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1350_ ( .A1(\us00\/_0752_ ), .A2(\us00\/_0640_ ), .B1(\us00\/_0568_ ), .B2(\us00\/_0175_ ), .Y(\us00\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1351_ ( .A(\us00\/_0076_ ), .B(\us00\/_0565_ ), .C(\us00\/_0567_ ), .D(\us00\/_0569_ ), .X(\us00\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us00/_1352_ ( .A1(\us00\/_0035_ ), .A2(\us00\/_0142_ ), .B1(\us00\/_0161_ ), .X(\us00\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1353_ ( .A(\us00\/_0099_ ), .B(\us00\/_0662_ ), .Y(\us00\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us00/_1354_ ( .A(\us00\/_0420_ ), .B(\us00\/_0571_ ), .C_N(\us00\/_0572_ ), .Y(\us00\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1355_ ( .A(\us00\/_0051_ ), .B(\us00\/_0747_ ), .Y(\us00\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1356_ ( .A(\us00\/_0574_ ), .B(\us00\/_0319_ ), .C(\us00\/_0320_ ), .D(\us00\/_0411_ ), .X(\us00\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1357_ ( .A(\us00\/_0736_ ), .B(\us00\/_0035_ ), .Y(\us00\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1358_ ( .A(\us00\/_0736_ ), .B(\us00\/_0030_ ), .Y(\us00\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1359_ ( .A(\us00\/_0298_ ), .B(\us00\/_0208_ ), .C(\us00\/_0577_ ), .D(\us00\/_0578_ ), .X(\us00\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1360_ ( .A1(\us00\/_0020_ ), .A2(\us00\/_0137_ ), .B1(\us00\/_0261_ ), .B2(\us00\/_0128_ ), .Y(\us00\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1361_ ( .A(\us00\/_0573_ ), .B(\us00\/_0576_ ), .C(\us00\/_0579_ ), .D(\us00\/_0580_ ), .X(\us00\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1362_ ( .A(\us00\/_0561_ ), .B(\us00\/_0563_ ), .C(\us00\/_0570_ ), .D(\us00\/_0581_ ), .X(\us00\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1363_ ( .A(\us00\/_0128_ ), .B(\us00\/_0193_ ), .X(\us00\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1364_ ( .A(\us00\/_0082_ ), .B(\us00\/_0162_ ), .X(\us00\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us00/_1365_ ( .A(\us00\/_0583_ ), .B(\us00\/_0584_ ), .C_N(\us00\/_0437_ ), .Y(\us00\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us00/_1366_ ( .A(\us00\/_0150_ ), .B(\us00\/_0118_ ), .C(\us00\/_0380_ ), .Y(\us00\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us00/_1367_ ( .A_N(\us00\/_0182_ ), .B(\us00\/_0587_ ), .C(\us00\/_0323_ ), .X(\us00\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1368_ ( .A1(\us00\/_0575_ ), .A2(\us00\/_0153_ ), .B1(\us00\/_0727_ ), .B2(\us00\/_0058_ ), .Y(\us00\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1369_ ( .A1(\us00\/_0218_ ), .A2(\us00\/_0064_ ), .B1(\us00\/_0134_ ), .B2(\us00\/_0255_ ), .Y(\us00\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1370_ ( .A(\us00\/_0585_ ), .B(\us00\/_0588_ ), .C(\us00\/_0589_ ), .D(\us00\/_0590_ ), .X(\us00\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us00/_1371_ ( .A1(\us00\/_0091_ ), .A2(\us00\/_0139_ ), .B1(\us00\/_0250_ ), .Y(\us00\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1372_ ( .A1(\us00\/_0092_ ), .A2(\us00\/_0739_ ), .B1(\us00\/_0324_ ), .B2(\us00\/_0247_ ), .Y(\us00\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1373_ ( .A1(\us00\/_0144_ ), .A2(\us00\/_0153_ ), .B1(\us00\/_0683_ ), .B2(\us00\/_0292_ ), .Y(\us00\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1374_ ( .A1(\us00\/_0091_ ), .A2(\us00\/_0218_ ), .B1(\us00\/_0330_ ), .B2(\us00\/_0292_ ), .Y(\us00\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1375_ ( .A(\us00\/_0592_ ), .B(\us00\/_0593_ ), .C(\us00\/_0594_ ), .D(\us00\/_0595_ ), .X(\us00\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1376_ ( .A(\us00\/_0218_ ), .B(\us00\/_0144_ ), .Y(\us00\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1377_ ( .A(\us00\/_0312_ ), .B(\us00\/_0598_ ), .Y(\us00\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1378_ ( .A(\us00\/_0575_ ), .B(\us00\/_0147_ ), .Y(\us00\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1379_ ( .A1(\us00\/_0293_ ), .A2(\us00\/_0137_ ), .B1(\us00\/_0093_ ), .B2(\us00\/_0739_ ), .Y(\us00\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1380_ ( .A1(\us00\/_0734_ ), .A2(\us00\/_0531_ ), .B1(\us00\/_0600_ ), .C1(\us00\/_0601_ ), .Y(\us00\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1381_ ( .A1(\us00\/_0153_ ), .A2(\us00\/_0261_ ), .B1(\us00\/_0599_ ), .C1(\us00\/_0602_ ), .Y(\us00\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1382_ ( .A(\us00\/_0591_ ), .B(\us00\/_0596_ ), .C(\us00\/_0174_ ), .D(\us00\/_0603_ ), .X(\us00\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1383_ ( .A(\us00\/_0247_ ), .B(\us00\/_0144_ ), .Y(\us00\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1384_ ( .A(\us00\/_0113_ ), .B(\us00\/_0017_ ), .Y(\us00\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1385_ ( .A(\us00\/_0381_ ), .B(\us00\/_0605_ ), .C(\us00\/_0361_ ), .D(\us00\/_0606_ ), .X(\us00\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1386_ ( .A1(\us00\/_0016_ ), .A2(\us00\/_0727_ ), .B1(\us00\/_0733_ ), .Y(\us00\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1387_ ( .A1(\us00\/_0586_ ), .A2(\us00\/_0159_ ), .B1(\us00\/_0082_ ), .B2(\us00\/_0750_ ), .Y(\us00\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1388_ ( .A1(\us00\/_0142_ ), .A2(\us00\/_0162_ ), .B1(\us00\/_0079_ ), .B2(\us00\/_0054_ ), .Y(\us00\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1389_ ( .A(\us00\/_0610_ ), .B(\us00\/_0611_ ), .C(\us00\/_0105_ ), .D(\us00\/_0106_ ), .X(\us00\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1390_ ( .A1(\us00\/_0094_ ), .A2(\us00\/_0302_ ), .B1(\us00\/_0324_ ), .B2(\us00\/_0089_ ), .Y(\us00\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1391_ ( .A(\us00\/_0607_ ), .B(\us00\/_0609_ ), .C(\us00\/_0612_ ), .D(\us00\/_0613_ ), .X(\us00\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1392_ ( .A(\us00\/_0041_ ), .B(\us00\/_0170_ ), .X(\us00\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1393_ ( .A(\us00\/_0554_ ), .B(\us00\/_0027_ ), .X(\us00\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1394_ ( .A(\us00\/_0027_ ), .B(\us00\/_0261_ ), .Y(\us00\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us00/_1395_ ( .A_N(\us00\/_0616_ ), .B(\us00\/_0617_ ), .Y(\us00\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1396_ ( .A1(\us00\/_0147_ ), .A2(\us00\/_0302_ ), .B1(\us00\/_0342_ ), .C1(\us00\/_0618_ ), .Y(\us00\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1397_ ( .A(\us00\/_0614_ ), .B(\us00\/_0272_ ), .C(\us00\/_0615_ ), .D(\us00\/_0620_ ), .X(\us00\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us00/_1398_ ( .A(\us00\/_0582_ ), .B(\us00\/_0604_ ), .C(\us00\/_0621_ ), .Y(\us00\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1399_ ( .A1(\us00\/_0084_ ), .A2(\us00\/_0134_ ), .B1(\us00\/_0089_ ), .Y(\us00\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1400_ ( .A1(\us00\/_0144_ ), .A2(\us00\/_0608_ ), .A3(\us00\/_0330_ ), .B1(\us00\/_0089_ ), .Y(\us00\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1401_ ( .A1(\us00\/_0197_ ), .A2(\us00\/_0130_ ), .A3(\us00\/_0110_ ), .B1(\us00\/_0094_ ), .Y(\us00\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1402_ ( .A(\us00\/_0432_ ), .B(\us00\/_0622_ ), .C(\us00\/_0623_ ), .D(\us00\/_0624_ ), .X(\us00\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us00/_1403_ ( .A1(\us00\/_0554_ ), .A2(\us00\/_0017_ ), .A3(\us00\/_0022_ ), .B1(\us00\/_0161_ ), .X(\us00\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us00/_1404_ ( .A_N(\us00\/_0269_ ), .B(\us00\/_0170_ ), .X(\us00\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1405_ ( .A1(\us00\/_0109_ ), .A2(\us00\/_0064_ ), .A3(\us00\/_0733_ ), .B1(\us00\/_0355_ ), .Y(\us00\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us00/_1406_ ( .A_N(\us00\/_0626_ ), .B(\us00\/_0627_ ), .C(\us00\/_0353_ ), .D(\us00\/_0628_ ), .X(\us00\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1407_ ( .A1(\us00\/_0091_ ), .A2(\us00\/_0110_ ), .A3(\us00\/_0176_ ), .B1(\us00\/_0139_ ), .Y(\us00\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1408_ ( .A1(\us00\/_0020_ ), .A2(\us00\/_0261_ ), .B1(\us00\/_0147_ ), .Y(\us00\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1409_ ( .A(\us00\/_0631_ ), .B(\us00\/_0344_ ), .C(\us00\/_0421_ ), .D(\us00\/_0632_ ), .X(\us00\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us00/_1410_ ( .A1(\us00\/_0325_ ), .A2(\us00\/_0734_ ), .B1(\us00\/_0038_ ), .C1(\us00\/_0113_ ), .X(\us00\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1411_ ( .A1(\us00\/_0134_ ), .A2(\us00\/_0114_ ), .B1(\us00\/_0221_ ), .C1(\us00\/_0634_ ), .Y(\us00\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us00/_1412_ ( .A(\us00\/_0119_ ), .B_N(\us00\/_0111_ ), .Y(\us00\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1413_ ( .A1(\us00\/_0032_ ), .A2(\us00\/_0113_ ), .B1(\us00\/_0636_ ), .C1(\us00\/_0400_ ), .Y(\us00\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1414_ ( .A1(\us00\/_0732_ ), .A2(\us00\/_0293_ ), .A3(\us00\/_0251_ ), .B1(\us00\/_0099_ ), .Y(\us00\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1415_ ( .A(\us00\/_0189_ ), .B(\us00\/_0635_ ), .C(\us00\/_0637_ ), .D(\us00\/_0638_ ), .X(\us00\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1416_ ( .A(\us00\/_0625_ ), .B(\us00\/_0630_ ), .C(\us00\/_0633_ ), .D(\us00\/_0639_ ), .X(\us00\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1417_ ( .A(\us00\/_0747_ ), .B(\us00\/_0738_ ), .X(\us00\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1418_ ( .A(\us00\/_0736_ ), .B(\us00\/_0731_ ), .X(\us00\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us00/_1419_ ( .A_N(\us00\/_0643_ ), .B(\us00\/_0577_ ), .Y(\us00\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1420_ ( .A1(\us00\/_0084_ ), .A2(\us00\/_0739_ ), .B1(\us00\/_0642_ ), .C1(\us00\/_0644_ ), .Y(\us00\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1421_ ( .A1(\us00\/_0050_ ), .A2(\us00\/_0249_ ), .B1(\us00\/_0194_ ), .C1(\us00\/_0738_ ), .Y(\us00\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1422_ ( .A(\us00\/_0646_ ), .B(\us00\/_0232_ ), .C(\us00\/_0417_ ), .D(\us00\/_0578_ ), .X(\us00\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1423_ ( .A1(\us00\/_0064_ ), .A2(\us00\/_0733_ ), .B1(\us00\/_0727_ ), .Y(\us00\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1424_ ( .A1(\us00\/_0193_ ), .A2(\us00\/_0276_ ), .B1(\us00\/_0727_ ), .Y(\us00\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1425_ ( .A(\us00\/_0645_ ), .B(\us00\/_0647_ ), .C(\us00\/_0648_ ), .D(\us00\/_0649_ ), .X(\us00\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1426_ ( .A1(\us00\/_0325_ ), .A2(\us00\/_0734_ ), .B1(\us00\/_0038_ ), .C1(\us00\/_0247_ ), .Y(\us00\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1427_ ( .A1(\us00\/_0249_ ), .A2(\us00\/_0205_ ), .B1(\us00\/_0412_ ), .C1(\us00\/_0247_ ), .Y(\us00\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1428_ ( .A(\us00\/_0652_ ), .B(\us00\/_0653_ ), .X(\us00\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1429_ ( .A1(\us00\/_0733_ ), .A2(\us00\/_0748_ ), .A3(\us00\/_0324_ ), .B1(\us00\/_0016_ ), .Y(\us00\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1430_ ( .A1(\us00\/_0640_ ), .A2(\us00\/_0193_ ), .A3(\us00\/_0091_ ), .B1(\us00\/_0016_ ), .Y(\us00\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1431_ ( .A1(\us00\/_0102_ ), .A2(\us00\/_0301_ ), .B1(\sa00\[3\] ), .C1(\us00\/_0247_ ), .Y(\us00\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1432_ ( .A(\us00\/_0654_ ), .B(\us00\/_0655_ ), .C(\us00\/_0656_ ), .D(\us00\/_0657_ ), .X(\us00\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1433_ ( .A1(\us00\/_0118_ ), .A2(\us00\/_0050_ ), .B1(\us00\/_0038_ ), .C1(\us00\/_0478_ ), .Y(\us00\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us00/_1434_ ( .A_N(\us00\/_0250_ ), .B(\us00\/_0465_ ), .C(\us00\/_0659_ ), .X(\us00\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1435_ ( .A1(\us00\/_0683_ ), .A2(\us00\/_0324_ ), .B1(\us00\/_0255_ ), .Y(\us00\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1436_ ( .A1(\us00\/_0032_ ), .A2(\us00\/_0193_ ), .A3(\us00\/_0047_ ), .B1(\us00\/_0255_ ), .Y(\us00\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1437_ ( .A1(\us00\/_0144_ ), .A2(\us00\/_0586_ ), .A3(\us00\/_0047_ ), .B1(\us00\/_0218_ ), .Y(\us00\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1438_ ( .A(\us00\/_0660_ ), .B(\us00\/_0661_ ), .C(\us00\/_0663_ ), .D(\us00\/_0664_ ), .X(\us00\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1439_ ( .A1(\us00\/_0091_ ), .A2(\us00\/_0276_ ), .B1(\us00\/_0060_ ), .Y(\us00\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1440_ ( .A1(\us00\/_0144_ ), .A2(\us00\/_0608_ ), .B1(\us00\/_0292_ ), .Y(\us00\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1441_ ( .A1(\us00\/_0412_ ), .A2(\us00\/_0038_ ), .B1(\us00\/_0102_ ), .C1(\us00\/_0060_ ), .Y(\us00\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1442_ ( .A1(\sa00\[1\] ), .A2(\us00\/_0734_ ), .B1(\us00\/_0109_ ), .C1(\us00\/_0292_ ), .Y(\us00\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1443_ ( .A(\us00\/_0666_ ), .B(\us00\/_0667_ ), .C(\us00\/_0668_ ), .D(\us00\/_0669_ ), .X(\us00\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1444_ ( .A(\us00\/_0650_ ), .B(\us00\/_0658_ ), .C(\us00\/_0665_ ), .D(\us00\/_0670_ ), .X(\us00\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us00/_1445_ ( .A(\us00\/_0641_ ), .B(\us00\/_0174_ ), .C(\us00\/_0671_ ), .Y(\us00\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us00/_1446_ ( .A(\us00\/_0049_ ), .B(\us00\/_0618_ ), .C_N(\us00\/_0052_ ), .Y(\us00\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us00/_1447_ ( .A(\us00\/_0239_ ), .Y(\us00\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1448_ ( .A(\us00\/_0705_ ), .B(\us00\/_0032_ ), .Y(\us00\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1449_ ( .A1(\us00\/_0054_ ), .A2(\us00\/_0732_ ), .B1(\us00\/_0035_ ), .B2(\us00\/_0705_ ), .Y(\us00\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1450_ ( .A1(\us00\/_0304_ ), .A2(\us00\/_0732_ ), .B1(\us00\/_0047_ ), .B2(\us00\/_0750_ ), .Y(\us00\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1451_ ( .A(\us00\/_0674_ ), .B(\us00\/_0675_ ), .C(\us00\/_0676_ ), .D(\us00\/_0677_ ), .X(\us00\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us00/_1452_ ( .A_N(\us00\/_0584_ ), .B(\us00\/_0283_ ), .X(\us00\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1453_ ( .A(\us00\/_0673_ ), .B(\us00\/_0678_ ), .C(\us00\/_0679_ ), .D(\us00\/_0508_ ), .X(\us00\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1454_ ( .A1(\us00\/_0016_ ), .A2(\us00\/_0733_ ), .B1(\us00\/_0355_ ), .B2(\us00\/_0092_ ), .Y(\us00\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1455_ ( .A(\us00\/_0681_ ), .B(\us00\/_0034_ ), .X(\us00\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us00/_1456_ ( .A1(\us00\/_0330_ ), .A2(\us00\/_0139_ ), .B1(\us00\/_0324_ ), .B2(\us00\/_0089_ ), .X(\us00\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1457_ ( .A1(\us00\/_0146_ ), .A2(\us00\/_0147_ ), .B1(\us00\/_0133_ ), .C1(\us00\/_0684_ ), .Y(\us00\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1458_ ( .A(\us00\/_0113_ ), .B(\us00\/_0251_ ), .Y(\us00\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us00/_1459_ ( .A_N(\us00\/_0463_ ), .B(\us00\/_0686_ ), .C(\us00\/_0383_ ), .D(\us00\/_0464_ ), .X(\us00\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1460_ ( .A1(\us00\/_0051_ ), .A2(\us00\/_0293_ ), .B1(\us00\/_0084_ ), .B2(\us00\/_0705_ ), .Y(\us00\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1461_ ( .A1(\us00\/_0017_ ), .A2(\us00\/_0072_ ), .B1(\us00\/_0134_ ), .B2(\us00\/_0078_ ), .Y(\us00\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1462_ ( .A(\us00\/_0687_ ), .B(\us00\/_0236_ ), .C(\us00\/_0688_ ), .D(\us00\/_0689_ ), .X(\us00\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1463_ ( .A(\us00\/_0680_ ), .B(\us00\/_0682_ ), .C(\us00\/_0685_ ), .D(\us00\/_0690_ ), .X(\us00\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us00/_1464_ ( .A1(\us00\/_0532_ ), .A2(\us00\/_0380_ ), .B1(\us00\/_0102_ ), .C1(\us00\/_0355_ ), .X(\us00\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us00/_1465_ ( .A(\us00\/_0692_ ), .B(\us00\/_0338_ ), .C(\us00\/_0644_ ), .Y(\us00\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1466_ ( .A(\us00\/_0016_ ), .B(\us00\/_0020_ ), .Y(\us00\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1467_ ( .A1(\us00\/_0032_ ), .A2(\us00\/_0137_ ), .B1(\us00\/_0279_ ), .B2(\us00\/_0094_ ), .Y(\us00\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1468_ ( .A1(\us00\/_0575_ ), .A2(\us00\/_0153_ ), .B1(\us00\/_0161_ ), .B2(\us00\/_0293_ ), .Y(\us00\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1469_ ( .A(\us00\/_0259_ ), .B(\us00\/_0695_ ), .C(\us00\/_0696_ ), .D(\us00\/_0697_ ), .X(\us00\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us00/_1470_ ( .A1(\us00\/_0255_ ), .A2(\us00\/_0640_ ), .B1(\us00\/_0016_ ), .B2(\us00\/_0193_ ), .X(\us00\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1471_ ( .A1(\us00\/_0060_ ), .A2(\us00\/_0176_ ), .B1(\us00\/_0699_ ), .C1(\us00\/_0177_ ), .Y(\us00\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1472_ ( .A1(\us00\/_0091_ ), .A2(\us00\/_0218_ ), .B1(\us00\/_0092_ ), .B2(\us00\/_0705_ ), .Y(\us00\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us00/_1473_ ( .A1(\us00\/_0705_ ), .A2(\us00\/_0683_ ), .B1(\us00\/_0093_ ), .B2(\us00\/_0114_ ), .Y(\us00\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us00/_1474_ ( .A1(\us00\/_0683_ ), .A2(\us00\/_0084_ ), .B1(\us00\/_0094_ ), .Y(\us00\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us00/_1475_ ( .A1(\us00\/_0249_ ), .A2(\us00\/_0205_ ), .B1(\us00\/_0038_ ), .C1(\us00\/_0292_ ), .Y(\us00\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1476_ ( .A(\us00\/_0701_ ), .B(\us00\/_0702_ ), .C(\us00\/_0703_ ), .D(\us00\/_0704_ ), .X(\us00\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1477_ ( .A(\us00\/_0693_ ), .B(\us00\/_0698_ ), .C(\us00\/_0700_ ), .D(\us00\/_0706_ ), .X(\us00\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us00/_1478_ ( .A1(\us00\/_0113_ ), .A2(\us00\/_0640_ ), .B1(\us00\/_0099_ ), .B2(\us00\/_0058_ ), .X(\us00\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us00/_1479_ ( .A(\us00\/_0407_ ), .B(\us00\/_0708_ ), .C(\us00\/_0529_ ), .Y(\us00\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1480_ ( .A(\us00\/_0568_ ), .B(\us00\/_0175_ ), .Y(\us00\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us00/_1481_ ( .A1(\us00\/_0247_ ), .A2(\us00\/_0114_ ), .A3(\us00\/_0051_ ), .B1(\us00\/_0130_ ), .Y(\us00\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1482_ ( .A(\us00\/_0709_ ), .B(\us00\/_0550_ ), .C(\us00\/_0710_ ), .D(\us00\/_0711_ ), .X(\us00\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us00/_1483_ ( .A1(\us00\/_0114_ ), .A2(\us00\/_0064_ ), .B1(\us00\/_0261_ ), .B2(\us00\/_0089_ ), .X(\us00\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1484_ ( .A1(\us00\/_0355_ ), .A2(\us00\/_0261_ ), .B1(\us00\/_0198_ ), .C1(\us00\/_0713_ ), .Y(\us00\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1485_ ( .A(\us00\/_0586_ ), .B(\us00\/_0478_ ), .Y(\us00\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us00/_1486_ ( .A_N(\us00\/_0541_ ), .B(\us00\/_0267_ ), .C(\us00\/_0715_ ), .D(\us00\/_0320_ ), .X(\us00\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1487_ ( .A(\us00\/_0586_ ), .B(\us00\/_0070_ ), .Y(\us00\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us00/_1488_ ( .A_N(\us00\/_0211_ ), .B(\us00\/_0155_ ), .C(\us00\/_0202_ ), .D(\us00\/_0718_ ), .X(\us00\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us00/_1489_ ( .A(\us00\/_0150_ ), .B(\us00\/_0205_ ), .C(\us00\/_0380_ ), .Y(\us00\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us00/_1490_ ( .A(\us00\/_0411_ ), .B(\us00\/_0720_ ), .X(\us00\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us00/_1491_ ( .A1(\us00\/_0017_ ), .A2(\us00\/_0022_ ), .B1(\us00\/_0078_ ), .X(\us00\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us00/_1492_ ( .A1(\us00\/_0134_ ), .A2(\us00\/_0738_ ), .B1(\us00\/_0101_ ), .C1(\us00\/_0722_ ), .Y(\us00\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1493_ ( .A(\us00\/_0717_ ), .B(\us00\/_0719_ ), .C(\us00\/_0721_ ), .D(\us00\/_0723_ ), .X(\us00\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us00/_1494_ ( .A(\us00\/_0739_ ), .B(\us00\/_0193_ ), .Y(\us00\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1495_ ( .A(\us00\/_0344_ ), .B(\us00\/_0184_ ), .C(\us00\/_0449_ ), .D(\us00\/_0725_ ), .X(\us00\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us00/_1496_ ( .A(\us00\/_0712_ ), .B(\us00\/_0714_ ), .C(\us00\/_0724_ ), .D(\us00\/_0726_ ), .X(\us00\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \us00/_1497_ ( .A(\us00\/_0691_ ), .B(\us00\/_0707_ ), .C(\us00\/_0728_ ), .Y(\us00\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \us01/_0753_ ( .A(\sa01\[2\] ), .B_N(\sa01\[3\] ), .Y(\us01\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \us01/_0755_ ( .A(\sa01\[1\] ), .B(\sa01\[0\] ), .X(\us01\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us01/_0756_ ( .A(\us01\/_0096_ ), .B(\us01\/_0118_ ), .X(\us01\/_0129_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0757_ ( .A(\sa01\[7\] ), .B(\sa01\[6\] ), .X(\us01\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_0758_ ( .A(\sa01\[4\] ), .B(\sa01\[5\] ), .Y(\us01\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0759_ ( .A(\us01\/_0140_ ), .B(\us01\/_0151_ ), .X(\us01\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0761_ ( .A(\us01\/_0129_ ), .B(\us01\/_0162_ ), .X(\us01\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0762_ ( .A(\us01\/_0096_ ), .X(\us01\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \us01/_0763_ ( .A(\sa01\[1\] ), .B_N(\sa01\[0\] ), .Y(\us01\/_0205_ ) );
sky130_fd_sc_hd__and3_1 \us01/_0765_ ( .A(\us01\/_0162_ ), .B(\us01\/_0194_ ), .C(\us01\/_0205_ ), .X(\us01\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us01/_0766_ ( .A(\us01\/_0183_ ), .SLEEP(\us01\/_0227_ ), .X(\us01\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \us01/_0767_ ( .A(\sa01\[0\] ), .B_N(\sa01\[1\] ), .Y(\us01\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_0768_ ( .A(\sa01\[2\] ), .B(\sa01\[3\] ), .Y(\us01\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0769_ ( .A(\us01\/_0249_ ), .B(\us01\/_0260_ ), .X(\us01\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0771_ ( .A(\us01\/_0271_ ), .X(\us01\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0772_ ( .A(\us01\/_0162_ ), .X(\us01\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_0773_ ( .A(\us01\/_0293_ ), .B(\us01\/_0304_ ), .Y(\us01\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us01/_0774_ ( .A(\sa01\[1\] ), .Y(\us01\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us01/_0776_ ( .A(\sa01\[0\] ), .Y(\us01\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0777_ ( .A(\sa01\[2\] ), .B(\sa01\[3\] ), .X(\us01\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0779_ ( .A(\us01\/_0358_ ), .X(\us01\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_0780_ ( .A1(\us01\/_0325_ ), .A2(\us01\/_0347_ ), .B1(\us01\/_0380_ ), .C1(\us01\/_0304_ ), .Y(\us01\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us01/_0781_ ( .A_N(\us01\/_0238_ ), .B(\us01\/_0314_ ), .C(\us01\/_0391_ ), .X(\us01\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us01/_0782_ ( .A(\sa01\[3\] ), .B_N(\sa01\[2\] ), .Y(\us01\/_0412_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0784_ ( .A(\us01\/_0412_ ), .B(\us01\/_0205_ ), .X(\us01\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \us01/_0787_ ( .A(\sa01\[5\] ), .B_N(\sa01\[4\] ), .Y(\us01\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0788_ ( .A(\us01\/_0467_ ), .B(\us01\/_0140_ ), .X(\us01\/_0478_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_0791_ ( .A(\us01\/_0134_ ), .B(\us01\/_0218_ ), .Y(\us01\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_0792_ ( .A(\us01\/_0478_ ), .B(\us01\/_0271_ ), .Y(\us01\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0793_ ( .A(\us01\/_0194_ ), .X(\us01\/_0532_ ) );
sky130_fd_sc_hd__and2_1 \us01/_0795_ ( .A(\us01\/_0249_ ), .B(\us01\/_0358_ ), .X(\us01\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0797_ ( .A(\us01\/_0554_ ), .X(\us01\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us01/_0798_ ( .A(\us01\/_0205_ ), .B(\us01\/_0358_ ), .X(\us01\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0800_ ( .A(\us01\/_0586_ ), .X(\us01\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_0801_ ( .A1(\us01\/_0532_ ), .A2(\us01\/_0575_ ), .A3(\us01\/_0608_ ), .B1(\us01\/_0218_ ), .Y(\us01\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us01/_0802_ ( .A(\us01\/_0401_ ), .B(\us01\/_0510_ ), .C(\us01\/_0521_ ), .D(\us01\/_0619_ ), .X(\us01\/_0629_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0803_ ( .A(\us01\/_0358_ ), .B(\sa01\[1\] ), .X(\us01\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0805_ ( .A(\us01\/_0205_ ), .B(\us01\/_0260_ ), .X(\us01\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0807_ ( .A(\us01\/_0662_ ), .X(\us01\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us01/_0808_ ( .A(\sa01\[6\] ), .B_N(\sa01\[7\] ), .Y(\us01\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \us01/_0809_ ( .A(\us01\/_0467_ ), .B(\us01\/_0694_ ), .X(\us01\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0811_ ( .A(\us01\/_0705_ ), .X(\us01\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_0812_ ( .A1(\us01\/_0640_ ), .A2(\us01\/_0293_ ), .A3(\us01\/_0683_ ), .B1(\us01\/_0727_ ), .Y(\us01\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_0813_ ( .A(\sa01\[1\] ), .B(\sa01\[0\] ), .Y(\us01\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0814_ ( .A(\us01\/_0730_ ), .B(\us01\/_0260_ ), .X(\us01\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0816_ ( .A(\us01\/_0731_ ), .X(\us01\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0817_ ( .A(\sa01\[0\] ), .X(\us01\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us01/_0818_ ( .A1(\us01\/_0325_ ), .A2(\us01\/_0734_ ), .B1(\us01\/_0412_ ), .X(\us01\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0819_ ( .A(\us01\/_0694_ ), .B(\us01\/_0151_ ), .X(\us01\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0821_ ( .A(\us01\/_0736_ ), .X(\us01\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0822_ ( .A(\us01\/_0738_ ), .X(\us01\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_0823_ ( .A1(\us01\/_0733_ ), .A2(\us01\/_0735_ ), .A3(\us01\/_0293_ ), .B1(\us01\/_0739_ ), .Y(\us01\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us01/_0824_ ( .A(\us01\/_0730_ ), .B_N(\us01\/_0358_ ), .Y(\us01\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_0825_ ( .A(\us01\/_0741_ ), .B(\us01\/_0739_ ), .Y(\us01\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_0827_ ( .A1(\us01\/_0118_ ), .A2(\us01\/_0205_ ), .B1(\us01\/_0532_ ), .C1(\us01\/_0739_ ), .Y(\us01\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us01/_0828_ ( .A(\us01\/_0729_ ), .B(\us01\/_0740_ ), .C(\us01\/_0742_ ), .D(\us01\/_0744_ ), .X(\us01\/_0745_ ) );
sky130_fd_sc_hd__and2_1 \us01/_0829_ ( .A(\us01\/_0412_ ), .B(\us01\/_0730_ ), .X(\us01\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0831_ ( .A(\us01\/_0746_ ), .X(\us01\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us01/_0832_ ( .A(\sa01\[4\] ), .B_N(\sa01\[5\] ), .Y(\us01\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0833_ ( .A(\us01\/_0749_ ), .B(\us01\/_0694_ ), .X(\us01\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0835_ ( .A(\us01\/_0750_ ), .X(\us01\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0836_ ( .A(\us01\/_0752_ ), .X(\us01\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0837_ ( .A(\us01\/_0118_ ), .B(\us01\/_0358_ ), .X(\us01\/_0017_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0839_ ( .A(\us01\/_0752_ ), .B(\us01\/_0017_ ), .X(\us01\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0840_ ( .A(\us01\/_0358_ ), .B(\us01\/_0325_ ), .X(\us01\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0842_ ( .A(\us01\/_0096_ ), .B(\us01\/_0205_ ), .X(\us01\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \us01/_0844_ ( .A1(\us01\/_0020_ ), .A2(\us01\/_0022_ ), .B1(\us01\/_0752_ ), .X(\us01\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_0845_ ( .A1(\us01\/_0748_ ), .A2(\us01\/_0016_ ), .B1(\us01\/_0019_ ), .C1(\us01\/_0024_ ), .Y(\us01\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \us01/_0846_ ( .A(\sa01\[4\] ), .B(\sa01\[5\] ), .X(\us01\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0847_ ( .A(\us01\/_0694_ ), .B(\us01\/_0026_ ), .X(\us01\/_0027_ ) );
sky130_fd_sc_hd__buf_2 \us01/_0849_ ( .A(\us01\/_0027_ ), .X(\us01\/_0029_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0850_ ( .A(\us01\/_0358_ ), .B(\us01\/_0730_ ), .X(\us01\/_0030_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_0853_ ( .A(\us01\/_0029_ ), .B(\us01\/_0030_ ), .Y(\us01\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_0854_ ( .A(\us01\/_0029_ ), .B(\us01\/_0735_ ), .Y(\us01\/_0034_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0855_ ( .A(\us01\/_0118_ ), .B(\us01\/_0260_ ), .X(\us01\/_0035_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0857_ ( .A(\us01\/_0027_ ), .B(\us01\/_0035_ ), .X(\us01\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0858_ ( .A(\us01\/_0260_ ), .X(\us01\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_0859_ ( .A(\us01\/_0038_ ), .B(\us01\/_0347_ ), .Y(\us01\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us01/_0860_ ( .A_N(\us01\/_0039_ ), .B(\us01\/_0027_ ), .X(\us01\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_0861_ ( .A(\us01\/_0037_ ), .B(\us01\/_0040_ ), .Y(\us01\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us01/_0862_ ( .A(\us01\/_0025_ ), .B(\us01\/_0033_ ), .C(\us01\/_0034_ ), .D(\us01\/_0041_ ), .X(\us01\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0863_ ( .A(\us01\/_0749_ ), .B(\us01\/_0140_ ), .X(\us01\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us01/_0865_ ( .A(\sa01\[0\] ), .B(\sa01\[2\] ), .C(\sa01\[3\] ), .X(\us01\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0866_ ( .A(\us01\/_0043_ ), .B(\us01\/_0045_ ), .X(\us01\/_0046_ ) );
sky130_fd_sc_hd__and2_1 \us01/_0867_ ( .A(\us01\/_0096_ ), .B(\us01\/_0249_ ), .X(\us01\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0869_ ( .A(\us01\/_0047_ ), .B(\us01\/_0043_ ), .X(\us01\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0870_ ( .A(\us01\/_0730_ ), .X(\us01\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0871_ ( .A(\us01\/_0043_ ), .X(\us01\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_0872_ ( .A1(\us01\/_0118_ ), .A2(\us01\/_0050_ ), .B1(\us01\/_0194_ ), .C1(\us01\/_0051_ ), .Y(\us01\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us01/_0873_ ( .A(\us01\/_0046_ ), .B(\us01\/_0049_ ), .C_N(\us01\/_0052_ ), .Y(\us01\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0874_ ( .A(\us01\/_0026_ ), .B(\us01\/_0140_ ), .X(\us01\/_0054_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_0877_ ( .A1(\us01\/_0532_ ), .A2(\us01\/_0575_ ), .B1(\us01\/_0292_ ), .Y(\us01\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0878_ ( .A(\us01\/_0412_ ), .B(\us01\/_0325_ ), .X(\us01\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0880_ ( .A(\us01\/_0051_ ), .X(\us01\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_0881_ ( .A1(\us01\/_0731_ ), .A2(\us01\/_0035_ ), .A3(\us01\/_0058_ ), .B1(\us01\/_0060_ ), .Y(\us01\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0882_ ( .A(\us01\/_0260_ ), .B(\sa01\[1\] ), .X(\us01\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0884_ ( .A(\us01\/_0062_ ), .X(\us01\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_0885_ ( .A1(\us01\/_0064_ ), .A2(\us01\/_0748_ ), .A3(\us01\/_0683_ ), .B1(\us01\/_0292_ ), .Y(\us01\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us01/_0886_ ( .A(\us01\/_0053_ ), .B(\us01\/_0057_ ), .C(\us01\/_0061_ ), .D(\us01\/_0065_ ), .X(\us01\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us01/_0887_ ( .A(\us01\/_0629_ ), .B(\us01\/_0745_ ), .C(\us01\/_0042_ ), .D(\us01\/_0066_ ), .X(\us01\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us01/_0889_ ( .A(\sa01\[7\] ), .B_N(\sa01\[6\] ), .Y(\us01\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0890_ ( .A(\us01\/_0069_ ), .B(\us01\/_0151_ ), .X(\us01\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0892_ ( .A(\us01\/_0070_ ), .X(\us01\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_0893_ ( .A1(\us01\/_0129_ ), .A2(\us01\/_0586_ ), .B1(\us01\/_0072_ ), .Y(\us01\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_0894_ ( .A1(\us01\/_0380_ ), .A2(\us01\/_0347_ ), .B1(\us01\/_0194_ ), .B2(\us01\/_0205_ ), .Y(\us01\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us01/_0895_ ( .A(\us01\/_0074_ ), .B_N(\us01\/_0070_ ), .Y(\us01\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us01/_0896_ ( .A(\us01\/_0073_ ), .SLEEP(\us01\/_0075_ ), .X(\us01\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us01/_0897_ ( .A(\us01\/_0467_ ), .B(\us01\/_0069_ ), .X(\us01\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0898_ ( .A(\us01\/_0077_ ), .X(\us01\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0899_ ( .A(\us01\/_0412_ ), .B(\us01\/_0118_ ), .X(\us01\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0901_ ( .A(\us01\/_0078_ ), .B(\us01\/_0079_ ), .X(\us01\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0902_ ( .A(\us01\/_0412_ ), .B(\us01\/_0249_ ), .X(\us01\/_0082_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0905_ ( .A(\us01\/_0280_ ), .B(\us01\/_0078_ ), .X(\us01\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us01/_0906_ ( .A1(\sa01\[0\] ), .A2(\us01\/_0325_ ), .B1(\us01\/_0260_ ), .Y(\us01\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us01/_0907_ ( .A_N(\us01\/_0086_ ), .B(\us01\/_0078_ ), .X(\us01\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us01/_0908_ ( .A(\us01\/_0081_ ), .B(\us01\/_0085_ ), .C(\us01\/_0087_ ), .Y(\us01\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0909_ ( .A(\us01\/_0072_ ), .X(\us01\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_0910_ ( .A1(\us01\/_0733_ ), .A2(\us01\/_0748_ ), .A3(\us01\/_0683_ ), .B1(\us01\/_0089_ ), .Y(\us01\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0911_ ( .A(\us01\/_0129_ ), .X(\us01\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0912_ ( .A(\us01\/_0017_ ), .X(\us01\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0913_ ( .A(\us01\/_0022_ ), .X(\us01\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0914_ ( .A(\us01\/_0078_ ), .X(\us01\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_0915_ ( .A1(\us01\/_0091_ ), .A2(\us01\/_0092_ ), .A3(\us01\/_0093_ ), .B1(\us01\/_0094_ ), .Y(\us01\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us01/_0916_ ( .A(\us01\/_0076_ ), .B(\us01\/_0088_ ), .C(\us01\/_0090_ ), .D(\us01\/_0095_ ), .X(\us01\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us01/_0917_ ( .A(\us01\/_0069_ ), .B(\us01\/_0026_ ), .X(\us01\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \us01/_0918_ ( .A(\us01\/_0098_ ), .X(\us01\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0919_ ( .A(\us01\/_0434_ ), .B(\us01\/_0099_ ), .X(\us01\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0920_ ( .A(\us01\/_0079_ ), .B(\us01\/_0098_ ), .X(\us01\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0921_ ( .A(\us01\/_0325_ ), .X(\us01\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_0922_ ( .A1(\us01\/_0102_ ), .A2(\us01\/_0734_ ), .B1(\us01\/_0038_ ), .C1(\us01\/_0099_ ), .Y(\us01\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us01/_0923_ ( .A(\us01\/_0100_ ), .B(\us01\/_0101_ ), .C_N(\us01\/_0103_ ), .Y(\us01\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_0924_ ( .A1(\us01\/_0554_ ), .A2(\us01\/_0586_ ), .B1(\us01\/_0099_ ), .Y(\us01\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_0925_ ( .A(\us01\/_0129_ ), .B(\us01\/_0099_ ), .Y(\us01\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0926_ ( .A(\us01\/_0105_ ), .B(\us01\/_0106_ ), .X(\us01\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0927_ ( .A(\us01\/_0412_ ), .X(\us01\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us01/_0928_ ( .A(\us01\/_0260_ ), .B(\sa01\[0\] ), .X(\us01\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0929_ ( .A(\us01\/_0069_ ), .B(\us01\/_0749_ ), .X(\us01\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0931_ ( .A(\us01\/_0111_ ), .X(\us01\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0932_ ( .A(\us01\/_0113_ ), .X(\us01\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_0933_ ( .A1(\us01\/_0109_ ), .A2(\us01\/_0110_ ), .B1(\us01\/_0114_ ), .Y(\us01\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us01/_0934_ ( .A(\us01\/_0022_ ), .Y(\us01\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us01/_0935_ ( .A(\us01\/_0554_ ), .Y(\us01\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us01/_0936_ ( .A1(\us01\/_0050_ ), .A2(\us01\/_0118_ ), .B1(\us01\/_0194_ ), .Y(\us01\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us01/_0937_ ( .A(\us01\/_0113_ ), .Y(\us01\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us01/_0938_ ( .A1(\us01\/_0116_ ), .A2(\us01\/_0117_ ), .A3(\us01\/_0119_ ), .B1(\us01\/_0120_ ), .X(\us01\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us01/_0939_ ( .A(\us01\/_0104_ ), .B(\us01\/_0108_ ), .C(\us01\/_0115_ ), .D(\us01\/_0121_ ), .X(\us01\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_0940_ ( .A(\sa01\[7\] ), .B(\sa01\[6\] ), .Y(\us01\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0941_ ( .A(\us01\/_0749_ ), .B(\us01\/_0123_ ), .X(\us01\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0943_ ( .A(\us01\/_0082_ ), .B(\us01\/_0124_ ), .X(\us01\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_0944_ ( .A(\us01\/_0271_ ), .B(\us01\/_0124_ ), .Y(\us01\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0945_ ( .A(\us01\/_0124_ ), .X(\us01\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0946_ ( .A(\us01\/_0260_ ), .B(\us01\/_0325_ ), .X(\us01\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_0948_ ( .A(\us01\/_0128_ ), .B(\us01\/_0130_ ), .Y(\us01\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_0949_ ( .A(\us01\/_0127_ ), .B(\us01\/_0132_ ), .Y(\us01\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us01/_0950_ ( .A(\us01\/_0434_ ), .X(\us01\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_0951_ ( .A(\us01\/_0134_ ), .B(\us01\/_0128_ ), .Y(\us01\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us01/_0952_ ( .A(\us01\/_0126_ ), .B(\us01\/_0133_ ), .C_N(\us01\/_0135_ ), .Y(\us01\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us01/_0953_ ( .A(\us01\/_0026_ ), .B(\us01\/_0123_ ), .X(\us01\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0955_ ( .A(\us01\/_0137_ ), .X(\us01\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_0956_ ( .A1(\us01\/_0110_ ), .A2(\us01\/_0293_ ), .A3(\us01\/_0280_ ), .B1(\us01\/_0139_ ), .Y(\us01\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0957_ ( .A(\us01\/_0096_ ), .B(\us01\/_0730_ ), .X(\us01\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0959_ ( .A(\us01\/_0142_ ), .X(\us01\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_0960_ ( .A1(\us01\/_0020_ ), .A2(\us01\/_0144_ ), .A3(\us01\/_0017_ ), .B1(\us01\/_0139_ ), .Y(\us01\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \us01/_0961_ ( .A(\sa01\[2\] ), .B(\us01\/_0050_ ), .C_N(\sa01\[3\] ), .Y(\us01\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0962_ ( .A(\us01\/_0128_ ), .X(\us01\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_0963_ ( .A1(\us01\/_0146_ ), .A2(\us01\/_0030_ ), .A3(\us01\/_0640_ ), .B1(\us01\/_0147_ ), .Y(\us01\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us01/_0964_ ( .A(\us01\/_0136_ ), .B(\us01\/_0141_ ), .C(\us01\/_0145_ ), .D(\us01\/_0148_ ), .X(\us01\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0965_ ( .A(\us01\/_0123_ ), .B(\us01\/_0151_ ), .X(\us01\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0967_ ( .A(\us01\/_0150_ ), .X(\us01\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \us01/_0968_ ( .A(\us01\/_0150_ ), .B(\us01\/_0062_ ), .X(\us01\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_0969_ ( .A(\us01\/_0079_ ), .B(\us01\/_0150_ ), .Y(\us01\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us01/_0970_ ( .A(\us01\/_0150_ ), .B(\us01\/_0412_ ), .C(\us01\/_0249_ ), .Y(\us01\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_0971_ ( .A(\us01\/_0155_ ), .B(\us01\/_0156_ ), .Y(\us01\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_0972_ ( .A1(\us01\/_0153_ ), .A2(\us01\/_0134_ ), .B1(\us01\/_0154_ ), .C1(\us01\/_0157_ ), .Y(\us01\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0973_ ( .A(\us01\/_0467_ ), .B(\us01\/_0123_ ), .X(\us01\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_0975_ ( .A(\us01\/_0159_ ), .X(\us01\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us01/_0976_ ( .A_N(\us01\/_0119_ ), .B(\us01\/_0161_ ), .X(\us01\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us01/_0977_ ( .A(\us01\/_0163_ ), .Y(\us01\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_0978_ ( .A1(\us01\/_0146_ ), .A2(\us01\/_0575_ ), .A3(\us01\/_0608_ ), .B1(\us01\/_0153_ ), .Y(\us01\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_0979_ ( .A1(\us01\/_0062_ ), .A2(\us01\/_0280_ ), .A3(\us01\/_0134_ ), .B1(\us01\/_0161_ ), .Y(\us01\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us01/_0980_ ( .A(\us01\/_0158_ ), .B(\us01\/_0164_ ), .C(\us01\/_0165_ ), .D(\us01\/_0166_ ), .X(\us01\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us01/_0981_ ( .A(\us01\/_0097_ ), .B(\us01\/_0122_ ), .C(\us01\/_0149_ ), .D(\us01\/_0167_ ), .X(\us01\/_0168_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0982_ ( .A(\us01\/_0662_ ), .B(\us01\/_0150_ ), .X(\us01\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_0983_ ( .A(\us01\/_0154_ ), .B(\us01\/_0169_ ), .Y(\us01\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us01/_0984_ ( .A(\us01\/_0123_ ), .B(\us01\/_0151_ ), .C(\us01\/_0038_ ), .X(\us01\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0985_ ( .A(\us01\/_0170_ ), .B(\us01\/_0171_ ), .X(\us01\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \us01/_0986_ ( .A(\us01\/_0172_ ), .Y(\us01\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \us01/_0987_ ( .A(\us01\/_0067_ ), .B(\us01\/_0168_ ), .C(\us01\/_0174_ ), .Y(\us01\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us01/_0988_ ( .A(\sa01\[1\] ), .B(\sa01\[0\] ), .Y(\us01\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us01/_0989_ ( .A(\us01\/_0175_ ), .B(\us01\/_0358_ ), .X(\us01\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0990_ ( .A(\us01\/_0176_ ), .B(\us01\/_0478_ ), .X(\us01\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_0991_ ( .A(\us01\/_0280_ ), .B(\us01\/_0113_ ), .Y(\us01\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0992_ ( .A(\us01\/_0111_ ), .B(\us01\/_0062_ ), .X(\us01\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0993_ ( .A(\us01\/_0111_ ), .B(\us01\/_0662_ ), .X(\us01\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_0994_ ( .A(\us01\/_0179_ ), .B(\us01\/_0180_ ), .Y(\us01\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0995_ ( .A(\us01\/_0054_ ), .B(\us01\/_0058_ ), .X(\us01\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us01/_0996_ ( .A(\us01\/_0182_ ), .Y(\us01\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us01/_0997_ ( .A_N(\us01\/_0177_ ), .B(\us01\/_0178_ ), .C(\us01\/_0181_ ), .D(\us01\/_0184_ ), .X(\us01\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0998_ ( .A(\us01\/_0098_ ), .B(\us01\/_0741_ ), .X(\us01\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us01/_0999_ ( .A(\us01\/_0047_ ), .B(\us01\/_0098_ ), .X(\us01\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us01/_1000_ ( .A(\us01\/_0186_ ), .B(\us01\/_0187_ ), .X(\us01\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1001_ ( .A(\us01\/_0188_ ), .Y(\us01\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1002_ ( .A(\us01\/_0738_ ), .B(\us01\/_0735_ ), .X(\us01\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1003_ ( .A(\us01\/_0271_ ), .B(\us01\/_0736_ ), .X(\us01\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_1004_ ( .A(\us01\/_0190_ ), .B(\us01\/_0191_ ), .Y(\us01\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us01/_1005_ ( .A(\us01\/_0096_ ), .B(\us01\/_0325_ ), .X(\us01\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1006_ ( .A1(\us01\/_0193_ ), .A2(\us01\/_0176_ ), .B1(\us01\/_0043_ ), .Y(\us01\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1007_ ( .A(\us01\/_0185_ ), .B(\us01\/_0189_ ), .C(\us01\/_0192_ ), .D(\us01\/_0195_ ), .X(\us01\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us01/_1008_ ( .A_N(\sa01\[3\] ), .B(\us01\/_0734_ ), .C(\sa01\[2\] ), .X(\us01\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1009_ ( .A(\us01\/_0137_ ), .B(\us01\/_0197_ ), .X(\us01\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_1010_ ( .A(\us01\/_0198_ ), .B(\us01\/_0040_ ), .Y(\us01\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1011_ ( .A(\us01\/_0293_ ), .B(\us01\/_0137_ ), .X(\us01\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1012_ ( .A(\us01\/_0200_ ), .Y(\us01\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1013_ ( .A(\us01\/_0137_ ), .B(\us01\/_0110_ ), .Y(\us01\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1014_ ( .A(\us01\/_0139_ ), .B(\us01\/_0020_ ), .Y(\us01\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1015_ ( .A(\us01\/_0199_ ), .B(\us01\/_0201_ ), .C(\us01\/_0202_ ), .D(\us01\/_0203_ ), .X(\us01\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us01/_1016_ ( .A1(\us01\/_0532_ ), .A2(\us01\/_0109_ ), .B1(\us01\/_0102_ ), .C1(\us01\/_0727_ ), .X(\us01\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1017_ ( .A(\us01\/_0022_ ), .B(\us01\/_0078_ ), .Y(\us01\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1018_ ( .A(\us01\/_0078_ ), .B(\us01\/_0142_ ), .Y(\us01\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1019_ ( .A(\us01\/_0207_ ), .B(\us01\/_0208_ ), .Y(\us01\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1020_ ( .A1(\us01\/_0094_ ), .A2(\us01\/_0176_ ), .B1(\us01\/_0206_ ), .C1(\us01\/_0209_ ), .Y(\us01\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1021_ ( .A(\us01\/_0662_ ), .B(\us01\/_0070_ ), .X(\us01\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us01/_1022_ ( .A(\us01\/_0731_ ), .B(\us01\/_0123_ ), .C(\us01\/_0749_ ), .Y(\us01\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us01/_1023_ ( .A(\us01\/_0731_ ), .B(\us01\/_0467_ ), .C(\us01\/_0069_ ), .Y(\us01\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us01/_1024_ ( .A_N(\us01\/_0211_ ), .B(\us01\/_0127_ ), .C(\us01\/_0212_ ), .D(\us01\/_0213_ ), .X(\us01\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1025_ ( .A(\us01\/_0137_ ), .Y(\us01\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1026_ ( .A(\us01\/_0128_ ), .B(\us01\/_0035_ ), .Y(\us01\/_0217_ ) );
sky130_fd_sc_hd__buf_2 \us01/_1027_ ( .A(\us01\/_0478_ ), .X(\us01\/_0218_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1028_ ( .A1(\us01\/_0159_ ), .A2(\us01\/_0746_ ), .B1(\us01\/_0434_ ), .B2(\us01\/_0218_ ), .Y(\us01\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us01/_1029_ ( .A1(\us01\/_0116_ ), .A2(\us01\/_0215_ ), .B1(\us01\/_0217_ ), .C1(\us01\/_0219_ ), .X(\us01\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1030_ ( .A(\us01\/_0113_ ), .B(\us01\/_0746_ ), .X(\us01\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us01/_1031_ ( .A1(\us01\/_0098_ ), .A2(\us01\/_0746_ ), .B1(\us01\/_0434_ ), .B2(\us01\/_0750_ ), .X(\us01\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1032_ ( .A1(\us01\/_0047_ ), .A2(\us01\/_0113_ ), .B1(\us01\/_0221_ ), .C1(\us01\/_0222_ ), .Y(\us01\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us01/_1033_ ( .A1(\us01\/_0129_ ), .A2(\us01\/_0162_ ), .B1(\us01\/_0271_ ), .B2(\us01\/_0705_ ), .X(\us01\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1034_ ( .A1(\us01\/_0093_ ), .A2(\us01\/_0738_ ), .B1(\us01\/_0081_ ), .C1(\us01\/_0224_ ), .Y(\us01\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1035_ ( .A(\us01\/_0214_ ), .B(\us01\/_0220_ ), .C(\us01\/_0223_ ), .D(\us01\/_0225_ ), .X(\us01\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1036_ ( .A(\us01\/_0196_ ), .B(\us01\/_0204_ ), .C(\us01\/_0210_ ), .D(\us01\/_0226_ ), .X(\us01\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1037_ ( .A(\us01\/_0111_ ), .B(\us01\/_0554_ ), .X(\us01\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1038_ ( .A(\us01\/_0229_ ), .Y(\us01\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1039_ ( .A(\us01\/_0111_ ), .B(\us01\/_0129_ ), .Y(\us01\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1040_ ( .A(\us01\/_0017_ ), .B(\us01\/_0738_ ), .Y(\us01\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1041_ ( .A(\us01\/_0030_ ), .B(\us01\/_0304_ ), .Y(\us01\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1042_ ( .A(\us01\/_0230_ ), .B(\us01\/_0231_ ), .C(\us01\/_0232_ ), .D(\us01\/_0233_ ), .X(\us01\/_0234_ ) );
sky130_fd_sc_hd__and2_1 \us01/_1043_ ( .A(\us01\/_0047_ ), .B(\us01\/_0478_ ), .X(\us01\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1044_ ( .A1(\us01\/_0129_ ), .A2(\us01\/_0554_ ), .B1(\us01\/_0137_ ), .Y(\us01\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us01/_1045_ ( .A(\us01\/_0235_ ), .B(\us01\/_0049_ ), .C_N(\us01\/_0236_ ), .Y(\us01\/_0237_ ) );
sky130_fd_sc_hd__and2_1 \us01/_1046_ ( .A(\us01\/_0047_ ), .B(\us01\/_0077_ ), .X(\us01\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1047_ ( .A(\us01\/_0070_ ), .B(\us01\/_0035_ ), .X(\us01\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us01/_1048_ ( .A1(\us01\/_0047_ ), .A2(\us01\/_0736_ ), .B1(\us01\/_0022_ ), .B2(\us01\/_0099_ ), .X(\us01\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us01/_1049_ ( .A(\us01\/_0239_ ), .B(\us01\/_0240_ ), .C(\us01\/_0241_ ), .Y(\us01\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1050_ ( .A(\us01\/_0554_ ), .B(\us01\/_0072_ ), .X(\us01\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us01/_1051_ ( .A1(\us01\/_0142_ ), .A2(\us01\/_0137_ ), .B1(\us01\/_0159_ ), .B2(\us01\/_0082_ ), .X(\us01\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1052_ ( .A1(\us01\/_0608_ ), .A2(\us01\/_0072_ ), .B1(\us01\/_0243_ ), .C1(\us01\/_0244_ ), .Y(\us01\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1053_ ( .A(\us01\/_0234_ ), .B(\us01\/_0237_ ), .C(\us01\/_0242_ ), .D(\us01\/_0245_ ), .X(\us01\/_0246_ ) );
sky130_fd_sc_hd__o21a_1 \us01/_1055_ ( .A1(\us01\/_0554_ ), .A2(\us01\/_0586_ ), .B1(\us01\/_0029_ ), .X(\us01\/_0248_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1056_ ( .A(\us01\/_0082_ ), .B(\us01\/_0478_ ), .X(\us01\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_1057_ ( .A(\us01\/_0079_ ), .X(\us01\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1058_ ( .A(\us01\/_0251_ ), .B(\us01\/_0478_ ), .X(\us01\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_1059_ ( .A(\us01\/_0250_ ), .B(\us01\/_0252_ ), .Y(\us01\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1060_ ( .A(\us01\/_0016_ ), .B(\us01\/_0064_ ), .Y(\us01\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_1061_ ( .A(\us01\/_0304_ ), .X(\us01\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1062_ ( .A(\us01\/_0255_ ), .B(\us01\/_0640_ ), .Y(\us01\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us01/_1063_ ( .A_N(\us01\/_0248_ ), .B(\us01\/_0253_ ), .C(\us01\/_0254_ ), .D(\us01\/_0256_ ), .X(\us01\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1064_ ( .A(\us01\/_0099_ ), .B(\us01\/_0110_ ), .X(\us01\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us01/_1065_ ( .A1(\us01\/_0161_ ), .A2(\us01\/_0130_ ), .B1(\us01\/_0258_ ), .Y(\us01\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1066_ ( .A(\us01\/_0194_ ), .B(\sa01\[1\] ), .X(\us01\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1068_ ( .A(\us01\/_0261_ ), .B(\us01\/_0153_ ), .Y(\us01\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us01/_1069_ ( .A_N(\us01\/_0154_ ), .B(\us01\/_0259_ ), .C(\us01\/_0263_ ), .X(\us01\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1070_ ( .A(\us01\/_0246_ ), .B(\us01\/_0174_ ), .C(\us01\/_0257_ ), .D(\us01\/_0264_ ), .X(\us01\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us01/_1071_ ( .A1(\us01\/_0261_ ), .A2(\us01\/_0554_ ), .B1(\us01\/_0159_ ), .X(\us01\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1072_ ( .A(\us01\/_0746_ ), .B(\us01\/_0150_ ), .Y(\us01\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1073_ ( .A(\us01\/_0175_ ), .Y(\us01\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us01/_1074_ ( .A(\us01\/_0412_ ), .B(\us01\/_0123_ ), .C(\us01\/_0151_ ), .X(\us01\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1075_ ( .A(\us01\/_0268_ ), .B(\us01\/_0269_ ), .Y(\us01\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us01/_1076_ ( .A_N(\us01\/_0266_ ), .B(\us01\/_0267_ ), .C(\us01\/_0270_ ), .X(\us01\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1077_ ( .A(\us01\/_0554_ ), .B(\us01\/_0150_ ), .X(\us01\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1078_ ( .A(\us01\/_0273_ ), .Y(\us01\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1079_ ( .A1(\us01\/_0734_ ), .A2(\us01\/_0325_ ), .B1(\us01\/_0380_ ), .Y(\us01\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1080_ ( .A(\us01\/_0275_ ), .Y(\us01\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1081_ ( .A(\us01\/_0276_ ), .B(\us01\/_0153_ ), .Y(\us01\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us01/_1082_ ( .A(\us01\/_0272_ ), .B(\us01\/_0274_ ), .C(\us01\/_0277_ ), .X(\us01\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_1083_ ( .A(\us01\/_0035_ ), .X(\us01\/_0279_ ) );
sky130_fd_sc_hd__buf_2 \us01/_1084_ ( .A(\us01\/_0082_ ), .X(\us01\/_0280_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1085_ ( .A1(\us01\/_0218_ ), .A2(\us01\/_0279_ ), .B1(\us01\/_0280_ ), .B2(\us01\/_0060_ ), .Y(\us01\/_0281_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1086_ ( .A1(\us01\/_0251_ ), .A2(\us01\/_0434_ ), .B1(\us01\/_0304_ ), .Y(\us01\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1087_ ( .A(\us01\/_0091_ ), .B(\us01\/_0292_ ), .Y(\us01\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1088_ ( .A1(\us01\/_0118_ ), .A2(\us01\/_0050_ ), .B1(\us01\/_0038_ ), .C1(\us01\/_0255_ ), .Y(\us01\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1089_ ( .A(\us01\/_0281_ ), .B(\us01\/_0283_ ), .C(\us01\/_0284_ ), .D(\us01\/_0285_ ), .X(\us01\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1090_ ( .A(\us01\/_0082_ ), .B(\us01\/_0027_ ), .X(\us01\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1091_ ( .A(\us01\/_0129_ ), .B(\us01\/_0027_ ), .X(\us01\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_1092_ ( .A(\us01\/_0287_ ), .B(\us01\/_0288_ ), .Y(\us01\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1093_ ( .A1(\us01\/_0752_ ), .A2(\us01\/_0683_ ), .B1(\us01\/_0093_ ), .B2(\us01\/_0029_ ), .Y(\us01\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1094_ ( .A1(\us01\/_0092_ ), .A2(\us01\/_0575_ ), .B1(\us01\/_0292_ ), .Y(\us01\/_0291_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_1095_ ( .A(\us01\/_0054_ ), .X(\us01\/_0292_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1096_ ( .A1(\us01\/_0218_ ), .A2(\us01\/_0662_ ), .B1(\us01\/_0280_ ), .B2(\us01\/_0292_ ), .Y(\us01\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1097_ ( .A(\us01\/_0289_ ), .B(\us01\/_0290_ ), .C(\us01\/_0291_ ), .D(\us01\/_0294_ ), .X(\us01\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1098_ ( .A(\us01\/_0750_ ), .B(\us01\/_0193_ ), .X(\us01\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1099_ ( .A(\us01\/_0705_ ), .B(\us01\/_0380_ ), .X(\us01\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1100_ ( .A(\us01\/_0752_ ), .B(\us01\/_0129_ ), .Y(\us01\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us01/_1101_ ( .A(\us01\/_0296_ ), .B(\us01\/_0297_ ), .C_N(\us01\/_0298_ ), .Y(\us01\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1102_ ( .A(\us01\/_0089_ ), .B(\us01\/_0532_ ), .Y(\us01\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1103_ ( .A(\sa01\[2\] ), .Y(\us01\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \us01/_1104_ ( .A(\us01\/_0301_ ), .B(\sa01\[3\] ), .C(\us01\/_0118_ ), .Y(\us01\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1105_ ( .A(\us01\/_0072_ ), .B(\us01\/_0302_ ), .X(\us01\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1106_ ( .A(\us01\/_0303_ ), .Y(\us01\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1107_ ( .A(\us01\/_0147_ ), .B(\us01\/_0302_ ), .Y(\us01\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1108_ ( .A(\us01\/_0299_ ), .B(\us01\/_0300_ ), .C(\us01\/_0305_ ), .D(\us01\/_0306_ ), .X(\us01\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1109_ ( .A(\us01\/_0278_ ), .B(\us01\/_0286_ ), .C(\us01\/_0295_ ), .D(\us01\/_0307_ ), .X(\us01\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us01/_1110_ ( .A(\us01\/_0228_ ), .B(\us01\/_0265_ ), .C(\us01\/_0308_ ), .Y(\us01\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1111_ ( .A(\us01\/_0235_ ), .Y(\us01\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1112_ ( .A(\us01\/_0478_ ), .B(\us01\/_0640_ ), .X(\us01\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1113_ ( .A(\us01\/_0310_ ), .Y(\us01\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1114_ ( .A(\us01\/_0022_ ), .B(\us01\/_0218_ ), .Y(\us01\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1115_ ( .A(\us01\/_0218_ ), .B(\us01\/_0030_ ), .Y(\us01\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1116_ ( .A(\us01\/_0309_ ), .B(\us01\/_0311_ ), .C(\us01\/_0312_ ), .D(\us01\/_0313_ ), .X(\us01\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1117_ ( .A(\us01\/_0218_ ), .B(\us01\/_0064_ ), .Y(\us01\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1118_ ( .A(\us01\/_0218_ ), .B(\us01\/_0683_ ), .Y(\us01\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1119_ ( .A(\us01\/_0315_ ), .B(\us01\/_0316_ ), .C(\us01\/_0317_ ), .D(\us01\/_0253_ ), .X(\us01\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1120_ ( .A(\us01\/_0047_ ), .B(\us01\/_0304_ ), .Y(\us01\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1121_ ( .A(\us01\/_0586_ ), .B(\us01\/_0162_ ), .Y(\us01\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1122_ ( .A(\us01\/_0319_ ), .B(\us01\/_0320_ ), .Y(\us01\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_1123_ ( .A(\us01\/_0321_ ), .B(\us01\/_0238_ ), .Y(\us01\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1124_ ( .A(\us01\/_0304_ ), .B(\us01\/_0062_ ), .Y(\us01\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_1125_ ( .A(\us01\/_0251_ ), .X(\us01\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1126_ ( .A1(\us01\/_0324_ ), .A2(\us01\/_0280_ ), .B1(\us01\/_0255_ ), .Y(\us01\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1127_ ( .A1(\us01\/_0050_ ), .A2(\us01\/_0205_ ), .B1(\us01\/_0109_ ), .C1(\us01\/_0255_ ), .Y(\us01\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1128_ ( .A(\us01\/_0322_ ), .B(\us01\/_0323_ ), .C(\us01\/_0326_ ), .D(\us01\/_0327_ ), .X(\us01\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1129_ ( .A1(\us01\/_0733_ ), .A2(\us01\/_0279_ ), .A3(\us01\/_0058_ ), .B1(\us01\/_0292_ ), .Y(\us01\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_1130_ ( .A(\us01\/_0047_ ), .X(\us01\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1131_ ( .A(\us01\/_0330_ ), .B(\us01\/_0292_ ), .Y(\us01\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1132_ ( .A(\us01\/_0054_ ), .B(\us01\/_0045_ ), .Y(\us01\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1133_ ( .A(\us01\/_0329_ ), .B(\us01\/_0331_ ), .C(\us01\/_0284_ ), .D(\us01\/_0332_ ), .X(\us01\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us01/_1134_ ( .A1(\us01\/_0249_ ), .A2(\us01\/_0205_ ), .B1(\us01\/_0532_ ), .C1(\us01\/_0060_ ), .X(\us01\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1135_ ( .A(\us01\/_0280_ ), .B(\us01\/_0060_ ), .Y(\us01\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1136_ ( .A(\us01\/_0324_ ), .B(\us01\/_0060_ ), .Y(\us01\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1137_ ( .A(\us01\/_0335_ ), .B(\us01\/_0337_ ), .Y(\us01\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1138_ ( .A1(\us01\/_0276_ ), .A2(\us01\/_0060_ ), .B1(\us01\/_0334_ ), .C1(\us01\/_0338_ ), .Y(\us01\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1139_ ( .A(\us01\/_0318_ ), .B(\us01\/_0328_ ), .C(\us01\/_0333_ ), .D(\us01\/_0339_ ), .X(\us01\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us01/_1140_ ( .A1(\us01\/_0746_ ), .A2(\us01\/_0134_ ), .B1(\us01\/_0128_ ), .X(\us01\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us01/_1141_ ( .A_N(\us01\/_0086_ ), .B(\us01\/_0128_ ), .X(\us01\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1142_ ( .A(\us01\/_0079_ ), .B(\us01\/_0124_ ), .X(\us01\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_1143_ ( .A(\us01\/_0126_ ), .B(\us01\/_0343_ ), .Y(\us01\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us01/_1144_ ( .A(\us01\/_0341_ ), .B(\us01\/_0342_ ), .C_N(\us01\/_0344_ ), .Y(\us01\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1146_ ( .A1(\us01\/_0193_ ), .A2(\us01\/_0092_ ), .A3(\us01\/_0330_ ), .B1(\us01\/_0147_ ), .Y(\us01\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1147_ ( .A1(\us01\/_0130_ ), .A2(\us01\/_0280_ ), .A3(\us01\/_0134_ ), .B1(\us01\/_0139_ ), .Y(\us01\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1148_ ( .A1(\us01\/_0144_ ), .A2(\us01\/_0608_ ), .A3(\us01\/_0092_ ), .B1(\us01\/_0139_ ), .Y(\us01\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1149_ ( .A(\us01\/_0345_ ), .B(\us01\/_0348_ ), .C(\us01\/_0349_ ), .D(\us01\/_0350_ ), .X(\us01\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us01/_1150_ ( .A(\us01\/_0150_ ), .B(\us01\/_0194_ ), .C(\us01\/_0249_ ), .X(\us01\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us01/_1151_ ( .A(\us01\/_0277_ ), .SLEEP(\us01\/_0352_ ), .X(\us01\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us01/_1152_ ( .A1(\us01\/_0268_ ), .A2(\us01\/_0171_ ), .B1(\us01\/_0157_ ), .Y(\us01\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us01/_1153_ ( .A(\us01\/_0161_ ), .X(\us01\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1154_ ( .A1(\us01\/_0279_ ), .A2(\us01\/_0280_ ), .B1(\us01\/_0355_ ), .Y(\us01\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1155_ ( .A1(\us01\/_0020_ ), .A2(\us01\/_0193_ ), .A3(\us01\/_0091_ ), .B1(\us01\/_0355_ ), .Y(\us01\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1156_ ( .A(\us01\/_0353_ ), .B(\us01\/_0354_ ), .C(\us01\/_0356_ ), .D(\us01\/_0357_ ), .X(\us01\/_0359_ ) );
sky130_fd_sc_hd__and2_1 \us01/_1157_ ( .A(\us01\/_0111_ ), .B(\us01\/_0586_ ), .X(\us01\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1158_ ( .A(\us01\/_0360_ ), .Y(\us01\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us01/_1159_ ( .A1(\us01\/_0119_ ), .A2(\us01\/_0120_ ), .B1(\us01\/_0230_ ), .C1(\us01\/_0361_ ), .X(\us01\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1160_ ( .A1(\us01\/_0662_ ), .A2(\us01\/_0251_ ), .A3(\us01\/_0134_ ), .B1(\us01\/_0114_ ), .Y(\us01\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1162_ ( .A1(\us01\/_0035_ ), .A2(\us01\/_0251_ ), .A3(\us01\/_0134_ ), .B1(\us01\/_0099_ ), .Y(\us01\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1163_ ( .A1(\us01\/_0193_ ), .A2(\us01\/_0608_ ), .B1(\us01\/_0099_ ), .Y(\us01\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1164_ ( .A(\us01\/_0362_ ), .B(\us01\/_0363_ ), .C(\us01\/_0365_ ), .D(\us01\/_0366_ ), .X(\us01\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1165_ ( .A1(\us01\/_0575_ ), .A2(\us01\/_0092_ ), .A3(\us01\/_0330_ ), .B1(\us01\/_0089_ ), .Y(\us01\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1166_ ( .A1(\us01\/_0586_ ), .A2(\us01\/_0017_ ), .A3(\us01\/_0330_ ), .B1(\us01\/_0094_ ), .Y(\us01\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \us01/_1167_ ( .A1(\us01\/_0293_ ), .A2(\us01\/_0134_ ), .B1(\us01\/_0089_ ), .Y(\us01\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1168_ ( .A1(\us01\/_0279_ ), .A2(\us01\/_0134_ ), .B1(\us01\/_0094_ ), .Y(\us01\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1169_ ( .A(\us01\/_0368_ ), .B(\us01\/_0370_ ), .C(\us01\/_0371_ ), .D(\us01\/_0372_ ), .X(\us01\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1170_ ( .A(\us01\/_0351_ ), .B(\us01\/_0359_ ), .C(\us01\/_0367_ ), .D(\us01\/_0373_ ), .X(\us01\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1171_ ( .A1(\us01\/_0102_ ), .A2(\us01\/_0347_ ), .B1(\us01\/_0109_ ), .C1(\us01\/_0029_ ), .Y(\us01\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1172_ ( .A1(\us01\/_0102_ ), .A2(\us01\/_0347_ ), .B1(\us01\/_0532_ ), .C1(\us01\/_0029_ ), .Y(\us01\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1173_ ( .A1(\us01\/_0050_ ), .A2(\us01\/_0249_ ), .B1(\us01\/_0380_ ), .C1(\us01\/_0029_ ), .Y(\us01\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1174_ ( .A(\us01\/_0041_ ), .B(\us01\/_0375_ ), .C(\us01\/_0376_ ), .D(\us01\/_0377_ ), .X(\us01\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1175_ ( .A(\us01\/_0047_ ), .B(\us01\/_0750_ ), .X(\us01\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1176_ ( .A(\us01\/_0379_ ), .Y(\us01\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1177_ ( .A(\us01\/_0016_ ), .B(\us01\/_0608_ ), .Y(\us01\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1178_ ( .A(\us01\/_0752_ ), .B(\us01\/_0554_ ), .Y(\us01\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1179_ ( .A1(\sa01\[1\] ), .A2(\us01\/_0734_ ), .B1(\us01\/_0109_ ), .C1(\us01\/_0016_ ), .Y(\us01\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1180_ ( .A(\us01\/_0381_ ), .B(\us01\/_0382_ ), .C(\us01\/_0383_ ), .D(\us01\/_0384_ ), .X(\us01\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us01/_1181_ ( .A(\us01\/_0086_ ), .B_N(\us01\/_0736_ ), .X(\us01\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1182_ ( .A1(\us01\/_0748_ ), .A2(\us01\/_0134_ ), .B1(\us01\/_0739_ ), .Y(\us01\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1183_ ( .A1(\us01\/_0118_ ), .A2(\us01\/_0249_ ), .B1(\us01\/_0109_ ), .C1(\us01\/_0739_ ), .Y(\us01\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1184_ ( .A1(\us01\/_0102_ ), .A2(\us01\/_0301_ ), .B1(\sa01\[3\] ), .C1(\us01\/_0739_ ), .Y(\us01\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1185_ ( .A(\us01\/_0386_ ), .B(\us01\/_0387_ ), .C(\us01\/_0388_ ), .D(\us01\/_0389_ ), .X(\us01\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1186_ ( .A(\us01\/_0020_ ), .Y(\us01\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1187_ ( .A(\us01\/_0727_ ), .Y(\us01\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1188_ ( .A(\us01\/_0727_ ), .B(\us01\/_0064_ ), .Y(\us01\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1189_ ( .A1(\us01\/_0102_ ), .A2(\us01\/_0734_ ), .B1(\us01\/_0532_ ), .C1(\us01\/_0727_ ), .Y(\us01\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us01/_1190_ ( .A1(\us01\/_0392_ ), .A2(\us01\/_0393_ ), .B1(\us01\/_0394_ ), .C1(\us01\/_0395_ ), .X(\us01\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1191_ ( .A(\us01\/_0378_ ), .B(\us01\/_0385_ ), .C(\us01\/_0390_ ), .D(\us01\/_0396_ ), .X(\us01\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us01/_1192_ ( .A(\us01\/_0340_ ), .B(\us01\/_0374_ ), .C(\us01\/_0397_ ), .Y(\us01\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1193_ ( .A(\us01\/_0077_ ), .B(\us01\/_0129_ ), .X(\us01\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_1194_ ( .A(\us01\/_0398_ ), .B(\us01\/_0239_ ), .Y(\us01\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1195_ ( .A(\us01\/_0022_ ), .B(\us01\/_0111_ ), .X(\us01\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us01/_1196_ ( .A_N(\us01\/_0400_ ), .B(\us01\/_0231_ ), .Y(\us01\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us01/_1197_ ( .A(\us01\/_0399_ ), .SLEEP(\us01\/_0402_ ), .X(\us01\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_1198_ ( .A(\us01\/_0746_ ), .B(\us01\/_0251_ ), .Y(\us01\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us01/_1199_ ( .A_N(\us01\/_0404_ ), .B(\us01\/_0752_ ), .Y(\us01\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us01/_1200_ ( .A(\us01\/_0467_ ), .B(\us01\/_0194_ ), .C(\us01\/_0694_ ), .X(\us01\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us01/_1201_ ( .A_N(\us01\/_0175_ ), .B(\us01\/_0406_ ), .X(\us01\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1202_ ( .A(\us01\/_0407_ ), .Y(\us01\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1203_ ( .A1(\us01\/_0094_ ), .A2(\us01\/_0197_ ), .B1(\us01\/_0114_ ), .B2(\us01\/_0640_ ), .Y(\us01\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1204_ ( .A(\us01\/_0403_ ), .B(\us01\/_0405_ ), .C(\us01\/_0408_ ), .D(\us01\/_0409_ ), .X(\us01\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1205_ ( .A(\us01\/_0030_ ), .B(\us01\/_0150_ ), .Y(\us01\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us01/_1206_ ( .A_N(\us01\/_0169_ ), .B(\us01\/_0289_ ), .C(\us01\/_0411_ ), .X(\us01\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us01/_1207_ ( .A1(\us01\/_0467_ ), .A2(\us01\/_0151_ ), .B1(\us01\/_0140_ ), .C1(\us01\/_0129_ ), .X(\us01\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1208_ ( .A1(\us01\/_0608_ ), .A2(\us01\/_0099_ ), .B1(\us01\/_0037_ ), .C1(\us01\/_0414_ ), .Y(\us01\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1209_ ( .A(\us01\/_0738_ ), .Y(\us01\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1210_ ( .A(\us01\/_0586_ ), .B(\us01\/_0736_ ), .Y(\us01\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1211_ ( .A1(\us01\/_0194_ ), .A2(\us01\/_0038_ ), .B1(\us01\/_0118_ ), .C1(\us01\/_0153_ ), .Y(\us01\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us01/_1212_ ( .A1(\us01\/_0416_ ), .A2(\us01\/_0117_ ), .B1(\us01\/_0417_ ), .C1(\us01\/_0418_ ), .X(\us01\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1213_ ( .A(\us01\/_0077_ ), .B(\us01\/_0035_ ), .X(\us01\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1214_ ( .A(\us01\/_0662_ ), .B(\us01\/_0124_ ), .Y(\us01\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1215_ ( .A(\us01\/_0030_ ), .B(\us01\/_0137_ ), .Y(\us01\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1216_ ( .A(\us01\/_0072_ ), .B(\us01\/_0731_ ), .Y(\us01\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us01/_1217_ ( .A_N(\us01\/_0420_ ), .B(\us01\/_0421_ ), .C(\us01\/_0422_ ), .D(\us01\/_0424_ ), .X(\us01\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1218_ ( .A(\us01\/_0413_ ), .B(\us01\/_0415_ ), .C(\us01\/_0419_ ), .D(\us01\/_0425_ ), .X(\us01\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us01/_1219_ ( .A(\us01\/_0355_ ), .B(\us01\/_0102_ ), .C(\us01\/_0109_ ), .Y(\us01\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1220_ ( .A(\us01\/_0077_ ), .B(\us01\/_0017_ ), .X(\us01\/_0428_ ) );
sky130_fd_sc_hd__and2_1 \us01/_1221_ ( .A(\us01\/_0077_ ), .B(\us01\/_0554_ ), .X(\us01\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us01/_1222_ ( .A1(\us01\/_0050_ ), .A2(\us01\/_0205_ ), .B1(\us01\/_0380_ ), .C1(\us01\/_0078_ ), .X(\us01\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us01/_1223_ ( .A(\us01\/_0428_ ), .B(\us01\/_0429_ ), .C(\us01\/_0430_ ), .Y(\us01\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us01/_1224_ ( .A_N(\us01\/_0209_ ), .B(\us01\/_0431_ ), .X(\us01\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us01/_1225_ ( .A1(\us01\/_0215_ ), .A2(\us01\/_0404_ ), .B1(\us01\/_0427_ ), .C1(\us01\/_0432_ ), .X(\us01\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1226_ ( .A(\us01\/_0043_ ), .B(\us01\/_0058_ ), .Y(\us01\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1227_ ( .A(\us01\/_0195_ ), .B(\us01\/_0233_ ), .C(\us01\/_0320_ ), .D(\us01\/_0435_ ), .X(\us01\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1228_ ( .A(\us01\/_0261_ ), .B(\us01\/_0738_ ), .Y(\us01\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1229_ ( .A1(\us01\/_0218_ ), .A2(\us01\/_0640_ ), .B1(\us01\/_0261_ ), .B2(\us01\/_0292_ ), .Y(\us01\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1230_ ( .A(\us01\/_0436_ ), .B(\us01\/_0394_ ), .C(\us01\/_0437_ ), .D(\us01\/_0438_ ), .X(\us01\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1231_ ( .A(\us01\/_0410_ ), .B(\us01\/_0426_ ), .C(\us01\/_0433_ ), .D(\us01\/_0439_ ), .X(\us01\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us01/_1232_ ( .A(\us01\/_0135_ ), .SLEEP(\us01\/_0273_ ), .X(\us01\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1233_ ( .A1(\us01\/_0279_ ), .A2(\us01\/_0134_ ), .B1(\us01\/_0099_ ), .Y(\us01\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1234_ ( .A(\us01\/_0441_ ), .B(\us01\/_0164_ ), .C(\us01\/_0270_ ), .D(\us01\/_0442_ ), .X(\us01\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1235_ ( .A(\us01\/_0051_ ), .B(\us01\/_0662_ ), .Y(\us01\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1236_ ( .A(\us01\/_0051_ ), .B(\us01\/_0271_ ), .Y(\us01\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1237_ ( .A(\us01\/_0444_ ), .B(\us01\/_0446_ ), .X(\us01\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1238_ ( .A(\us01\/_0193_ ), .B(\us01\/_0304_ ), .X(\us01\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1239_ ( .A(\us01\/_0448_ ), .Y(\us01\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1240_ ( .A(\us01\/_0162_ ), .B(\us01\/_0130_ ), .X(\us01\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1241_ ( .A(\us01\/_0450_ ), .Y(\us01\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1242_ ( .A1(\us01\/_0129_ ), .A2(\us01\/_0554_ ), .B1(\us01\/_0043_ ), .Y(\us01\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1243_ ( .A(\us01\/_0447_ ), .B(\us01\/_0449_ ), .C(\us01\/_0451_ ), .D(\us01\/_0452_ ), .X(\us01\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1244_ ( .A(\us01\/_0292_ ), .B(\us01\/_0064_ ), .Y(\us01\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us01/_1245_ ( .A_N(\us01\/_0248_ ), .B(\us01\/_0454_ ), .C(\us01\/_0254_ ), .D(\us01\/_0256_ ), .X(\us01\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1246_ ( .A1(\us01\/_0330_ ), .A2(\us01\/_0099_ ), .B1(\us01\/_0134_ ), .B2(\us01\/_0705_ ), .Y(\us01\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1247_ ( .A1(\us01\/_0748_ ), .A2(\us01\/_0738_ ), .B1(\us01\/_0092_ ), .B2(\us01\/_0752_ ), .Y(\us01\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1248_ ( .A1(\us01\/_0072_ ), .A2(\us01\/_0035_ ), .B1(\us01\/_0748_ ), .B2(\us01\/_0292_ ), .Y(\us01\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1249_ ( .A1(\us01\/_0748_ ), .A2(\us01\/_0251_ ), .B1(\us01\/_0029_ ), .Y(\us01\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1250_ ( .A(\us01\/_0457_ ), .B(\us01\/_0458_ ), .C(\us01\/_0459_ ), .D(\us01\/_0460_ ), .X(\us01\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1251_ ( .A(\us01\/_0443_ ), .B(\us01\/_0453_ ), .C(\us01\/_0455_ ), .D(\us01\/_0461_ ), .X(\us01\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1252_ ( .A(\us01\/_0705_ ), .B(\us01\/_0079_ ), .X(\us01\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1253_ ( .A(\us01\/_0586_ ), .B(\us01\/_0124_ ), .Y(\us01\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1254_ ( .A(\us01\/_0218_ ), .B(\us01\/_0746_ ), .Y(\us01\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us01/_1255_ ( .A_N(\us01\/_0463_ ), .B(\us01\/_0464_ ), .C(\us01\/_0465_ ), .X(\us01\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us01/_1256_ ( .A1(\us01\/_0271_ ), .A2(\us01\/_0072_ ), .B1(\us01\/_0142_ ), .B2(\us01\/_0027_ ), .X(\us01\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1257_ ( .A1(\us01\/_0144_ ), .A2(\us01\/_0099_ ), .B1(\us01\/_0360_ ), .C1(\us01\/_0468_ ), .Y(\us01\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us01/_1258_ ( .A1(\us01\/_0662_ ), .A2(\us01\/_0251_ ), .B1(\us01\/_0218_ ), .X(\us01\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1259_ ( .A1(\us01\/_0575_ ), .A2(\us01\/_0292_ ), .B1(\us01\/_0379_ ), .C1(\us01\/_0470_ ), .Y(\us01\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1260_ ( .A(\us01\/_0466_ ), .B(\us01\/_0469_ ), .C(\us01\/_0471_ ), .D(\us01\/_0305_ ), .X(\us01\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us01/_1261_ ( .A1(\us01\/_0029_ ), .A2(\us01\/_0683_ ), .B1(\us01\/_0324_ ), .B2(\us01\/_0292_ ), .X(\us01\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1262_ ( .A(\us01\/_0280_ ), .B(\us01\/_0099_ ), .X(\us01\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us01/_1263_ ( .A1(\us01\/_0092_ ), .A2(\us01\/_0029_ ), .B1(\us01\/_0474_ ), .X(\us01\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us01/_1264_ ( .A(\us01\/_0075_ ), .B(\us01\/_0473_ ), .C(\us01\/_0475_ ), .Y(\us01\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1265_ ( .A1(\us01\/_0279_ ), .A2(\us01\/_0255_ ), .B1(\us01\/_0280_ ), .B2(\us01\/_0060_ ), .Y(\us01\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1266_ ( .A1(\us01\/_0093_ ), .A2(\us01\/_0292_ ), .B1(\us01\/_0134_ ), .B2(\us01\/_0114_ ), .Y(\us01\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1267_ ( .A1(\us01\/_0161_ ), .A2(\us01\/_0030_ ), .B1(\us01\/_0324_ ), .B2(\us01\/_0147_ ), .Y(\us01\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1268_ ( .A1(\us01\/_0054_ ), .A2(\us01\/_0731_ ), .B1(\us01\/_0748_ ), .B2(\us01\/_0304_ ), .Y(\us01\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1269_ ( .A(\us01\/_0477_ ), .B(\us01\/_0479_ ), .C(\us01\/_0480_ ), .D(\us01\/_0481_ ), .X(\us01\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1270_ ( .A(\us01\/_0161_ ), .B(\us01\/_0064_ ), .Y(\us01\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us01/_1271_ ( .A(\us01\/_0731_ ), .B(\us01\/_0123_ ), .C(\us01\/_0467_ ), .Y(\us01\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1272_ ( .A(\us01\/_0483_ ), .B(\us01\/_0484_ ), .Y(\us01\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1273_ ( .A(\us01\/_0297_ ), .Y(\us01\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us01/_1274_ ( .A_N(\us01\/_0485_ ), .B(\us01\/_0181_ ), .C(\us01\/_0486_ ), .D(\us01\/_0386_ ), .X(\us01\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1275_ ( .A(\us01\/_0472_ ), .B(\us01\/_0476_ ), .C(\us01\/_0482_ ), .D(\us01\/_0487_ ), .X(\us01\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \us01/_1276_ ( .A(\us01\/_0440_ ), .B(\us01\/_0462_ ), .C(\us01\/_0488_ ), .Y(\us01\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1277_ ( .A(\us01\/_0403_ ), .B(\us01\/_0230_ ), .C(\us01\/_0451_ ), .D(\us01\/_0361_ ), .X(\us01\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1278_ ( .A1(\us01\/_0118_ ), .A2(\us01\/_0050_ ), .B1(\us01\/_0109_ ), .C1(\us01\/_0139_ ), .Y(\us01\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1279_ ( .A(\us01\/_0447_ ), .B(\us01\/_0437_ ), .C(\us01\/_0491_ ), .D(\us01\/_0427_ ), .X(\us01\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1280_ ( .A1(\us01\/_0280_ ), .A2(\us01\/_0255_ ), .B1(\us01\/_0608_ ), .B2(\us01\/_0029_ ), .Y(\us01\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1281_ ( .A1(\us01\/_0144_ ), .A2(\us01\/_0147_ ), .B1(\us01\/_0355_ ), .B2(\us01\/_0093_ ), .Y(\us01\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1282_ ( .A1(\us01\/_0705_ ), .A2(\us01\/_0279_ ), .B1(\us01\/_0330_ ), .B2(\us01\/_0029_ ), .Y(\us01\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1283_ ( .A1(\us01\/_0279_ ), .A2(\us01\/_0280_ ), .B1(\us01\/_0114_ ), .Y(\us01\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1284_ ( .A(\us01\/_0493_ ), .B(\us01\/_0494_ ), .C(\us01\/_0495_ ), .D(\us01\/_0496_ ), .X(\us01\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1285_ ( .A1(\us01\/_0134_ ), .A2(\us01\/_0137_ ), .B1(\us01\/_0355_ ), .B2(\us01\/_0575_ ), .Y(\us01\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1286_ ( .A1(\us01\/_0099_ ), .A2(\us01\/_0733_ ), .B1(\us01\/_0093_ ), .B2(\us01\/_0218_ ), .Y(\us01\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1287_ ( .A(\us01\/_0147_ ), .B(\us01\/_0640_ ), .Y(\us01\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1288_ ( .A1(\us01\/_0153_ ), .A2(\us01\/_0292_ ), .B1(\us01\/_0748_ ), .Y(\us01\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1289_ ( .A(\us01\/_0498_ ), .B(\us01\/_0500_ ), .C(\us01\/_0501_ ), .D(\us01\/_0502_ ), .X(\us01\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1290_ ( .A(\us01\/_0490_ ), .B(\us01\/_0492_ ), .C(\us01\/_0497_ ), .D(\us01\/_0503_ ), .X(\us01\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us01/_1291_ ( .A_N(\us01\/_0275_ ), .B(\us01\/_0705_ ), .X(\us01\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1292_ ( .A(\us01\/_0505_ ), .Y(\us01\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1293_ ( .A(\us01\/_0380_ ), .B(\us01\/_0347_ ), .X(\us01\/_0507_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1294_ ( .A1(\us01\/_0507_ ), .A2(\us01\/_0093_ ), .B1(\us01\/_0292_ ), .Y(\us01\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1295_ ( .A(\us01\/_0322_ ), .B(\us01\/_0277_ ), .C(\us01\/_0506_ ), .D(\us01\/_0508_ ), .X(\us01\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1296_ ( .A(\us01\/_0280_ ), .B(\us01\/_0705_ ), .X(\us01\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1297_ ( .A1(\us01\/_0733_ ), .A2(\us01\/_0114_ ), .B1(\us01\/_0429_ ), .C1(\us01\/_0511_ ), .Y(\us01\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_1298_ ( .A(\us01\/_0019_ ), .B(\us01\/_0024_ ), .Y(\us01\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1299_ ( .A(\us01\/_0512_ ), .B(\us01\/_0513_ ), .C(\us01\/_0742_ ), .D(\us01\/_0306_ ), .X(\us01\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1300_ ( .A1(\us01\/_0532_ ), .A2(\us01\/_0089_ ), .B1(\us01\/_0154_ ), .C1(\us01\/_0169_ ), .Y(\us01\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us01/_1301_ ( .A1(\us01\/_0749_ ), .A2(\us01\/_0026_ ), .B1(\us01\/_0069_ ), .C1(\us01\/_0030_ ), .X(\us01\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us01/_1302_ ( .A1(\us01\/_0324_ ), .A2(\us01\/_0355_ ), .B1(\us01\/_0330_ ), .B2(\us01\/_0727_ ), .X(\us01\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us01/_1303_ ( .A(\us01\/_0133_ ), .B(\us01\/_0516_ ), .C(\us01\/_0517_ ), .Y(\us01\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1304_ ( .A(\us01\/_0509_ ), .B(\us01\/_0514_ ), .C(\us01\/_0515_ ), .D(\us01\/_0518_ ), .X(\us01\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1305_ ( .A(\us01\/_0746_ ), .B(\us01\/_0072_ ), .Y(\us01\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1306_ ( .A1(\us01\/_0082_ ), .A2(\us01\/_0070_ ), .B1(\us01\/_0043_ ), .B2(\us01\/_0193_ ), .Y(\us01\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1307_ ( .A(\us01\/_0311_ ), .B(\us01\/_0520_ ), .C(\us01\/_0332_ ), .D(\us01\/_0522_ ), .X(\us01\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1308_ ( .A(\us01\/_0129_ ), .B(\us01\/_0218_ ), .X(\us01\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_1309_ ( .A(\us01\/_0235_ ), .B(\us01\/_0524_ ), .Y(\us01\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us01/_1310_ ( .A(\us01\/_0081_ ), .B(\us01\/_0085_ ), .Y(\us01\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1311_ ( .A1(\us01\/_0051_ ), .A2(\us01\/_0045_ ), .B1(\us01\/_0130_ ), .B2(\us01\/_0094_ ), .Y(\us01\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1312_ ( .A(\us01\/_0523_ ), .B(\us01\/_0525_ ), .C(\us01\/_0526_ ), .D(\us01\/_0527_ ), .X(\us01\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us01/_1313_ ( .A_N(\us01\/_0250_ ), .B(\us01\/_0521_ ), .Y(\us01\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1314_ ( .A(\us01\/_0128_ ), .B(\us01\/_0020_ ), .X(\us01\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1315_ ( .A(\us01\/_0530_ ), .Y(\us01\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1316_ ( .A(\us01\/_0099_ ), .B(\us01\/_0058_ ), .X(\us01\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1317_ ( .A(\us01\/_0533_ ), .Y(\us01\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us01/_1318_ ( .A_N(\us01\/_0529_ ), .B(\us01\/_0531_ ), .C(\us01\/_0534_ ), .D(\us01\/_0192_ ), .X(\us01\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1319_ ( .A(\us01\/_0434_ ), .B(\us01\/_0078_ ), .X(\us01\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us01/_1320_ ( .A1(\us01\/_0750_ ), .A2(\us01\/_0079_ ), .B1(\us01\/_0129_ ), .B2(\us01\/_0705_ ), .X(\us01\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1321_ ( .A1(\us01\/_0161_ ), .A2(\us01\/_0030_ ), .B1(\us01\/_0536_ ), .C1(\us01\/_0537_ ), .Y(\us01\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us01/_1322_ ( .A1(\us01\/_0746_ ), .A2(\us01\/_0162_ ), .B1(\us01\/_0079_ ), .B2(\us01\/_0043_ ), .X(\us01\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1323_ ( .A1(\us01\/_0093_ ), .A2(\us01\/_0029_ ), .B1(\us01\/_0240_ ), .C1(\us01\/_0539_ ), .Y(\us01\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1324_ ( .A(\us01\/_0434_ ), .B(\us01\/_0043_ ), .X(\us01\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us01/_1325_ ( .A1(\us01\/_0142_ ), .A2(\us01\/_0150_ ), .B1(\us01\/_0022_ ), .B2(\us01\/_0137_ ), .X(\us01\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1326_ ( .A1(\us01\/_0279_ ), .A2(\us01\/_0051_ ), .B1(\us01\/_0541_ ), .C1(\us01\/_0542_ ), .Y(\us01\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1327_ ( .A(\us01\/_0159_ ), .B(\us01\/_0035_ ), .X(\us01\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us01/_1328_ ( .A1(\us01\/_0271_ ), .A2(\us01\/_0434_ ), .B1(\us01\/_0027_ ), .X(\us01\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1329_ ( .A1(\us01\/_0091_ ), .A2(\us01\/_0128_ ), .B1(\us01\/_0545_ ), .C1(\us01\/_0546_ ), .Y(\us01\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1330_ ( .A(\us01\/_0538_ ), .B(\us01\/_0540_ ), .C(\us01\/_0544_ ), .D(\us01\/_0547_ ), .X(\us01\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1331_ ( .A(\us01\/_0099_ ), .B(\us01\/_0193_ ), .X(\us01\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us01/_1332_ ( .A(\us01\/_0549_ ), .B(\us01\/_0186_ ), .C(\us01\/_0187_ ), .Y(\us01\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1333_ ( .A(\us01\/_0062_ ), .B(\us01\/_0347_ ), .C(\us01\/_0749_ ), .D(\us01\/_0694_ ), .X(\us01\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1334_ ( .A1(\us01\/_0130_ ), .A2(\us01\/_0218_ ), .B1(\us01\/_0551_ ), .C1(\us01\/_0101_ ), .Y(\us01\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1335_ ( .A(\us01\/_0139_ ), .B(\us01\/_0640_ ), .Y(\us01\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1336_ ( .A1(\us01\/_0752_ ), .A2(\us01\/_0662_ ), .B1(\us01\/_0280_ ), .B2(\us01\/_0099_ ), .Y(\us01\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1337_ ( .A(\us01\/_0550_ ), .B(\us01\/_0552_ ), .C(\us01\/_0553_ ), .D(\us01\/_0555_ ), .X(\us01\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1338_ ( .A(\us01\/_0528_ ), .B(\us01\/_0535_ ), .C(\us01\/_0548_ ), .D(\us01\/_0556_ ), .X(\us01\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us01/_1339_ ( .A(\us01\/_0504_ ), .B(\us01\/_0519_ ), .C(\us01\/_0557_ ), .Y(\us01\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1340_ ( .A(\us01\/_0054_ ), .B(\us01\/_0507_ ), .X(\us01\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us01/_1341_ ( .A_N(\us01\/_0558_ ), .B(\us01\/_0408_ ), .C(\us01\/_0451_ ), .D(\us01\/_0452_ ), .X(\us01\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1342_ ( .A(\us01\/_0549_ ), .Y(\us01\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1343_ ( .A(\us01\/_0559_ ), .B(\us01\/_0403_ ), .C(\us01\/_0560_ ), .D(\us01\/_0371_ ), .X(\us01\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1344_ ( .A(\us01\/_0181_ ), .B(\us01\/_0178_ ), .X(\us01\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1345_ ( .A(\us01\/_0562_ ), .B(\us01\/_0552_ ), .C(\us01\/_0553_ ), .D(\us01\/_0555_ ), .X(\us01\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1346_ ( .A(\us01\/_0029_ ), .B(\us01\/_0020_ ), .Y(\us01\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1347_ ( .A(\us01\/_0051_ ), .B(\us01\/_0130_ ), .X(\us01\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1348_ ( .A(\us01\/_0566_ ), .Y(\us01\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1349_ ( .A(\us01\/_0159_ ), .B(\us01\/_0412_ ), .X(\us01\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1350_ ( .A1(\us01\/_0752_ ), .A2(\us01\/_0640_ ), .B1(\us01\/_0568_ ), .B2(\us01\/_0175_ ), .Y(\us01\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1351_ ( .A(\us01\/_0076_ ), .B(\us01\/_0565_ ), .C(\us01\/_0567_ ), .D(\us01\/_0569_ ), .X(\us01\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us01/_1352_ ( .A1(\us01\/_0035_ ), .A2(\us01\/_0142_ ), .B1(\us01\/_0161_ ), .X(\us01\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1353_ ( .A(\us01\/_0099_ ), .B(\us01\/_0662_ ), .Y(\us01\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us01/_1354_ ( .A(\us01\/_0420_ ), .B(\us01\/_0571_ ), .C_N(\us01\/_0572_ ), .Y(\us01\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1355_ ( .A(\us01\/_0051_ ), .B(\us01\/_0746_ ), .Y(\us01\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1356_ ( .A(\us01\/_0574_ ), .B(\us01\/_0319_ ), .C(\us01\/_0320_ ), .D(\us01\/_0411_ ), .X(\us01\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1357_ ( .A(\us01\/_0736_ ), .B(\us01\/_0035_ ), .Y(\us01\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1358_ ( .A(\us01\/_0736_ ), .B(\us01\/_0030_ ), .Y(\us01\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1359_ ( .A(\us01\/_0298_ ), .B(\us01\/_0208_ ), .C(\us01\/_0577_ ), .D(\us01\/_0578_ ), .X(\us01\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1360_ ( .A1(\us01\/_0020_ ), .A2(\us01\/_0137_ ), .B1(\us01\/_0261_ ), .B2(\us01\/_0128_ ), .Y(\us01\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1361_ ( .A(\us01\/_0573_ ), .B(\us01\/_0576_ ), .C(\us01\/_0579_ ), .D(\us01\/_0580_ ), .X(\us01\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1362_ ( .A(\us01\/_0561_ ), .B(\us01\/_0563_ ), .C(\us01\/_0570_ ), .D(\us01\/_0581_ ), .X(\us01\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1363_ ( .A(\us01\/_0128_ ), .B(\us01\/_0193_ ), .X(\us01\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1364_ ( .A(\us01\/_0082_ ), .B(\us01\/_0162_ ), .X(\us01\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us01/_1365_ ( .A(\us01\/_0583_ ), .B(\us01\/_0584_ ), .C_N(\us01\/_0437_ ), .Y(\us01\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us01/_1366_ ( .A(\us01\/_0150_ ), .B(\us01\/_0118_ ), .C(\us01\/_0380_ ), .Y(\us01\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us01/_1367_ ( .A_N(\us01\/_0182_ ), .B(\us01\/_0587_ ), .C(\us01\/_0323_ ), .X(\us01\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1368_ ( .A1(\us01\/_0575_ ), .A2(\us01\/_0153_ ), .B1(\us01\/_0727_ ), .B2(\us01\/_0058_ ), .Y(\us01\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1369_ ( .A1(\us01\/_0218_ ), .A2(\us01\/_0064_ ), .B1(\us01\/_0134_ ), .B2(\us01\/_0255_ ), .Y(\us01\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1370_ ( .A(\us01\/_0585_ ), .B(\us01\/_0588_ ), .C(\us01\/_0589_ ), .D(\us01\/_0590_ ), .X(\us01\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us01/_1371_ ( .A1(\us01\/_0091_ ), .A2(\us01\/_0139_ ), .B1(\us01\/_0250_ ), .Y(\us01\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1372_ ( .A1(\us01\/_0092_ ), .A2(\us01\/_0739_ ), .B1(\us01\/_0324_ ), .B2(\us01\/_0029_ ), .Y(\us01\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1373_ ( .A1(\us01\/_0144_ ), .A2(\us01\/_0153_ ), .B1(\us01\/_0683_ ), .B2(\us01\/_0292_ ), .Y(\us01\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1374_ ( .A1(\us01\/_0091_ ), .A2(\us01\/_0218_ ), .B1(\us01\/_0330_ ), .B2(\us01\/_0292_ ), .Y(\us01\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1375_ ( .A(\us01\/_0592_ ), .B(\us01\/_0593_ ), .C(\us01\/_0594_ ), .D(\us01\/_0595_ ), .X(\us01\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1376_ ( .A(\us01\/_0218_ ), .B(\us01\/_0144_ ), .Y(\us01\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1377_ ( .A(\us01\/_0312_ ), .B(\us01\/_0598_ ), .Y(\us01\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1378_ ( .A(\us01\/_0575_ ), .B(\us01\/_0147_ ), .Y(\us01\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1379_ ( .A1(\us01\/_0293_ ), .A2(\us01\/_0137_ ), .B1(\us01\/_0093_ ), .B2(\us01\/_0739_ ), .Y(\us01\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1380_ ( .A1(\us01\/_0734_ ), .A2(\us01\/_0531_ ), .B1(\us01\/_0600_ ), .C1(\us01\/_0601_ ), .Y(\us01\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1381_ ( .A1(\us01\/_0153_ ), .A2(\us01\/_0261_ ), .B1(\us01\/_0599_ ), .C1(\us01\/_0602_ ), .Y(\us01\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1382_ ( .A(\us01\/_0591_ ), .B(\us01\/_0596_ ), .C(\us01\/_0174_ ), .D(\us01\/_0603_ ), .X(\us01\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1383_ ( .A(\us01\/_0029_ ), .B(\us01\/_0144_ ), .Y(\us01\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1384_ ( .A(\us01\/_0113_ ), .B(\us01\/_0017_ ), .Y(\us01\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1385_ ( .A(\us01\/_0381_ ), .B(\us01\/_0605_ ), .C(\us01\/_0361_ ), .D(\us01\/_0606_ ), .X(\us01\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1386_ ( .A1(\us01\/_0016_ ), .A2(\us01\/_0727_ ), .B1(\us01\/_0733_ ), .Y(\us01\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1387_ ( .A1(\us01\/_0586_ ), .A2(\us01\/_0159_ ), .B1(\us01\/_0082_ ), .B2(\us01\/_0750_ ), .Y(\us01\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1388_ ( .A1(\us01\/_0142_ ), .A2(\us01\/_0162_ ), .B1(\us01\/_0079_ ), .B2(\us01\/_0054_ ), .Y(\us01\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1389_ ( .A(\us01\/_0610_ ), .B(\us01\/_0611_ ), .C(\us01\/_0105_ ), .D(\us01\/_0106_ ), .X(\us01\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1390_ ( .A1(\us01\/_0094_ ), .A2(\us01\/_0302_ ), .B1(\us01\/_0324_ ), .B2(\us01\/_0089_ ), .Y(\us01\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1391_ ( .A(\us01\/_0607_ ), .B(\us01\/_0609_ ), .C(\us01\/_0612_ ), .D(\us01\/_0613_ ), .X(\us01\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1392_ ( .A(\us01\/_0041_ ), .B(\us01\/_0170_ ), .X(\us01\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1393_ ( .A(\us01\/_0554_ ), .B(\us01\/_0027_ ), .X(\us01\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1394_ ( .A(\us01\/_0027_ ), .B(\us01\/_0261_ ), .Y(\us01\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us01/_1395_ ( .A_N(\us01\/_0616_ ), .B(\us01\/_0617_ ), .Y(\us01\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1396_ ( .A1(\us01\/_0147_ ), .A2(\us01\/_0302_ ), .B1(\us01\/_0342_ ), .C1(\us01\/_0618_ ), .Y(\us01\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1397_ ( .A(\us01\/_0614_ ), .B(\us01\/_0272_ ), .C(\us01\/_0615_ ), .D(\us01\/_0620_ ), .X(\us01\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us01/_1398_ ( .A(\us01\/_0582_ ), .B(\us01\/_0604_ ), .C(\us01\/_0621_ ), .Y(\us01\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1399_ ( .A1(\us01\/_0280_ ), .A2(\us01\/_0134_ ), .B1(\us01\/_0089_ ), .Y(\us01\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1400_ ( .A1(\us01\/_0144_ ), .A2(\us01\/_0608_ ), .A3(\us01\/_0330_ ), .B1(\us01\/_0089_ ), .Y(\us01\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1401_ ( .A1(\us01\/_0197_ ), .A2(\us01\/_0130_ ), .A3(\us01\/_0110_ ), .B1(\us01\/_0094_ ), .Y(\us01\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1402_ ( .A(\us01\/_0432_ ), .B(\us01\/_0622_ ), .C(\us01\/_0623_ ), .D(\us01\/_0624_ ), .X(\us01\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us01/_1403_ ( .A1(\us01\/_0554_ ), .A2(\us01\/_0017_ ), .A3(\us01\/_0022_ ), .B1(\us01\/_0161_ ), .X(\us01\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us01/_1404_ ( .A_N(\us01\/_0269_ ), .B(\us01\/_0170_ ), .X(\us01\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1405_ ( .A1(\us01\/_0109_ ), .A2(\us01\/_0064_ ), .A3(\us01\/_0733_ ), .B1(\us01\/_0355_ ), .Y(\us01\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us01/_1406_ ( .A_N(\us01\/_0626_ ), .B(\us01\/_0627_ ), .C(\us01\/_0353_ ), .D(\us01\/_0628_ ), .X(\us01\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1407_ ( .A1(\us01\/_0091_ ), .A2(\us01\/_0110_ ), .A3(\us01\/_0176_ ), .B1(\us01\/_0139_ ), .Y(\us01\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1408_ ( .A1(\us01\/_0020_ ), .A2(\us01\/_0261_ ), .B1(\us01\/_0147_ ), .Y(\us01\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1409_ ( .A(\us01\/_0631_ ), .B(\us01\/_0344_ ), .C(\us01\/_0421_ ), .D(\us01\/_0632_ ), .X(\us01\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us01/_1410_ ( .A1(\us01\/_0325_ ), .A2(\us01\/_0734_ ), .B1(\us01\/_0038_ ), .C1(\us01\/_0113_ ), .X(\us01\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1411_ ( .A1(\us01\/_0134_ ), .A2(\us01\/_0114_ ), .B1(\us01\/_0221_ ), .C1(\us01\/_0634_ ), .Y(\us01\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us01/_1412_ ( .A(\us01\/_0119_ ), .B_N(\us01\/_0111_ ), .Y(\us01\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1413_ ( .A1(\us01\/_0030_ ), .A2(\us01\/_0113_ ), .B1(\us01\/_0636_ ), .C1(\us01\/_0400_ ), .Y(\us01\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1414_ ( .A1(\us01\/_0731_ ), .A2(\us01\/_0293_ ), .A3(\us01\/_0251_ ), .B1(\us01\/_0099_ ), .Y(\us01\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1415_ ( .A(\us01\/_0189_ ), .B(\us01\/_0635_ ), .C(\us01\/_0637_ ), .D(\us01\/_0638_ ), .X(\us01\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1416_ ( .A(\us01\/_0625_ ), .B(\us01\/_0630_ ), .C(\us01\/_0633_ ), .D(\us01\/_0639_ ), .X(\us01\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1417_ ( .A(\us01\/_0746_ ), .B(\us01\/_0738_ ), .X(\us01\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1418_ ( .A(\us01\/_0736_ ), .B(\us01\/_0731_ ), .X(\us01\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us01/_1419_ ( .A_N(\us01\/_0643_ ), .B(\us01\/_0577_ ), .Y(\us01\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1420_ ( .A1(\us01\/_0280_ ), .A2(\us01\/_0739_ ), .B1(\us01\/_0642_ ), .C1(\us01\/_0644_ ), .Y(\us01\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1421_ ( .A1(\us01\/_0050_ ), .A2(\us01\/_0249_ ), .B1(\us01\/_0194_ ), .C1(\us01\/_0738_ ), .Y(\us01\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1422_ ( .A(\us01\/_0646_ ), .B(\us01\/_0232_ ), .C(\us01\/_0417_ ), .D(\us01\/_0578_ ), .X(\us01\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1423_ ( .A1(\us01\/_0064_ ), .A2(\us01\/_0733_ ), .B1(\us01\/_0727_ ), .Y(\us01\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1424_ ( .A1(\us01\/_0193_ ), .A2(\us01\/_0276_ ), .B1(\us01\/_0727_ ), .Y(\us01\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1425_ ( .A(\us01\/_0645_ ), .B(\us01\/_0647_ ), .C(\us01\/_0648_ ), .D(\us01\/_0649_ ), .X(\us01\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1426_ ( .A1(\us01\/_0325_ ), .A2(\us01\/_0734_ ), .B1(\us01\/_0038_ ), .C1(\us01\/_0029_ ), .Y(\us01\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1427_ ( .A1(\us01\/_0249_ ), .A2(\us01\/_0205_ ), .B1(\us01\/_0412_ ), .C1(\us01\/_0029_ ), .Y(\us01\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1428_ ( .A(\us01\/_0652_ ), .B(\us01\/_0653_ ), .X(\us01\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1429_ ( .A1(\us01\/_0733_ ), .A2(\us01\/_0748_ ), .A3(\us01\/_0324_ ), .B1(\us01\/_0016_ ), .Y(\us01\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1430_ ( .A1(\us01\/_0640_ ), .A2(\us01\/_0193_ ), .A3(\us01\/_0091_ ), .B1(\us01\/_0016_ ), .Y(\us01\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1431_ ( .A1(\us01\/_0102_ ), .A2(\us01\/_0301_ ), .B1(\sa01\[3\] ), .C1(\us01\/_0029_ ), .Y(\us01\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1432_ ( .A(\us01\/_0654_ ), .B(\us01\/_0655_ ), .C(\us01\/_0656_ ), .D(\us01\/_0657_ ), .X(\us01\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1433_ ( .A1(\us01\/_0118_ ), .A2(\us01\/_0050_ ), .B1(\us01\/_0038_ ), .C1(\us01\/_0478_ ), .Y(\us01\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us01/_1434_ ( .A_N(\us01\/_0250_ ), .B(\us01\/_0465_ ), .C(\us01\/_0659_ ), .X(\us01\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1435_ ( .A1(\us01\/_0683_ ), .A2(\us01\/_0324_ ), .B1(\us01\/_0255_ ), .Y(\us01\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1436_ ( .A1(\us01\/_0030_ ), .A2(\us01\/_0193_ ), .A3(\us01\/_0047_ ), .B1(\us01\/_0255_ ), .Y(\us01\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1437_ ( .A1(\us01\/_0144_ ), .A2(\us01\/_0586_ ), .A3(\us01\/_0047_ ), .B1(\us01\/_0218_ ), .Y(\us01\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1438_ ( .A(\us01\/_0660_ ), .B(\us01\/_0661_ ), .C(\us01\/_0663_ ), .D(\us01\/_0664_ ), .X(\us01\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1439_ ( .A1(\us01\/_0091_ ), .A2(\us01\/_0276_ ), .B1(\us01\/_0060_ ), .Y(\us01\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1440_ ( .A1(\us01\/_0144_ ), .A2(\us01\/_0608_ ), .B1(\us01\/_0292_ ), .Y(\us01\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1441_ ( .A1(\us01\/_0412_ ), .A2(\us01\/_0038_ ), .B1(\us01\/_0102_ ), .C1(\us01\/_0060_ ), .Y(\us01\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1442_ ( .A1(\sa01\[1\] ), .A2(\us01\/_0734_ ), .B1(\us01\/_0109_ ), .C1(\us01\/_0292_ ), .Y(\us01\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1443_ ( .A(\us01\/_0666_ ), .B(\us01\/_0667_ ), .C(\us01\/_0668_ ), .D(\us01\/_0669_ ), .X(\us01\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1444_ ( .A(\us01\/_0650_ ), .B(\us01\/_0658_ ), .C(\us01\/_0665_ ), .D(\us01\/_0670_ ), .X(\us01\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us01/_1445_ ( .A(\us01\/_0641_ ), .B(\us01\/_0174_ ), .C(\us01\/_0671_ ), .Y(\us01\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us01/_1446_ ( .A(\us01\/_0049_ ), .B(\us01\/_0618_ ), .C_N(\us01\/_0052_ ), .Y(\us01\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us01/_1447_ ( .A(\us01\/_0239_ ), .Y(\us01\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1448_ ( .A(\us01\/_0705_ ), .B(\us01\/_0030_ ), .Y(\us01\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1449_ ( .A1(\us01\/_0054_ ), .A2(\us01\/_0731_ ), .B1(\us01\/_0035_ ), .B2(\us01\/_0705_ ), .Y(\us01\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1450_ ( .A1(\us01\/_0304_ ), .A2(\us01\/_0731_ ), .B1(\us01\/_0047_ ), .B2(\us01\/_0750_ ), .Y(\us01\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1451_ ( .A(\us01\/_0674_ ), .B(\us01\/_0675_ ), .C(\us01\/_0676_ ), .D(\us01\/_0677_ ), .X(\us01\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us01/_1452_ ( .A_N(\us01\/_0584_ ), .B(\us01\/_0283_ ), .X(\us01\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1453_ ( .A(\us01\/_0673_ ), .B(\us01\/_0678_ ), .C(\us01\/_0679_ ), .D(\us01\/_0508_ ), .X(\us01\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1454_ ( .A1(\us01\/_0016_ ), .A2(\us01\/_0733_ ), .B1(\us01\/_0355_ ), .B2(\us01\/_0092_ ), .Y(\us01\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1455_ ( .A(\us01\/_0681_ ), .B(\us01\/_0034_ ), .X(\us01\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us01/_1456_ ( .A1(\us01\/_0330_ ), .A2(\us01\/_0139_ ), .B1(\us01\/_0324_ ), .B2(\us01\/_0089_ ), .X(\us01\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1457_ ( .A1(\us01\/_0146_ ), .A2(\us01\/_0147_ ), .B1(\us01\/_0133_ ), .C1(\us01\/_0684_ ), .Y(\us01\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1458_ ( .A(\us01\/_0113_ ), .B(\us01\/_0251_ ), .Y(\us01\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us01/_1459_ ( .A_N(\us01\/_0463_ ), .B(\us01\/_0686_ ), .C(\us01\/_0383_ ), .D(\us01\/_0464_ ), .X(\us01\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1460_ ( .A1(\us01\/_0051_ ), .A2(\us01\/_0293_ ), .B1(\us01\/_0280_ ), .B2(\us01\/_0705_ ), .Y(\us01\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1461_ ( .A1(\us01\/_0017_ ), .A2(\us01\/_0072_ ), .B1(\us01\/_0134_ ), .B2(\us01\/_0078_ ), .Y(\us01\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1462_ ( .A(\us01\/_0687_ ), .B(\us01\/_0236_ ), .C(\us01\/_0688_ ), .D(\us01\/_0689_ ), .X(\us01\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1463_ ( .A(\us01\/_0680_ ), .B(\us01\/_0682_ ), .C(\us01\/_0685_ ), .D(\us01\/_0690_ ), .X(\us01\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us01/_1464_ ( .A1(\us01\/_0532_ ), .A2(\us01\/_0380_ ), .B1(\us01\/_0102_ ), .C1(\us01\/_0355_ ), .X(\us01\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us01/_1465_ ( .A(\us01\/_0692_ ), .B(\us01\/_0338_ ), .C(\us01\/_0644_ ), .Y(\us01\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1466_ ( .A(\us01\/_0016_ ), .B(\us01\/_0020_ ), .Y(\us01\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1467_ ( .A1(\us01\/_0030_ ), .A2(\us01\/_0137_ ), .B1(\us01\/_0279_ ), .B2(\us01\/_0094_ ), .Y(\us01\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1468_ ( .A1(\us01\/_0575_ ), .A2(\us01\/_0153_ ), .B1(\us01\/_0161_ ), .B2(\us01\/_0293_ ), .Y(\us01\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1469_ ( .A(\us01\/_0259_ ), .B(\us01\/_0695_ ), .C(\us01\/_0696_ ), .D(\us01\/_0697_ ), .X(\us01\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us01/_1470_ ( .A1(\us01\/_0255_ ), .A2(\us01\/_0640_ ), .B1(\us01\/_0016_ ), .B2(\us01\/_0193_ ), .X(\us01\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1471_ ( .A1(\us01\/_0060_ ), .A2(\us01\/_0176_ ), .B1(\us01\/_0699_ ), .C1(\us01\/_0177_ ), .Y(\us01\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1472_ ( .A1(\us01\/_0091_ ), .A2(\us01\/_0218_ ), .B1(\us01\/_0092_ ), .B2(\us01\/_0705_ ), .Y(\us01\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us01/_1473_ ( .A1(\us01\/_0705_ ), .A2(\us01\/_0683_ ), .B1(\us01\/_0093_ ), .B2(\us01\/_0114_ ), .Y(\us01\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us01/_1474_ ( .A1(\us01\/_0683_ ), .A2(\us01\/_0280_ ), .B1(\us01\/_0094_ ), .Y(\us01\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us01/_1475_ ( .A1(\us01\/_0249_ ), .A2(\us01\/_0205_ ), .B1(\us01\/_0038_ ), .C1(\us01\/_0292_ ), .Y(\us01\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1476_ ( .A(\us01\/_0701_ ), .B(\us01\/_0702_ ), .C(\us01\/_0703_ ), .D(\us01\/_0704_ ), .X(\us01\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1477_ ( .A(\us01\/_0693_ ), .B(\us01\/_0698_ ), .C(\us01\/_0700_ ), .D(\us01\/_0706_ ), .X(\us01\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us01/_1478_ ( .A1(\us01\/_0113_ ), .A2(\us01\/_0640_ ), .B1(\us01\/_0099_ ), .B2(\us01\/_0058_ ), .X(\us01\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us01/_1479_ ( .A(\us01\/_0407_ ), .B(\us01\/_0708_ ), .C(\us01\/_0529_ ), .Y(\us01\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1480_ ( .A(\us01\/_0568_ ), .B(\us01\/_0175_ ), .Y(\us01\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us01/_1481_ ( .A1(\us01\/_0029_ ), .A2(\us01\/_0114_ ), .A3(\us01\/_0051_ ), .B1(\us01\/_0130_ ), .Y(\us01\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1482_ ( .A(\us01\/_0709_ ), .B(\us01\/_0550_ ), .C(\us01\/_0710_ ), .D(\us01\/_0711_ ), .X(\us01\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us01/_1483_ ( .A1(\us01\/_0114_ ), .A2(\us01\/_0064_ ), .B1(\us01\/_0261_ ), .B2(\us01\/_0089_ ), .X(\us01\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1484_ ( .A1(\us01\/_0355_ ), .A2(\us01\/_0261_ ), .B1(\us01\/_0198_ ), .C1(\us01\/_0713_ ), .Y(\us01\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1485_ ( .A(\us01\/_0586_ ), .B(\us01\/_0478_ ), .Y(\us01\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us01/_1486_ ( .A_N(\us01\/_0541_ ), .B(\us01\/_0267_ ), .C(\us01\/_0715_ ), .D(\us01\/_0320_ ), .X(\us01\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1487_ ( .A(\us01\/_0586_ ), .B(\us01\/_0070_ ), .Y(\us01\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us01/_1488_ ( .A_N(\us01\/_0211_ ), .B(\us01\/_0155_ ), .C(\us01\/_0202_ ), .D(\us01\/_0718_ ), .X(\us01\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us01/_1489_ ( .A(\us01\/_0150_ ), .B(\us01\/_0205_ ), .C(\us01\/_0380_ ), .Y(\us01\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us01/_1490_ ( .A(\us01\/_0411_ ), .B(\us01\/_0720_ ), .X(\us01\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us01/_1491_ ( .A1(\us01\/_0017_ ), .A2(\us01\/_0022_ ), .B1(\us01\/_0078_ ), .X(\us01\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us01/_1492_ ( .A1(\us01\/_0134_ ), .A2(\us01\/_0738_ ), .B1(\us01\/_0101_ ), .C1(\us01\/_0722_ ), .Y(\us01\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1493_ ( .A(\us01\/_0717_ ), .B(\us01\/_0719_ ), .C(\us01\/_0721_ ), .D(\us01\/_0723_ ), .X(\us01\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us01/_1494_ ( .A(\us01\/_0739_ ), .B(\us01\/_0193_ ), .Y(\us01\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1495_ ( .A(\us01\/_0344_ ), .B(\us01\/_0184_ ), .C(\us01\/_0449_ ), .D(\us01\/_0725_ ), .X(\us01\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us01/_1496_ ( .A(\us01\/_0712_ ), .B(\us01\/_0714_ ), .C(\us01\/_0724_ ), .D(\us01\/_0726_ ), .X(\us01\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \us01/_1497_ ( .A(\us01\/_0691_ ), .B(\us01\/_0707_ ), .C(\us01\/_0728_ ), .Y(\us01\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \us02/_0753_ ( .A(\sa02\[2\] ), .B_N(\sa02\[3\] ), .Y(\us02\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \us02/_0755_ ( .A(\sa02\[1\] ), .B(\sa02\[0\] ), .X(\us02\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us02/_0756_ ( .A(\us02\/_0096_ ), .B(\us02\/_0118_ ), .X(\us02\/_0129_ ) );
sky130_fd_sc_hd__and2_1 \us02/_0757_ ( .A(\sa02\[7\] ), .B(\sa02\[6\] ), .X(\us02\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_0758_ ( .A(\sa02\[4\] ), .B(\sa02\[5\] ), .Y(\us02\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0759_ ( .A(\us02\/_0140_ ), .B(\us02\/_0151_ ), .X(\us02\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0761_ ( .A(\us02\/_0129_ ), .B(\us02\/_0162_ ), .X(\us02\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0762_ ( .A(\us02\/_0096_ ), .X(\us02\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \us02/_0763_ ( .A(\sa02\[1\] ), .B_N(\sa02\[0\] ), .Y(\us02\/_0205_ ) );
sky130_fd_sc_hd__and3_1 \us02/_0765_ ( .A(\us02\/_0162_ ), .B(\us02\/_0194_ ), .C(\us02\/_0205_ ), .X(\us02\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us02/_0766_ ( .A(\us02\/_0183_ ), .SLEEP(\us02\/_0227_ ), .X(\us02\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \us02/_0767_ ( .A(\sa02\[0\] ), .B_N(\sa02\[1\] ), .Y(\us02\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_0768_ ( .A(\sa02\[2\] ), .B(\sa02\[3\] ), .Y(\us02\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0769_ ( .A(\us02\/_0249_ ), .B(\us02\/_0260_ ), .X(\us02\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0771_ ( .A(\us02\/_0271_ ), .X(\us02\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0772_ ( .A(\us02\/_0162_ ), .X(\us02\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_0773_ ( .A(\us02\/_0293_ ), .B(\us02\/_0304_ ), .Y(\us02\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us02/_0774_ ( .A(\sa02\[1\] ), .Y(\us02\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us02/_0776_ ( .A(\sa02\[0\] ), .Y(\us02\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0777_ ( .A(\sa02\[2\] ), .B(\sa02\[3\] ), .X(\us02\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0779_ ( .A(\us02\/_0358_ ), .X(\us02\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_0780_ ( .A1(\us02\/_0325_ ), .A2(\us02\/_0347_ ), .B1(\us02\/_0380_ ), .C1(\us02\/_0304_ ), .Y(\us02\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us02/_0781_ ( .A_N(\us02\/_0238_ ), .B(\us02\/_0314_ ), .C(\us02\/_0391_ ), .X(\us02\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us02/_0782_ ( .A(\sa02\[3\] ), .B_N(\sa02\[2\] ), .Y(\us02\/_0412_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0784_ ( .A(\us02\/_0412_ ), .B(\us02\/_0205_ ), .X(\us02\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \us02/_0787_ ( .A(\sa02\[5\] ), .B_N(\sa02\[4\] ), .Y(\us02\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0788_ ( .A(\us02\/_0467_ ), .B(\us02\/_0140_ ), .X(\us02\/_0478_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_0791_ ( .A(\us02\/_0134_ ), .B(\us02\/_0218_ ), .Y(\us02\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_0792_ ( .A(\us02\/_0478_ ), .B(\us02\/_0271_ ), .Y(\us02\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0793_ ( .A(\us02\/_0194_ ), .X(\us02\/_0532_ ) );
sky130_fd_sc_hd__and2_1 \us02/_0795_ ( .A(\us02\/_0249_ ), .B(\us02\/_0358_ ), .X(\us02\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0797_ ( .A(\us02\/_0554_ ), .X(\us02\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us02/_0798_ ( .A(\us02\/_0205_ ), .B(\us02\/_0358_ ), .X(\us02\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0800_ ( .A(\us02\/_0586_ ), .X(\us02\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_0801_ ( .A1(\us02\/_0532_ ), .A2(\us02\/_0575_ ), .A3(\us02\/_0608_ ), .B1(\us02\/_0218_ ), .Y(\us02\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us02/_0802_ ( .A(\us02\/_0401_ ), .B(\us02\/_0510_ ), .C(\us02\/_0521_ ), .D(\us02\/_0619_ ), .X(\us02\/_0629_ ) );
sky130_fd_sc_hd__and2_1 \us02/_0803_ ( .A(\us02\/_0358_ ), .B(\sa02\[1\] ), .X(\us02\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0805_ ( .A(\us02\/_0205_ ), .B(\us02\/_0260_ ), .X(\us02\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0807_ ( .A(\us02\/_0662_ ), .X(\us02\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us02/_0808_ ( .A(\sa02\[6\] ), .B_N(\sa02\[7\] ), .Y(\us02\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \us02/_0809_ ( .A(\us02\/_0467_ ), .B(\us02\/_0694_ ), .X(\us02\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0811_ ( .A(\us02\/_0705_ ), .X(\us02\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_0812_ ( .A1(\us02\/_0640_ ), .A2(\us02\/_0293_ ), .A3(\us02\/_0683_ ), .B1(\us02\/_0727_ ), .Y(\us02\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_0813_ ( .A(\sa02\[1\] ), .B(\sa02\[0\] ), .Y(\us02\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0814_ ( .A(\us02\/_0730_ ), .B(\us02\/_0260_ ), .X(\us02\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0816_ ( .A(\us02\/_0731_ ), .X(\us02\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0817_ ( .A(\sa02\[0\] ), .X(\us02\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us02/_0818_ ( .A1(\us02\/_0325_ ), .A2(\us02\/_0734_ ), .B1(\us02\/_0412_ ), .X(\us02\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0819_ ( .A(\us02\/_0694_ ), .B(\us02\/_0151_ ), .X(\us02\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0821_ ( .A(\us02\/_0736_ ), .X(\us02\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0822_ ( .A(\us02\/_0738_ ), .X(\us02\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_0823_ ( .A1(\us02\/_0733_ ), .A2(\us02\/_0735_ ), .A3(\us02\/_0293_ ), .B1(\us02\/_0739_ ), .Y(\us02\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us02/_0824_ ( .A(\us02\/_0730_ ), .B_N(\us02\/_0358_ ), .Y(\us02\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_0825_ ( .A(\us02\/_0741_ ), .B(\us02\/_0739_ ), .Y(\us02\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_0827_ ( .A1(\us02\/_0118_ ), .A2(\us02\/_0205_ ), .B1(\us02\/_0532_ ), .C1(\us02\/_0739_ ), .Y(\us02\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us02/_0828_ ( .A(\us02\/_0729_ ), .B(\us02\/_0740_ ), .C(\us02\/_0742_ ), .D(\us02\/_0744_ ), .X(\us02\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0829_ ( .A(\us02\/_0412_ ), .B(\us02\/_0730_ ), .X(\us02\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0831_ ( .A(\us02\/_0746_ ), .X(\us02\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us02/_0832_ ( .A(\sa02\[4\] ), .B_N(\sa02\[5\] ), .Y(\us02\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0833_ ( .A(\us02\/_0749_ ), .B(\us02\/_0694_ ), .X(\us02\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0835_ ( .A(\us02\/_0750_ ), .X(\us02\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0836_ ( .A(\us02\/_0752_ ), .X(\us02\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0837_ ( .A(\us02\/_0118_ ), .B(\us02\/_0358_ ), .X(\us02\/_0017_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0839_ ( .A(\us02\/_0752_ ), .B(\us02\/_0017_ ), .X(\us02\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0840_ ( .A(\us02\/_0358_ ), .B(\us02\/_0325_ ), .X(\us02\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0842_ ( .A(\us02\/_0096_ ), .B(\us02\/_0205_ ), .X(\us02\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \us02/_0844_ ( .A1(\us02\/_0020_ ), .A2(\us02\/_0022_ ), .B1(\us02\/_0752_ ), .X(\us02\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_0845_ ( .A1(\us02\/_0748_ ), .A2(\us02\/_0016_ ), .B1(\us02\/_0019_ ), .C1(\us02\/_0024_ ), .Y(\us02\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \us02/_0846_ ( .A(\sa02\[4\] ), .B(\sa02\[5\] ), .X(\us02\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0847_ ( .A(\us02\/_0694_ ), .B(\us02\/_0026_ ), .X(\us02\/_0027_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0850_ ( .A(\us02\/_0358_ ), .B(\us02\/_0730_ ), .X(\us02\/_0030_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0852_ ( .A(\us02\/_0030_ ), .X(\us02\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_0853_ ( .A(\us02\/_0247_ ), .B(\us02\/_0032_ ), .Y(\us02\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_0854_ ( .A(\us02\/_0247_ ), .B(\us02\/_0735_ ), .Y(\us02\/_0034_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0855_ ( .A(\us02\/_0118_ ), .B(\us02\/_0260_ ), .X(\us02\/_0035_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0857_ ( .A(\us02\/_0027_ ), .B(\us02\/_0035_ ), .X(\us02\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0858_ ( .A(\us02\/_0260_ ), .X(\us02\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_0859_ ( .A(\us02\/_0038_ ), .B(\us02\/_0347_ ), .Y(\us02\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us02/_0860_ ( .A_N(\us02\/_0039_ ), .B(\us02\/_0027_ ), .X(\us02\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_0861_ ( .A(\us02\/_0037_ ), .B(\us02\/_0040_ ), .Y(\us02\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us02/_0862_ ( .A(\us02\/_0025_ ), .B(\us02\/_0033_ ), .C(\us02\/_0034_ ), .D(\us02\/_0041_ ), .X(\us02\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0863_ ( .A(\us02\/_0749_ ), .B(\us02\/_0140_ ), .X(\us02\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us02/_0865_ ( .A(\sa02\[0\] ), .B(\sa02\[2\] ), .C(\sa02\[3\] ), .X(\us02\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0866_ ( .A(\us02\/_0043_ ), .B(\us02\/_0045_ ), .X(\us02\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0867_ ( .A(\us02\/_0096_ ), .B(\us02\/_0249_ ), .X(\us02\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0869_ ( .A(\us02\/_0047_ ), .B(\us02\/_0043_ ), .X(\us02\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0870_ ( .A(\us02\/_0730_ ), .X(\us02\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0871_ ( .A(\us02\/_0043_ ), .X(\us02\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_0872_ ( .A1(\us02\/_0118_ ), .A2(\us02\/_0050_ ), .B1(\us02\/_0194_ ), .C1(\us02\/_0051_ ), .Y(\us02\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us02/_0873_ ( .A(\us02\/_0046_ ), .B(\us02\/_0049_ ), .C_N(\us02\/_0052_ ), .Y(\us02\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0874_ ( .A(\us02\/_0026_ ), .B(\us02\/_0140_ ), .X(\us02\/_0054_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0876_ ( .A(\us02\/_0054_ ), .X(\us02\/_0056_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_0877_ ( .A1(\us02\/_0532_ ), .A2(\us02\/_0575_ ), .B1(\us02\/_0056_ ), .Y(\us02\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0878_ ( .A(\us02\/_0412_ ), .B(\us02\/_0325_ ), .X(\us02\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0880_ ( .A(\us02\/_0051_ ), .X(\us02\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_0881_ ( .A1(\us02\/_0731_ ), .A2(\us02\/_0035_ ), .A3(\us02\/_0058_ ), .B1(\us02\/_0060_ ), .Y(\us02\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0882_ ( .A(\us02\/_0260_ ), .B(\sa02\[1\] ), .X(\us02\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0884_ ( .A(\us02\/_0062_ ), .X(\us02\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_0885_ ( .A1(\us02\/_0064_ ), .A2(\us02\/_0748_ ), .A3(\us02\/_0683_ ), .B1(\us02\/_0056_ ), .Y(\us02\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us02/_0886_ ( .A(\us02\/_0053_ ), .B(\us02\/_0057_ ), .C(\us02\/_0061_ ), .D(\us02\/_0065_ ), .X(\us02\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us02/_0887_ ( .A(\us02\/_0629_ ), .B(\us02\/_0745_ ), .C(\us02\/_0042_ ), .D(\us02\/_0066_ ), .X(\us02\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us02/_0889_ ( .A(\sa02\[7\] ), .B_N(\sa02\[6\] ), .Y(\us02\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0890_ ( .A(\us02\/_0069_ ), .B(\us02\/_0151_ ), .X(\us02\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0892_ ( .A(\us02\/_0070_ ), .X(\us02\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_0893_ ( .A1(\us02\/_0129_ ), .A2(\us02\/_0586_ ), .B1(\us02\/_0072_ ), .Y(\us02\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_0894_ ( .A1(\us02\/_0380_ ), .A2(\us02\/_0347_ ), .B1(\us02\/_0194_ ), .B2(\us02\/_0205_ ), .Y(\us02\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us02/_0895_ ( .A(\us02\/_0074_ ), .B_N(\us02\/_0070_ ), .Y(\us02\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us02/_0896_ ( .A(\us02\/_0073_ ), .SLEEP(\us02\/_0075_ ), .X(\us02\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us02/_0897_ ( .A(\us02\/_0467_ ), .B(\us02\/_0069_ ), .X(\us02\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0898_ ( .A(\us02\/_0077_ ), .X(\us02\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0899_ ( .A(\us02\/_0412_ ), .B(\us02\/_0118_ ), .X(\us02\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0901_ ( .A(\us02\/_0078_ ), .B(\us02\/_0079_ ), .X(\us02\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0902_ ( .A(\us02\/_0412_ ), .B(\us02\/_0249_ ), .X(\us02\/_0082_ ) );
sky130_fd_sc_hd__buf_2 \us02/_0904_ ( .A(\us02\/_0082_ ), .X(\us02\/_0084_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0905_ ( .A(\us02\/_0084_ ), .B(\us02\/_0078_ ), .X(\us02\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us02/_0906_ ( .A1(\sa02\[0\] ), .A2(\us02\/_0325_ ), .B1(\us02\/_0260_ ), .Y(\us02\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us02/_0907_ ( .A_N(\us02\/_0086_ ), .B(\us02\/_0078_ ), .X(\us02\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us02/_0908_ ( .A(\us02\/_0081_ ), .B(\us02\/_0085_ ), .C(\us02\/_0087_ ), .Y(\us02\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0909_ ( .A(\us02\/_0072_ ), .X(\us02\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_0910_ ( .A1(\us02\/_0733_ ), .A2(\us02\/_0748_ ), .A3(\us02\/_0683_ ), .B1(\us02\/_0089_ ), .Y(\us02\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0911_ ( .A(\us02\/_0129_ ), .X(\us02\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0912_ ( .A(\us02\/_0017_ ), .X(\us02\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0913_ ( .A(\us02\/_0022_ ), .X(\us02\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0914_ ( .A(\us02\/_0078_ ), .X(\us02\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_0915_ ( .A1(\us02\/_0091_ ), .A2(\us02\/_0092_ ), .A3(\us02\/_0093_ ), .B1(\us02\/_0094_ ), .Y(\us02\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us02/_0916_ ( .A(\us02\/_0076_ ), .B(\us02\/_0088_ ), .C(\us02\/_0090_ ), .D(\us02\/_0095_ ), .X(\us02\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us02/_0917_ ( .A(\us02\/_0069_ ), .B(\us02\/_0026_ ), .X(\us02\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \us02/_0918_ ( .A(\us02\/_0098_ ), .X(\us02\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0919_ ( .A(\us02\/_0434_ ), .B(\us02\/_0099_ ), .X(\us02\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0920_ ( .A(\us02\/_0079_ ), .B(\us02\/_0098_ ), .X(\us02\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0921_ ( .A(\us02\/_0325_ ), .X(\us02\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_0922_ ( .A1(\us02\/_0102_ ), .A2(\us02\/_0734_ ), .B1(\us02\/_0038_ ), .C1(\us02\/_0099_ ), .Y(\us02\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us02/_0923_ ( .A(\us02\/_0100_ ), .B(\us02\/_0101_ ), .C_N(\us02\/_0103_ ), .Y(\us02\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_0924_ ( .A1(\us02\/_0554_ ), .A2(\us02\/_0586_ ), .B1(\us02\/_0099_ ), .Y(\us02\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_0925_ ( .A(\us02\/_0129_ ), .B(\us02\/_0099_ ), .Y(\us02\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0926_ ( .A(\us02\/_0105_ ), .B(\us02\/_0106_ ), .X(\us02\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0927_ ( .A(\us02\/_0412_ ), .X(\us02\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us02/_0928_ ( .A(\us02\/_0260_ ), .B(\sa02\[0\] ), .X(\us02\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0929_ ( .A(\us02\/_0069_ ), .B(\us02\/_0749_ ), .X(\us02\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0931_ ( .A(\us02\/_0111_ ), .X(\us02\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0932_ ( .A(\us02\/_0113_ ), .X(\us02\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_0933_ ( .A1(\us02\/_0109_ ), .A2(\us02\/_0110_ ), .B1(\us02\/_0114_ ), .Y(\us02\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us02/_0934_ ( .A(\us02\/_0022_ ), .Y(\us02\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us02/_0935_ ( .A(\us02\/_0554_ ), .Y(\us02\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us02/_0936_ ( .A1(\us02\/_0050_ ), .A2(\us02\/_0118_ ), .B1(\us02\/_0194_ ), .Y(\us02\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us02/_0937_ ( .A(\us02\/_0113_ ), .Y(\us02\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us02/_0938_ ( .A1(\us02\/_0116_ ), .A2(\us02\/_0117_ ), .A3(\us02\/_0119_ ), .B1(\us02\/_0120_ ), .X(\us02\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us02/_0939_ ( .A(\us02\/_0104_ ), .B(\us02\/_0108_ ), .C(\us02\/_0115_ ), .D(\us02\/_0121_ ), .X(\us02\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_0940_ ( .A(\sa02\[7\] ), .B(\sa02\[6\] ), .Y(\us02\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0941_ ( .A(\us02\/_0749_ ), .B(\us02\/_0123_ ), .X(\us02\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0943_ ( .A(\us02\/_0082_ ), .B(\us02\/_0124_ ), .X(\us02\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_0944_ ( .A(\us02\/_0271_ ), .B(\us02\/_0124_ ), .Y(\us02\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0945_ ( .A(\us02\/_0124_ ), .X(\us02\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0946_ ( .A(\us02\/_0260_ ), .B(\us02\/_0325_ ), .X(\us02\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_0948_ ( .A(\us02\/_0128_ ), .B(\us02\/_0130_ ), .Y(\us02\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_0949_ ( .A(\us02\/_0127_ ), .B(\us02\/_0132_ ), .Y(\us02\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us02/_0950_ ( .A(\us02\/_0434_ ), .X(\us02\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_0951_ ( .A(\us02\/_0134_ ), .B(\us02\/_0128_ ), .Y(\us02\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us02/_0952_ ( .A(\us02\/_0126_ ), .B(\us02\/_0133_ ), .C_N(\us02\/_0135_ ), .Y(\us02\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us02/_0953_ ( .A(\us02\/_0026_ ), .B(\us02\/_0123_ ), .X(\us02\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0955_ ( .A(\us02\/_0137_ ), .X(\us02\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_0956_ ( .A1(\us02\/_0110_ ), .A2(\us02\/_0293_ ), .A3(\us02\/_0084_ ), .B1(\us02\/_0139_ ), .Y(\us02\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0957_ ( .A(\us02\/_0096_ ), .B(\us02\/_0730_ ), .X(\us02\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0959_ ( .A(\us02\/_0142_ ), .X(\us02\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_0960_ ( .A1(\us02\/_0020_ ), .A2(\us02\/_0144_ ), .A3(\us02\/_0017_ ), .B1(\us02\/_0139_ ), .Y(\us02\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \us02/_0961_ ( .A(\sa02\[2\] ), .B(\us02\/_0050_ ), .C_N(\sa02\[3\] ), .Y(\us02\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0962_ ( .A(\us02\/_0128_ ), .X(\us02\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_0963_ ( .A1(\us02\/_0146_ ), .A2(\us02\/_0032_ ), .A3(\us02\/_0640_ ), .B1(\us02\/_0147_ ), .Y(\us02\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us02/_0964_ ( .A(\us02\/_0136_ ), .B(\us02\/_0141_ ), .C(\us02\/_0145_ ), .D(\us02\/_0148_ ), .X(\us02\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0965_ ( .A(\us02\/_0123_ ), .B(\us02\/_0151_ ), .X(\us02\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0967_ ( .A(\us02\/_0150_ ), .X(\us02\/_0153_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0968_ ( .A(\us02\/_0150_ ), .B(\us02\/_0062_ ), .X(\us02\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_0969_ ( .A(\us02\/_0079_ ), .B(\us02\/_0150_ ), .Y(\us02\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us02/_0970_ ( .A(\us02\/_0150_ ), .B(\us02\/_0412_ ), .C(\us02\/_0249_ ), .Y(\us02\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_0971_ ( .A(\us02\/_0155_ ), .B(\us02\/_0156_ ), .Y(\us02\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_0972_ ( .A1(\us02\/_0153_ ), .A2(\us02\/_0134_ ), .B1(\us02\/_0154_ ), .C1(\us02\/_0157_ ), .Y(\us02\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0973_ ( .A(\us02\/_0467_ ), .B(\us02\/_0123_ ), .X(\us02\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_0975_ ( .A(\us02\/_0159_ ), .X(\us02\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us02/_0976_ ( .A_N(\us02\/_0119_ ), .B(\us02\/_0161_ ), .X(\us02\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us02/_0977_ ( .A(\us02\/_0163_ ), .Y(\us02\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_0978_ ( .A1(\us02\/_0146_ ), .A2(\us02\/_0575_ ), .A3(\us02\/_0608_ ), .B1(\us02\/_0153_ ), .Y(\us02\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_0979_ ( .A1(\us02\/_0062_ ), .A2(\us02\/_0084_ ), .A3(\us02\/_0134_ ), .B1(\us02\/_0161_ ), .Y(\us02\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us02/_0980_ ( .A(\us02\/_0158_ ), .B(\us02\/_0164_ ), .C(\us02\/_0165_ ), .D(\us02\/_0166_ ), .X(\us02\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us02/_0981_ ( .A(\us02\/_0097_ ), .B(\us02\/_0122_ ), .C(\us02\/_0149_ ), .D(\us02\/_0167_ ), .X(\us02\/_0168_ ) );
sky130_fd_sc_hd__and2_1 \us02/_0982_ ( .A(\us02\/_0662_ ), .B(\us02\/_0150_ ), .X(\us02\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_0983_ ( .A(\us02\/_0154_ ), .B(\us02\/_0169_ ), .Y(\us02\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us02/_0984_ ( .A(\us02\/_0123_ ), .B(\us02\/_0151_ ), .C(\us02\/_0038_ ), .X(\us02\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0985_ ( .A(\us02\/_0170_ ), .B(\us02\/_0171_ ), .X(\us02\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \us02/_0986_ ( .A(\us02\/_0172_ ), .Y(\us02\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \us02/_0987_ ( .A(\us02\/_0067_ ), .B(\us02\/_0168_ ), .C(\us02\/_0174_ ), .Y(\us02\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us02/_0988_ ( .A(\sa02\[1\] ), .B(\sa02\[0\] ), .Y(\us02\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us02/_0989_ ( .A(\us02\/_0175_ ), .B(\us02\/_0358_ ), .X(\us02\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0990_ ( .A(\us02\/_0176_ ), .B(\us02\/_0478_ ), .X(\us02\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_0991_ ( .A(\us02\/_0084_ ), .B(\us02\/_0113_ ), .Y(\us02\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0992_ ( .A(\us02\/_0111_ ), .B(\us02\/_0062_ ), .X(\us02\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0993_ ( .A(\us02\/_0111_ ), .B(\us02\/_0662_ ), .X(\us02\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_0994_ ( .A(\us02\/_0179_ ), .B(\us02\/_0180_ ), .Y(\us02\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0995_ ( .A(\us02\/_0054_ ), .B(\us02\/_0058_ ), .X(\us02\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us02/_0996_ ( .A(\us02\/_0182_ ), .Y(\us02\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us02/_0997_ ( .A_N(\us02\/_0177_ ), .B(\us02\/_0178_ ), .C(\us02\/_0181_ ), .D(\us02\/_0184_ ), .X(\us02\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0998_ ( .A(\us02\/_0098_ ), .B(\us02\/_0741_ ), .X(\us02\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us02/_0999_ ( .A(\us02\/_0047_ ), .B(\us02\/_0098_ ), .X(\us02\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us02/_1000_ ( .A(\us02\/_0186_ ), .B(\us02\/_0187_ ), .X(\us02\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1001_ ( .A(\us02\/_0188_ ), .Y(\us02\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1002_ ( .A(\us02\/_0738_ ), .B(\us02\/_0735_ ), .X(\us02\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1003_ ( .A(\us02\/_0271_ ), .B(\us02\/_0736_ ), .X(\us02\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_1004_ ( .A(\us02\/_0190_ ), .B(\us02\/_0191_ ), .Y(\us02\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us02/_1005_ ( .A(\us02\/_0096_ ), .B(\us02\/_0325_ ), .X(\us02\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1006_ ( .A1(\us02\/_0193_ ), .A2(\us02\/_0176_ ), .B1(\us02\/_0043_ ), .Y(\us02\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1007_ ( .A(\us02\/_0185_ ), .B(\us02\/_0189_ ), .C(\us02\/_0192_ ), .D(\us02\/_0195_ ), .X(\us02\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us02/_1008_ ( .A_N(\sa02\[3\] ), .B(\us02\/_0734_ ), .C(\sa02\[2\] ), .X(\us02\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1009_ ( .A(\us02\/_0137_ ), .B(\us02\/_0197_ ), .X(\us02\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_1010_ ( .A(\us02\/_0198_ ), .B(\us02\/_0040_ ), .Y(\us02\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1011_ ( .A(\us02\/_0293_ ), .B(\us02\/_0137_ ), .X(\us02\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1012_ ( .A(\us02\/_0200_ ), .Y(\us02\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1013_ ( .A(\us02\/_0137_ ), .B(\us02\/_0110_ ), .Y(\us02\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1014_ ( .A(\us02\/_0139_ ), .B(\us02\/_0020_ ), .Y(\us02\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1015_ ( .A(\us02\/_0199_ ), .B(\us02\/_0201_ ), .C(\us02\/_0202_ ), .D(\us02\/_0203_ ), .X(\us02\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us02/_1016_ ( .A1(\us02\/_0532_ ), .A2(\us02\/_0109_ ), .B1(\us02\/_0102_ ), .C1(\us02\/_0727_ ), .X(\us02\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1017_ ( .A(\us02\/_0022_ ), .B(\us02\/_0078_ ), .Y(\us02\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1018_ ( .A(\us02\/_0078_ ), .B(\us02\/_0142_ ), .Y(\us02\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1019_ ( .A(\us02\/_0207_ ), .B(\us02\/_0208_ ), .Y(\us02\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1020_ ( .A1(\us02\/_0094_ ), .A2(\us02\/_0176_ ), .B1(\us02\/_0206_ ), .C1(\us02\/_0209_ ), .Y(\us02\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1021_ ( .A(\us02\/_0662_ ), .B(\us02\/_0070_ ), .X(\us02\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us02/_1022_ ( .A(\us02\/_0731_ ), .B(\us02\/_0123_ ), .C(\us02\/_0749_ ), .Y(\us02\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us02/_1023_ ( .A(\us02\/_0731_ ), .B(\us02\/_0467_ ), .C(\us02\/_0069_ ), .Y(\us02\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us02/_1024_ ( .A_N(\us02\/_0211_ ), .B(\us02\/_0127_ ), .C(\us02\/_0212_ ), .D(\us02\/_0213_ ), .X(\us02\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1025_ ( .A(\us02\/_0137_ ), .Y(\us02\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1026_ ( .A(\us02\/_0128_ ), .B(\us02\/_0035_ ), .Y(\us02\/_0217_ ) );
sky130_fd_sc_hd__buf_2 \us02/_1027_ ( .A(\us02\/_0478_ ), .X(\us02\/_0218_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1028_ ( .A1(\us02\/_0159_ ), .A2(\us02\/_0746_ ), .B1(\us02\/_0434_ ), .B2(\us02\/_0218_ ), .Y(\us02\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us02/_1029_ ( .A1(\us02\/_0116_ ), .A2(\us02\/_0215_ ), .B1(\us02\/_0217_ ), .C1(\us02\/_0219_ ), .X(\us02\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1030_ ( .A(\us02\/_0113_ ), .B(\us02\/_0746_ ), .X(\us02\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us02/_1031_ ( .A1(\us02\/_0098_ ), .A2(\us02\/_0746_ ), .B1(\us02\/_0434_ ), .B2(\us02\/_0750_ ), .X(\us02\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1032_ ( .A1(\us02\/_0047_ ), .A2(\us02\/_0113_ ), .B1(\us02\/_0221_ ), .C1(\us02\/_0222_ ), .Y(\us02\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us02/_1033_ ( .A1(\us02\/_0129_ ), .A2(\us02\/_0162_ ), .B1(\us02\/_0271_ ), .B2(\us02\/_0705_ ), .X(\us02\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1034_ ( .A1(\us02\/_0093_ ), .A2(\us02\/_0738_ ), .B1(\us02\/_0081_ ), .C1(\us02\/_0224_ ), .Y(\us02\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1035_ ( .A(\us02\/_0214_ ), .B(\us02\/_0220_ ), .C(\us02\/_0223_ ), .D(\us02\/_0225_ ), .X(\us02\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1036_ ( .A(\us02\/_0196_ ), .B(\us02\/_0204_ ), .C(\us02\/_0210_ ), .D(\us02\/_0226_ ), .X(\us02\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1037_ ( .A(\us02\/_0111_ ), .B(\us02\/_0554_ ), .X(\us02\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1038_ ( .A(\us02\/_0229_ ), .Y(\us02\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1039_ ( .A(\us02\/_0111_ ), .B(\us02\/_0129_ ), .Y(\us02\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1040_ ( .A(\us02\/_0017_ ), .B(\us02\/_0738_ ), .Y(\us02\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1041_ ( .A(\us02\/_0030_ ), .B(\us02\/_0304_ ), .Y(\us02\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1042_ ( .A(\us02\/_0230_ ), .B(\us02\/_0231_ ), .C(\us02\/_0232_ ), .D(\us02\/_0233_ ), .X(\us02\/_0234_ ) );
sky130_fd_sc_hd__and2_1 \us02/_1043_ ( .A(\us02\/_0047_ ), .B(\us02\/_0478_ ), .X(\us02\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1044_ ( .A1(\us02\/_0129_ ), .A2(\us02\/_0554_ ), .B1(\us02\/_0137_ ), .Y(\us02\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us02/_1045_ ( .A(\us02\/_0235_ ), .B(\us02\/_0049_ ), .C_N(\us02\/_0236_ ), .Y(\us02\/_0237_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1046_ ( .A(\us02\/_0047_ ), .B(\us02\/_0077_ ), .X(\us02\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1047_ ( .A(\us02\/_0070_ ), .B(\us02\/_0035_ ), .X(\us02\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us02/_1048_ ( .A1(\us02\/_0047_ ), .A2(\us02\/_0736_ ), .B1(\us02\/_0022_ ), .B2(\us02\/_0099_ ), .X(\us02\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us02/_1049_ ( .A(\us02\/_0239_ ), .B(\us02\/_0240_ ), .C(\us02\/_0241_ ), .Y(\us02\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1050_ ( .A(\us02\/_0554_ ), .B(\us02\/_0072_ ), .X(\us02\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us02/_1051_ ( .A1(\us02\/_0142_ ), .A2(\us02\/_0137_ ), .B1(\us02\/_0159_ ), .B2(\us02\/_0082_ ), .X(\us02\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1052_ ( .A1(\us02\/_0608_ ), .A2(\us02\/_0072_ ), .B1(\us02\/_0243_ ), .C1(\us02\/_0244_ ), .Y(\us02\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1053_ ( .A(\us02\/_0234_ ), .B(\us02\/_0237_ ), .C(\us02\/_0242_ ), .D(\us02\/_0245_ ), .X(\us02\/_0246_ ) );
sky130_fd_sc_hd__buf_2 \us02/_1054_ ( .A(\us02\/_0027_ ), .X(\us02\/_0247_ ) );
sky130_fd_sc_hd__o21a_1 \us02/_1055_ ( .A1(\us02\/_0554_ ), .A2(\us02\/_0586_ ), .B1(\us02\/_0247_ ), .X(\us02\/_0248_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1056_ ( .A(\us02\/_0082_ ), .B(\us02\/_0478_ ), .X(\us02\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_1057_ ( .A(\us02\/_0079_ ), .X(\us02\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1058_ ( .A(\us02\/_0251_ ), .B(\us02\/_0478_ ), .X(\us02\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_1059_ ( .A(\us02\/_0250_ ), .B(\us02\/_0252_ ), .Y(\us02\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1060_ ( .A(\us02\/_0016_ ), .B(\us02\/_0064_ ), .Y(\us02\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_1061_ ( .A(\us02\/_0304_ ), .X(\us02\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1062_ ( .A(\us02\/_0255_ ), .B(\us02\/_0640_ ), .Y(\us02\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us02/_1063_ ( .A_N(\us02\/_0248_ ), .B(\us02\/_0253_ ), .C(\us02\/_0254_ ), .D(\us02\/_0256_ ), .X(\us02\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1064_ ( .A(\us02\/_0099_ ), .B(\us02\/_0110_ ), .X(\us02\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us02/_1065_ ( .A1(\us02\/_0161_ ), .A2(\us02\/_0130_ ), .B1(\us02\/_0258_ ), .Y(\us02\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1066_ ( .A(\us02\/_0194_ ), .B(\sa02\[1\] ), .X(\us02\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1068_ ( .A(\us02\/_0261_ ), .B(\us02\/_0153_ ), .Y(\us02\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us02/_1069_ ( .A_N(\us02\/_0154_ ), .B(\us02\/_0259_ ), .C(\us02\/_0263_ ), .X(\us02\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1070_ ( .A(\us02\/_0246_ ), .B(\us02\/_0174_ ), .C(\us02\/_0257_ ), .D(\us02\/_0264_ ), .X(\us02\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us02/_1071_ ( .A1(\us02\/_0261_ ), .A2(\us02\/_0554_ ), .B1(\us02\/_0159_ ), .X(\us02\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1072_ ( .A(\us02\/_0746_ ), .B(\us02\/_0150_ ), .Y(\us02\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1073_ ( .A(\us02\/_0175_ ), .Y(\us02\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us02/_1074_ ( .A(\us02\/_0412_ ), .B(\us02\/_0123_ ), .C(\us02\/_0151_ ), .X(\us02\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1075_ ( .A(\us02\/_0268_ ), .B(\us02\/_0269_ ), .Y(\us02\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us02/_1076_ ( .A_N(\us02\/_0266_ ), .B(\us02\/_0267_ ), .C(\us02\/_0270_ ), .X(\us02\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1077_ ( .A(\us02\/_0554_ ), .B(\us02\/_0150_ ), .X(\us02\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1078_ ( .A(\us02\/_0273_ ), .Y(\us02\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1079_ ( .A1(\us02\/_0734_ ), .A2(\us02\/_0325_ ), .B1(\us02\/_0380_ ), .Y(\us02\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1080_ ( .A(\us02\/_0275_ ), .Y(\us02\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1081_ ( .A(\us02\/_0276_ ), .B(\us02\/_0153_ ), .Y(\us02\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us02/_1082_ ( .A(\us02\/_0272_ ), .B(\us02\/_0274_ ), .C(\us02\/_0277_ ), .X(\us02\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_1083_ ( .A(\us02\/_0035_ ), .X(\us02\/_0279_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1085_ ( .A1(\us02\/_0218_ ), .A2(\us02\/_0279_ ), .B1(\us02\/_0084_ ), .B2(\us02\/_0060_ ), .Y(\us02\/_0281_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1086_ ( .A1(\us02\/_0251_ ), .A2(\us02\/_0434_ ), .B1(\us02\/_0304_ ), .Y(\us02\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1087_ ( .A(\us02\/_0091_ ), .B(\us02\/_0056_ ), .Y(\us02\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1088_ ( .A1(\us02\/_0118_ ), .A2(\us02\/_0050_ ), .B1(\us02\/_0038_ ), .C1(\us02\/_0255_ ), .Y(\us02\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1089_ ( .A(\us02\/_0281_ ), .B(\us02\/_0283_ ), .C(\us02\/_0284_ ), .D(\us02\/_0285_ ), .X(\us02\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1090_ ( .A(\us02\/_0082_ ), .B(\us02\/_0027_ ), .X(\us02\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1091_ ( .A(\us02\/_0129_ ), .B(\us02\/_0027_ ), .X(\us02\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_1092_ ( .A(\us02\/_0287_ ), .B(\us02\/_0288_ ), .Y(\us02\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1093_ ( .A1(\us02\/_0752_ ), .A2(\us02\/_0683_ ), .B1(\us02\/_0093_ ), .B2(\us02\/_0247_ ), .Y(\us02\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1094_ ( .A1(\us02\/_0092_ ), .A2(\us02\/_0575_ ), .B1(\us02\/_0056_ ), .Y(\us02\/_0291_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1096_ ( .A1(\us02\/_0218_ ), .A2(\us02\/_0662_ ), .B1(\us02\/_0084_ ), .B2(\us02\/_0056_ ), .Y(\us02\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1097_ ( .A(\us02\/_0289_ ), .B(\us02\/_0290_ ), .C(\us02\/_0291_ ), .D(\us02\/_0294_ ), .X(\us02\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1098_ ( .A(\us02\/_0750_ ), .B(\us02\/_0193_ ), .X(\us02\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1099_ ( .A(\us02\/_0705_ ), .B(\us02\/_0380_ ), .X(\us02\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1100_ ( .A(\us02\/_0752_ ), .B(\us02\/_0129_ ), .Y(\us02\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us02/_1101_ ( .A(\us02\/_0296_ ), .B(\us02\/_0297_ ), .C_N(\us02\/_0298_ ), .Y(\us02\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1102_ ( .A(\us02\/_0089_ ), .B(\us02\/_0532_ ), .Y(\us02\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1103_ ( .A(\sa02\[2\] ), .Y(\us02\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \us02/_1104_ ( .A(\us02\/_0301_ ), .B(\sa02\[3\] ), .C(\us02\/_0118_ ), .Y(\us02\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1105_ ( .A(\us02\/_0072_ ), .B(\us02\/_0302_ ), .X(\us02\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1106_ ( .A(\us02\/_0303_ ), .Y(\us02\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1107_ ( .A(\us02\/_0147_ ), .B(\us02\/_0302_ ), .Y(\us02\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1108_ ( .A(\us02\/_0299_ ), .B(\us02\/_0300_ ), .C(\us02\/_0305_ ), .D(\us02\/_0306_ ), .X(\us02\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1109_ ( .A(\us02\/_0278_ ), .B(\us02\/_0286_ ), .C(\us02\/_0295_ ), .D(\us02\/_0307_ ), .X(\us02\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us02/_1110_ ( .A(\us02\/_0228_ ), .B(\us02\/_0265_ ), .C(\us02\/_0308_ ), .Y(\us02\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1111_ ( .A(\us02\/_0235_ ), .Y(\us02\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1112_ ( .A(\us02\/_0478_ ), .B(\us02\/_0640_ ), .X(\us02\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1113_ ( .A(\us02\/_0310_ ), .Y(\us02\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1114_ ( .A(\us02\/_0022_ ), .B(\us02\/_0218_ ), .Y(\us02\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1115_ ( .A(\us02\/_0218_ ), .B(\us02\/_0032_ ), .Y(\us02\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1116_ ( .A(\us02\/_0309_ ), .B(\us02\/_0311_ ), .C(\us02\/_0312_ ), .D(\us02\/_0313_ ), .X(\us02\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1117_ ( .A(\us02\/_0218_ ), .B(\us02\/_0064_ ), .Y(\us02\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1118_ ( .A(\us02\/_0218_ ), .B(\us02\/_0683_ ), .Y(\us02\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1119_ ( .A(\us02\/_0315_ ), .B(\us02\/_0316_ ), .C(\us02\/_0317_ ), .D(\us02\/_0253_ ), .X(\us02\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1120_ ( .A(\us02\/_0047_ ), .B(\us02\/_0304_ ), .Y(\us02\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1121_ ( .A(\us02\/_0586_ ), .B(\us02\/_0162_ ), .Y(\us02\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1122_ ( .A(\us02\/_0319_ ), .B(\us02\/_0320_ ), .Y(\us02\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_1123_ ( .A(\us02\/_0321_ ), .B(\us02\/_0238_ ), .Y(\us02\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1124_ ( .A(\us02\/_0304_ ), .B(\us02\/_0062_ ), .Y(\us02\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_1125_ ( .A(\us02\/_0251_ ), .X(\us02\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1126_ ( .A1(\us02\/_0324_ ), .A2(\us02\/_0084_ ), .B1(\us02\/_0255_ ), .Y(\us02\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1127_ ( .A1(\us02\/_0050_ ), .A2(\us02\/_0205_ ), .B1(\us02\/_0109_ ), .C1(\us02\/_0255_ ), .Y(\us02\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1128_ ( .A(\us02\/_0322_ ), .B(\us02\/_0323_ ), .C(\us02\/_0326_ ), .D(\us02\/_0327_ ), .X(\us02\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1129_ ( .A1(\us02\/_0733_ ), .A2(\us02\/_0279_ ), .A3(\us02\/_0058_ ), .B1(\us02\/_0056_ ), .Y(\us02\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_1130_ ( .A(\us02\/_0047_ ), .X(\us02\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1131_ ( .A(\us02\/_0330_ ), .B(\us02\/_0056_ ), .Y(\us02\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1132_ ( .A(\us02\/_0054_ ), .B(\us02\/_0045_ ), .Y(\us02\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1133_ ( .A(\us02\/_0329_ ), .B(\us02\/_0331_ ), .C(\us02\/_0284_ ), .D(\us02\/_0332_ ), .X(\us02\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us02/_1134_ ( .A1(\us02\/_0249_ ), .A2(\us02\/_0205_ ), .B1(\us02\/_0532_ ), .C1(\us02\/_0060_ ), .X(\us02\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1135_ ( .A(\us02\/_0084_ ), .B(\us02\/_0060_ ), .Y(\us02\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1136_ ( .A(\us02\/_0324_ ), .B(\us02\/_0060_ ), .Y(\us02\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1137_ ( .A(\us02\/_0335_ ), .B(\us02\/_0337_ ), .Y(\us02\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1138_ ( .A1(\us02\/_0276_ ), .A2(\us02\/_0060_ ), .B1(\us02\/_0334_ ), .C1(\us02\/_0338_ ), .Y(\us02\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1139_ ( .A(\us02\/_0318_ ), .B(\us02\/_0328_ ), .C(\us02\/_0333_ ), .D(\us02\/_0339_ ), .X(\us02\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us02/_1140_ ( .A1(\us02\/_0746_ ), .A2(\us02\/_0134_ ), .B1(\us02\/_0128_ ), .X(\us02\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us02/_1141_ ( .A_N(\us02\/_0086_ ), .B(\us02\/_0128_ ), .X(\us02\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1142_ ( .A(\us02\/_0079_ ), .B(\us02\/_0124_ ), .X(\us02\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_1143_ ( .A(\us02\/_0126_ ), .B(\us02\/_0343_ ), .Y(\us02\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us02/_1144_ ( .A(\us02\/_0341_ ), .B(\us02\/_0342_ ), .C_N(\us02\/_0344_ ), .Y(\us02\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1146_ ( .A1(\us02\/_0193_ ), .A2(\us02\/_0092_ ), .A3(\us02\/_0330_ ), .B1(\us02\/_0147_ ), .Y(\us02\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1147_ ( .A1(\us02\/_0130_ ), .A2(\us02\/_0084_ ), .A3(\us02\/_0134_ ), .B1(\us02\/_0139_ ), .Y(\us02\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1148_ ( .A1(\us02\/_0144_ ), .A2(\us02\/_0608_ ), .A3(\us02\/_0092_ ), .B1(\us02\/_0139_ ), .Y(\us02\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1149_ ( .A(\us02\/_0345_ ), .B(\us02\/_0348_ ), .C(\us02\/_0349_ ), .D(\us02\/_0350_ ), .X(\us02\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us02/_1150_ ( .A(\us02\/_0150_ ), .B(\us02\/_0194_ ), .C(\us02\/_0249_ ), .X(\us02\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us02/_1151_ ( .A(\us02\/_0277_ ), .SLEEP(\us02\/_0352_ ), .X(\us02\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us02/_1152_ ( .A1(\us02\/_0268_ ), .A2(\us02\/_0171_ ), .B1(\us02\/_0157_ ), .Y(\us02\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us02/_1153_ ( .A(\us02\/_0161_ ), .X(\us02\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1154_ ( .A1(\us02\/_0279_ ), .A2(\us02\/_0084_ ), .B1(\us02\/_0355_ ), .Y(\us02\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1155_ ( .A1(\us02\/_0020_ ), .A2(\us02\/_0193_ ), .A3(\us02\/_0091_ ), .B1(\us02\/_0355_ ), .Y(\us02\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1156_ ( .A(\us02\/_0353_ ), .B(\us02\/_0354_ ), .C(\us02\/_0356_ ), .D(\us02\/_0357_ ), .X(\us02\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1157_ ( .A(\us02\/_0111_ ), .B(\us02\/_0586_ ), .X(\us02\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1158_ ( .A(\us02\/_0360_ ), .Y(\us02\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us02/_1159_ ( .A1(\us02\/_0119_ ), .A2(\us02\/_0120_ ), .B1(\us02\/_0230_ ), .C1(\us02\/_0361_ ), .X(\us02\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1160_ ( .A1(\us02\/_0662_ ), .A2(\us02\/_0251_ ), .A3(\us02\/_0134_ ), .B1(\us02\/_0114_ ), .Y(\us02\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1162_ ( .A1(\us02\/_0035_ ), .A2(\us02\/_0251_ ), .A3(\us02\/_0134_ ), .B1(\us02\/_0099_ ), .Y(\us02\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1163_ ( .A1(\us02\/_0193_ ), .A2(\us02\/_0608_ ), .B1(\us02\/_0099_ ), .Y(\us02\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1164_ ( .A(\us02\/_0362_ ), .B(\us02\/_0363_ ), .C(\us02\/_0365_ ), .D(\us02\/_0366_ ), .X(\us02\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1165_ ( .A1(\us02\/_0575_ ), .A2(\us02\/_0092_ ), .A3(\us02\/_0330_ ), .B1(\us02\/_0089_ ), .Y(\us02\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1166_ ( .A1(\us02\/_0586_ ), .A2(\us02\/_0017_ ), .A3(\us02\/_0330_ ), .B1(\us02\/_0094_ ), .Y(\us02\/_0370_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1167_ ( .A1(\us02\/_0293_ ), .A2(\us02\/_0134_ ), .B1(\us02\/_0089_ ), .Y(\us02\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1168_ ( .A1(\us02\/_0279_ ), .A2(\us02\/_0134_ ), .B1(\us02\/_0094_ ), .Y(\us02\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1169_ ( .A(\us02\/_0368_ ), .B(\us02\/_0370_ ), .C(\us02\/_0371_ ), .D(\us02\/_0372_ ), .X(\us02\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1170_ ( .A(\us02\/_0351_ ), .B(\us02\/_0359_ ), .C(\us02\/_0367_ ), .D(\us02\/_0373_ ), .X(\us02\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1171_ ( .A1(\us02\/_0102_ ), .A2(\us02\/_0347_ ), .B1(\us02\/_0109_ ), .C1(\us02\/_0247_ ), .Y(\us02\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1172_ ( .A1(\us02\/_0102_ ), .A2(\us02\/_0347_ ), .B1(\us02\/_0532_ ), .C1(\us02\/_0247_ ), .Y(\us02\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1173_ ( .A1(\us02\/_0050_ ), .A2(\us02\/_0249_ ), .B1(\us02\/_0380_ ), .C1(\us02\/_0247_ ), .Y(\us02\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1174_ ( .A(\us02\/_0041_ ), .B(\us02\/_0375_ ), .C(\us02\/_0376_ ), .D(\us02\/_0377_ ), .X(\us02\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1175_ ( .A(\us02\/_0047_ ), .B(\us02\/_0750_ ), .X(\us02\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1176_ ( .A(\us02\/_0379_ ), .Y(\us02\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1177_ ( .A(\us02\/_0016_ ), .B(\us02\/_0608_ ), .Y(\us02\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1178_ ( .A(\us02\/_0752_ ), .B(\us02\/_0554_ ), .Y(\us02\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1179_ ( .A1(\sa02\[1\] ), .A2(\us02\/_0734_ ), .B1(\us02\/_0109_ ), .C1(\us02\/_0016_ ), .Y(\us02\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1180_ ( .A(\us02\/_0381_ ), .B(\us02\/_0382_ ), .C(\us02\/_0383_ ), .D(\us02\/_0384_ ), .X(\us02\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us02/_1181_ ( .A(\us02\/_0086_ ), .B_N(\us02\/_0736_ ), .X(\us02\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1182_ ( .A1(\us02\/_0748_ ), .A2(\us02\/_0134_ ), .B1(\us02\/_0739_ ), .Y(\us02\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1183_ ( .A1(\us02\/_0118_ ), .A2(\us02\/_0249_ ), .B1(\us02\/_0109_ ), .C1(\us02\/_0739_ ), .Y(\us02\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1184_ ( .A1(\us02\/_0102_ ), .A2(\us02\/_0301_ ), .B1(\sa02\[3\] ), .C1(\us02\/_0739_ ), .Y(\us02\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1185_ ( .A(\us02\/_0386_ ), .B(\us02\/_0387_ ), .C(\us02\/_0388_ ), .D(\us02\/_0389_ ), .X(\us02\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1186_ ( .A(\us02\/_0020_ ), .Y(\us02\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1187_ ( .A(\us02\/_0727_ ), .Y(\us02\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1188_ ( .A(\us02\/_0727_ ), .B(\us02\/_0064_ ), .Y(\us02\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1189_ ( .A1(\us02\/_0102_ ), .A2(\us02\/_0734_ ), .B1(\us02\/_0532_ ), .C1(\us02\/_0727_ ), .Y(\us02\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us02/_1190_ ( .A1(\us02\/_0392_ ), .A2(\us02\/_0393_ ), .B1(\us02\/_0394_ ), .C1(\us02\/_0395_ ), .X(\us02\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1191_ ( .A(\us02\/_0378_ ), .B(\us02\/_0385_ ), .C(\us02\/_0390_ ), .D(\us02\/_0396_ ), .X(\us02\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us02/_1192_ ( .A(\us02\/_0340_ ), .B(\us02\/_0374_ ), .C(\us02\/_0397_ ), .Y(\us02\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1193_ ( .A(\us02\/_0077_ ), .B(\us02\/_0129_ ), .X(\us02\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_1194_ ( .A(\us02\/_0398_ ), .B(\us02\/_0239_ ), .Y(\us02\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1195_ ( .A(\us02\/_0022_ ), .B(\us02\/_0111_ ), .X(\us02\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us02/_1196_ ( .A_N(\us02\/_0400_ ), .B(\us02\/_0231_ ), .Y(\us02\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us02/_1197_ ( .A(\us02\/_0399_ ), .SLEEP(\us02\/_0402_ ), .X(\us02\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_1198_ ( .A(\us02\/_0746_ ), .B(\us02\/_0251_ ), .Y(\us02\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us02/_1199_ ( .A_N(\us02\/_0404_ ), .B(\us02\/_0752_ ), .Y(\us02\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us02/_1200_ ( .A(\us02\/_0467_ ), .B(\us02\/_0194_ ), .C(\us02\/_0694_ ), .X(\us02\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us02/_1201_ ( .A_N(\us02\/_0175_ ), .B(\us02\/_0406_ ), .X(\us02\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1202_ ( .A(\us02\/_0407_ ), .Y(\us02\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1203_ ( .A1(\us02\/_0094_ ), .A2(\us02\/_0197_ ), .B1(\us02\/_0114_ ), .B2(\us02\/_0640_ ), .Y(\us02\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1204_ ( .A(\us02\/_0403_ ), .B(\us02\/_0405_ ), .C(\us02\/_0408_ ), .D(\us02\/_0409_ ), .X(\us02\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1205_ ( .A(\us02\/_0030_ ), .B(\us02\/_0150_ ), .Y(\us02\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us02/_1206_ ( .A_N(\us02\/_0169_ ), .B(\us02\/_0289_ ), .C(\us02\/_0411_ ), .X(\us02\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us02/_1207_ ( .A1(\us02\/_0467_ ), .A2(\us02\/_0151_ ), .B1(\us02\/_0140_ ), .C1(\us02\/_0129_ ), .X(\us02\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1208_ ( .A1(\us02\/_0608_ ), .A2(\us02\/_0099_ ), .B1(\us02\/_0037_ ), .C1(\us02\/_0414_ ), .Y(\us02\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1209_ ( .A(\us02\/_0738_ ), .Y(\us02\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1210_ ( .A(\us02\/_0586_ ), .B(\us02\/_0736_ ), .Y(\us02\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1211_ ( .A1(\us02\/_0194_ ), .A2(\us02\/_0038_ ), .B1(\us02\/_0118_ ), .C1(\us02\/_0153_ ), .Y(\us02\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us02/_1212_ ( .A1(\us02\/_0416_ ), .A2(\us02\/_0117_ ), .B1(\us02\/_0417_ ), .C1(\us02\/_0418_ ), .X(\us02\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1213_ ( .A(\us02\/_0077_ ), .B(\us02\/_0035_ ), .X(\us02\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1214_ ( .A(\us02\/_0662_ ), .B(\us02\/_0124_ ), .Y(\us02\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1215_ ( .A(\us02\/_0030_ ), .B(\us02\/_0137_ ), .Y(\us02\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1216_ ( .A(\us02\/_0072_ ), .B(\us02\/_0731_ ), .Y(\us02\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us02/_1217_ ( .A_N(\us02\/_0420_ ), .B(\us02\/_0421_ ), .C(\us02\/_0422_ ), .D(\us02\/_0424_ ), .X(\us02\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1218_ ( .A(\us02\/_0413_ ), .B(\us02\/_0415_ ), .C(\us02\/_0419_ ), .D(\us02\/_0425_ ), .X(\us02\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us02/_1219_ ( .A(\us02\/_0355_ ), .B(\us02\/_0102_ ), .C(\us02\/_0109_ ), .Y(\us02\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1220_ ( .A(\us02\/_0077_ ), .B(\us02\/_0017_ ), .X(\us02\/_0428_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1221_ ( .A(\us02\/_0077_ ), .B(\us02\/_0554_ ), .X(\us02\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us02/_1222_ ( .A1(\us02\/_0050_ ), .A2(\us02\/_0205_ ), .B1(\us02\/_0380_ ), .C1(\us02\/_0078_ ), .X(\us02\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us02/_1223_ ( .A(\us02\/_0428_ ), .B(\us02\/_0429_ ), .C(\us02\/_0430_ ), .Y(\us02\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us02/_1224_ ( .A_N(\us02\/_0209_ ), .B(\us02\/_0431_ ), .X(\us02\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us02/_1225_ ( .A1(\us02\/_0215_ ), .A2(\us02\/_0404_ ), .B1(\us02\/_0427_ ), .C1(\us02\/_0432_ ), .X(\us02\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1226_ ( .A(\us02\/_0043_ ), .B(\us02\/_0058_ ), .Y(\us02\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1227_ ( .A(\us02\/_0195_ ), .B(\us02\/_0233_ ), .C(\us02\/_0320_ ), .D(\us02\/_0435_ ), .X(\us02\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1228_ ( .A(\us02\/_0261_ ), .B(\us02\/_0738_ ), .Y(\us02\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1229_ ( .A1(\us02\/_0218_ ), .A2(\us02\/_0640_ ), .B1(\us02\/_0261_ ), .B2(\us02\/_0056_ ), .Y(\us02\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1230_ ( .A(\us02\/_0436_ ), .B(\us02\/_0394_ ), .C(\us02\/_0437_ ), .D(\us02\/_0438_ ), .X(\us02\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1231_ ( .A(\us02\/_0410_ ), .B(\us02\/_0426_ ), .C(\us02\/_0433_ ), .D(\us02\/_0439_ ), .X(\us02\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us02/_1232_ ( .A(\us02\/_0135_ ), .SLEEP(\us02\/_0273_ ), .X(\us02\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1233_ ( .A1(\us02\/_0279_ ), .A2(\us02\/_0134_ ), .B1(\us02\/_0099_ ), .Y(\us02\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1234_ ( .A(\us02\/_0441_ ), .B(\us02\/_0164_ ), .C(\us02\/_0270_ ), .D(\us02\/_0442_ ), .X(\us02\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1235_ ( .A(\us02\/_0051_ ), .B(\us02\/_0662_ ), .Y(\us02\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1236_ ( .A(\us02\/_0051_ ), .B(\us02\/_0271_ ), .Y(\us02\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1237_ ( .A(\us02\/_0444_ ), .B(\us02\/_0446_ ), .X(\us02\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1238_ ( .A(\us02\/_0193_ ), .B(\us02\/_0304_ ), .X(\us02\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1239_ ( .A(\us02\/_0448_ ), .Y(\us02\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1240_ ( .A(\us02\/_0162_ ), .B(\us02\/_0130_ ), .X(\us02\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1241_ ( .A(\us02\/_0450_ ), .Y(\us02\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1242_ ( .A1(\us02\/_0129_ ), .A2(\us02\/_0554_ ), .B1(\us02\/_0043_ ), .Y(\us02\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1243_ ( .A(\us02\/_0447_ ), .B(\us02\/_0449_ ), .C(\us02\/_0451_ ), .D(\us02\/_0452_ ), .X(\us02\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1244_ ( .A(\us02\/_0056_ ), .B(\us02\/_0064_ ), .Y(\us02\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us02/_1245_ ( .A_N(\us02\/_0248_ ), .B(\us02\/_0454_ ), .C(\us02\/_0254_ ), .D(\us02\/_0256_ ), .X(\us02\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1246_ ( .A1(\us02\/_0330_ ), .A2(\us02\/_0099_ ), .B1(\us02\/_0134_ ), .B2(\us02\/_0705_ ), .Y(\us02\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1247_ ( .A1(\us02\/_0748_ ), .A2(\us02\/_0738_ ), .B1(\us02\/_0092_ ), .B2(\us02\/_0752_ ), .Y(\us02\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1248_ ( .A1(\us02\/_0072_ ), .A2(\us02\/_0035_ ), .B1(\us02\/_0748_ ), .B2(\us02\/_0056_ ), .Y(\us02\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1249_ ( .A1(\us02\/_0748_ ), .A2(\us02\/_0251_ ), .B1(\us02\/_0247_ ), .Y(\us02\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1250_ ( .A(\us02\/_0457_ ), .B(\us02\/_0458_ ), .C(\us02\/_0459_ ), .D(\us02\/_0460_ ), .X(\us02\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1251_ ( .A(\us02\/_0443_ ), .B(\us02\/_0453_ ), .C(\us02\/_0455_ ), .D(\us02\/_0461_ ), .X(\us02\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1252_ ( .A(\us02\/_0705_ ), .B(\us02\/_0079_ ), .X(\us02\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1253_ ( .A(\us02\/_0586_ ), .B(\us02\/_0124_ ), .Y(\us02\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1254_ ( .A(\us02\/_0218_ ), .B(\us02\/_0746_ ), .Y(\us02\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us02/_1255_ ( .A_N(\us02\/_0463_ ), .B(\us02\/_0464_ ), .C(\us02\/_0465_ ), .X(\us02\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us02/_1256_ ( .A1(\us02\/_0271_ ), .A2(\us02\/_0072_ ), .B1(\us02\/_0142_ ), .B2(\us02\/_0027_ ), .X(\us02\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1257_ ( .A1(\us02\/_0144_ ), .A2(\us02\/_0099_ ), .B1(\us02\/_0360_ ), .C1(\us02\/_0468_ ), .Y(\us02\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us02/_1258_ ( .A1(\us02\/_0662_ ), .A2(\us02\/_0251_ ), .B1(\us02\/_0218_ ), .X(\us02\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1259_ ( .A1(\us02\/_0575_ ), .A2(\us02\/_0056_ ), .B1(\us02\/_0379_ ), .C1(\us02\/_0470_ ), .Y(\us02\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1260_ ( .A(\us02\/_0466_ ), .B(\us02\/_0469_ ), .C(\us02\/_0471_ ), .D(\us02\/_0305_ ), .X(\us02\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us02/_1261_ ( .A1(\us02\/_0247_ ), .A2(\us02\/_0683_ ), .B1(\us02\/_0324_ ), .B2(\us02\/_0056_ ), .X(\us02\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1262_ ( .A(\us02\/_0084_ ), .B(\us02\/_0099_ ), .X(\us02\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us02/_1263_ ( .A1(\us02\/_0092_ ), .A2(\us02\/_0247_ ), .B1(\us02\/_0474_ ), .X(\us02\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us02/_1264_ ( .A(\us02\/_0075_ ), .B(\us02\/_0473_ ), .C(\us02\/_0475_ ), .Y(\us02\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1265_ ( .A1(\us02\/_0279_ ), .A2(\us02\/_0255_ ), .B1(\us02\/_0084_ ), .B2(\us02\/_0060_ ), .Y(\us02\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1266_ ( .A1(\us02\/_0093_ ), .A2(\us02\/_0056_ ), .B1(\us02\/_0134_ ), .B2(\us02\/_0114_ ), .Y(\us02\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1267_ ( .A1(\us02\/_0161_ ), .A2(\us02\/_0032_ ), .B1(\us02\/_0324_ ), .B2(\us02\/_0147_ ), .Y(\us02\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1268_ ( .A1(\us02\/_0054_ ), .A2(\us02\/_0731_ ), .B1(\us02\/_0748_ ), .B2(\us02\/_0304_ ), .Y(\us02\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1269_ ( .A(\us02\/_0477_ ), .B(\us02\/_0479_ ), .C(\us02\/_0480_ ), .D(\us02\/_0481_ ), .X(\us02\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1270_ ( .A(\us02\/_0161_ ), .B(\us02\/_0064_ ), .Y(\us02\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us02/_1271_ ( .A(\us02\/_0731_ ), .B(\us02\/_0123_ ), .C(\us02\/_0467_ ), .Y(\us02\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1272_ ( .A(\us02\/_0483_ ), .B(\us02\/_0484_ ), .Y(\us02\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1273_ ( .A(\us02\/_0297_ ), .Y(\us02\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us02/_1274_ ( .A_N(\us02\/_0485_ ), .B(\us02\/_0181_ ), .C(\us02\/_0486_ ), .D(\us02\/_0386_ ), .X(\us02\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1275_ ( .A(\us02\/_0472_ ), .B(\us02\/_0476_ ), .C(\us02\/_0482_ ), .D(\us02\/_0487_ ), .X(\us02\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \us02/_1276_ ( .A(\us02\/_0440_ ), .B(\us02\/_0462_ ), .C(\us02\/_0488_ ), .Y(\us02\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1277_ ( .A(\us02\/_0403_ ), .B(\us02\/_0230_ ), .C(\us02\/_0451_ ), .D(\us02\/_0361_ ), .X(\us02\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1278_ ( .A1(\us02\/_0118_ ), .A2(\us02\/_0050_ ), .B1(\us02\/_0109_ ), .C1(\us02\/_0139_ ), .Y(\us02\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1279_ ( .A(\us02\/_0447_ ), .B(\us02\/_0437_ ), .C(\us02\/_0491_ ), .D(\us02\/_0427_ ), .X(\us02\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1280_ ( .A1(\us02\/_0084_ ), .A2(\us02\/_0255_ ), .B1(\us02\/_0608_ ), .B2(\us02\/_0247_ ), .Y(\us02\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1281_ ( .A1(\us02\/_0144_ ), .A2(\us02\/_0147_ ), .B1(\us02\/_0355_ ), .B2(\us02\/_0093_ ), .Y(\us02\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1282_ ( .A1(\us02\/_0705_ ), .A2(\us02\/_0279_ ), .B1(\us02\/_0330_ ), .B2(\us02\/_0247_ ), .Y(\us02\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1283_ ( .A1(\us02\/_0279_ ), .A2(\us02\/_0084_ ), .B1(\us02\/_0114_ ), .Y(\us02\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1284_ ( .A(\us02\/_0493_ ), .B(\us02\/_0494_ ), .C(\us02\/_0495_ ), .D(\us02\/_0496_ ), .X(\us02\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1285_ ( .A1(\us02\/_0134_ ), .A2(\us02\/_0137_ ), .B1(\us02\/_0355_ ), .B2(\us02\/_0575_ ), .Y(\us02\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1286_ ( .A1(\us02\/_0099_ ), .A2(\us02\/_0733_ ), .B1(\us02\/_0093_ ), .B2(\us02\/_0218_ ), .Y(\us02\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1287_ ( .A(\us02\/_0147_ ), .B(\us02\/_0640_ ), .Y(\us02\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1288_ ( .A1(\us02\/_0153_ ), .A2(\us02\/_0056_ ), .B1(\us02\/_0748_ ), .Y(\us02\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1289_ ( .A(\us02\/_0498_ ), .B(\us02\/_0500_ ), .C(\us02\/_0501_ ), .D(\us02\/_0502_ ), .X(\us02\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1290_ ( .A(\us02\/_0490_ ), .B(\us02\/_0492_ ), .C(\us02\/_0497_ ), .D(\us02\/_0503_ ), .X(\us02\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us02/_1291_ ( .A_N(\us02\/_0275_ ), .B(\us02\/_0705_ ), .X(\us02\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1292_ ( .A(\us02\/_0505_ ), .Y(\us02\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1293_ ( .A(\us02\/_0380_ ), .B(\us02\/_0347_ ), .X(\us02\/_0507_ ) );
sky130_fd_sc_hd__o21ai_1 \us02/_1294_ ( .A1(\us02\/_0507_ ), .A2(\us02\/_0093_ ), .B1(\us02\/_0056_ ), .Y(\us02\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1295_ ( .A(\us02\/_0322_ ), .B(\us02\/_0277_ ), .C(\us02\/_0506_ ), .D(\us02\/_0508_ ), .X(\us02\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1296_ ( .A(\us02\/_0084_ ), .B(\us02\/_0705_ ), .X(\us02\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1297_ ( .A1(\us02\/_0733_ ), .A2(\us02\/_0114_ ), .B1(\us02\/_0429_ ), .C1(\us02\/_0511_ ), .Y(\us02\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_1298_ ( .A(\us02\/_0019_ ), .B(\us02\/_0024_ ), .Y(\us02\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1299_ ( .A(\us02\/_0512_ ), .B(\us02\/_0513_ ), .C(\us02\/_0742_ ), .D(\us02\/_0306_ ), .X(\us02\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1300_ ( .A1(\us02\/_0532_ ), .A2(\us02\/_0089_ ), .B1(\us02\/_0154_ ), .C1(\us02\/_0169_ ), .Y(\us02\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us02/_1301_ ( .A1(\us02\/_0749_ ), .A2(\us02\/_0026_ ), .B1(\us02\/_0069_ ), .C1(\us02\/_0032_ ), .X(\us02\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us02/_1302_ ( .A1(\us02\/_0324_ ), .A2(\us02\/_0355_ ), .B1(\us02\/_0330_ ), .B2(\us02\/_0727_ ), .X(\us02\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us02/_1303_ ( .A(\us02\/_0133_ ), .B(\us02\/_0516_ ), .C(\us02\/_0517_ ), .Y(\us02\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1304_ ( .A(\us02\/_0509_ ), .B(\us02\/_0514_ ), .C(\us02\/_0515_ ), .D(\us02\/_0518_ ), .X(\us02\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1305_ ( .A(\us02\/_0746_ ), .B(\us02\/_0072_ ), .Y(\us02\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1306_ ( .A1(\us02\/_0082_ ), .A2(\us02\/_0070_ ), .B1(\us02\/_0043_ ), .B2(\us02\/_0193_ ), .Y(\us02\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1307_ ( .A(\us02\/_0311_ ), .B(\us02\/_0520_ ), .C(\us02\/_0332_ ), .D(\us02\/_0522_ ), .X(\us02\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1308_ ( .A(\us02\/_0129_ ), .B(\us02\/_0218_ ), .X(\us02\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_1309_ ( .A(\us02\/_0235_ ), .B(\us02\/_0524_ ), .Y(\us02\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us02/_1310_ ( .A(\us02\/_0081_ ), .B(\us02\/_0085_ ), .Y(\us02\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1311_ ( .A1(\us02\/_0051_ ), .A2(\us02\/_0045_ ), .B1(\us02\/_0130_ ), .B2(\us02\/_0094_ ), .Y(\us02\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1312_ ( .A(\us02\/_0523_ ), .B(\us02\/_0525_ ), .C(\us02\/_0526_ ), .D(\us02\/_0527_ ), .X(\us02\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us02/_1313_ ( .A_N(\us02\/_0250_ ), .B(\us02\/_0521_ ), .Y(\us02\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1314_ ( .A(\us02\/_0128_ ), .B(\us02\/_0020_ ), .X(\us02\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1315_ ( .A(\us02\/_0530_ ), .Y(\us02\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1316_ ( .A(\us02\/_0099_ ), .B(\us02\/_0058_ ), .X(\us02\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1317_ ( .A(\us02\/_0533_ ), .Y(\us02\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us02/_1318_ ( .A_N(\us02\/_0529_ ), .B(\us02\/_0531_ ), .C(\us02\/_0534_ ), .D(\us02\/_0192_ ), .X(\us02\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1319_ ( .A(\us02\/_0434_ ), .B(\us02\/_0078_ ), .X(\us02\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us02/_1320_ ( .A1(\us02\/_0750_ ), .A2(\us02\/_0079_ ), .B1(\us02\/_0129_ ), .B2(\us02\/_0705_ ), .X(\us02\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1321_ ( .A1(\us02\/_0161_ ), .A2(\us02\/_0032_ ), .B1(\us02\/_0536_ ), .C1(\us02\/_0537_ ), .Y(\us02\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us02/_1322_ ( .A1(\us02\/_0746_ ), .A2(\us02\/_0162_ ), .B1(\us02\/_0079_ ), .B2(\us02\/_0043_ ), .X(\us02\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1323_ ( .A1(\us02\/_0093_ ), .A2(\us02\/_0247_ ), .B1(\us02\/_0240_ ), .C1(\us02\/_0539_ ), .Y(\us02\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1324_ ( .A(\us02\/_0434_ ), .B(\us02\/_0043_ ), .X(\us02\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us02/_1325_ ( .A1(\us02\/_0142_ ), .A2(\us02\/_0150_ ), .B1(\us02\/_0022_ ), .B2(\us02\/_0137_ ), .X(\us02\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1326_ ( .A1(\us02\/_0279_ ), .A2(\us02\/_0051_ ), .B1(\us02\/_0541_ ), .C1(\us02\/_0542_ ), .Y(\us02\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1327_ ( .A(\us02\/_0159_ ), .B(\us02\/_0035_ ), .X(\us02\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us02/_1328_ ( .A1(\us02\/_0271_ ), .A2(\us02\/_0434_ ), .B1(\us02\/_0027_ ), .X(\us02\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1329_ ( .A1(\us02\/_0091_ ), .A2(\us02\/_0128_ ), .B1(\us02\/_0545_ ), .C1(\us02\/_0546_ ), .Y(\us02\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1330_ ( .A(\us02\/_0538_ ), .B(\us02\/_0540_ ), .C(\us02\/_0544_ ), .D(\us02\/_0547_ ), .X(\us02\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1331_ ( .A(\us02\/_0099_ ), .B(\us02\/_0193_ ), .X(\us02\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us02/_1332_ ( .A(\us02\/_0549_ ), .B(\us02\/_0186_ ), .C(\us02\/_0187_ ), .Y(\us02\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1333_ ( .A(\us02\/_0062_ ), .B(\us02\/_0347_ ), .C(\us02\/_0749_ ), .D(\us02\/_0694_ ), .X(\us02\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1334_ ( .A1(\us02\/_0130_ ), .A2(\us02\/_0218_ ), .B1(\us02\/_0551_ ), .C1(\us02\/_0101_ ), .Y(\us02\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1335_ ( .A(\us02\/_0139_ ), .B(\us02\/_0640_ ), .Y(\us02\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1336_ ( .A1(\us02\/_0752_ ), .A2(\us02\/_0662_ ), .B1(\us02\/_0084_ ), .B2(\us02\/_0099_ ), .Y(\us02\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1337_ ( .A(\us02\/_0550_ ), .B(\us02\/_0552_ ), .C(\us02\/_0553_ ), .D(\us02\/_0555_ ), .X(\us02\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1338_ ( .A(\us02\/_0528_ ), .B(\us02\/_0535_ ), .C(\us02\/_0548_ ), .D(\us02\/_0556_ ), .X(\us02\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us02/_1339_ ( .A(\us02\/_0504_ ), .B(\us02\/_0519_ ), .C(\us02\/_0557_ ), .Y(\us02\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1340_ ( .A(\us02\/_0054_ ), .B(\us02\/_0507_ ), .X(\us02\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us02/_1341_ ( .A_N(\us02\/_0558_ ), .B(\us02\/_0408_ ), .C(\us02\/_0451_ ), .D(\us02\/_0452_ ), .X(\us02\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1342_ ( .A(\us02\/_0549_ ), .Y(\us02\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1343_ ( .A(\us02\/_0559_ ), .B(\us02\/_0403_ ), .C(\us02\/_0560_ ), .D(\us02\/_0371_ ), .X(\us02\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1344_ ( .A(\us02\/_0181_ ), .B(\us02\/_0178_ ), .X(\us02\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1345_ ( .A(\us02\/_0562_ ), .B(\us02\/_0552_ ), .C(\us02\/_0553_ ), .D(\us02\/_0555_ ), .X(\us02\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1346_ ( .A(\us02\/_0247_ ), .B(\us02\/_0020_ ), .Y(\us02\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1347_ ( .A(\us02\/_0051_ ), .B(\us02\/_0130_ ), .X(\us02\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1348_ ( .A(\us02\/_0566_ ), .Y(\us02\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1349_ ( .A(\us02\/_0159_ ), .B(\us02\/_0412_ ), .X(\us02\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1350_ ( .A1(\us02\/_0752_ ), .A2(\us02\/_0640_ ), .B1(\us02\/_0568_ ), .B2(\us02\/_0175_ ), .Y(\us02\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1351_ ( .A(\us02\/_0076_ ), .B(\us02\/_0565_ ), .C(\us02\/_0567_ ), .D(\us02\/_0569_ ), .X(\us02\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us02/_1352_ ( .A1(\us02\/_0035_ ), .A2(\us02\/_0142_ ), .B1(\us02\/_0161_ ), .X(\us02\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1353_ ( .A(\us02\/_0099_ ), .B(\us02\/_0662_ ), .Y(\us02\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us02/_1354_ ( .A(\us02\/_0420_ ), .B(\us02\/_0571_ ), .C_N(\us02\/_0572_ ), .Y(\us02\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1355_ ( .A(\us02\/_0051_ ), .B(\us02\/_0746_ ), .Y(\us02\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1356_ ( .A(\us02\/_0574_ ), .B(\us02\/_0319_ ), .C(\us02\/_0320_ ), .D(\us02\/_0411_ ), .X(\us02\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1357_ ( .A(\us02\/_0736_ ), .B(\us02\/_0035_ ), .Y(\us02\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1358_ ( .A(\us02\/_0736_ ), .B(\us02\/_0030_ ), .Y(\us02\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1359_ ( .A(\us02\/_0298_ ), .B(\us02\/_0208_ ), .C(\us02\/_0577_ ), .D(\us02\/_0578_ ), .X(\us02\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1360_ ( .A1(\us02\/_0020_ ), .A2(\us02\/_0137_ ), .B1(\us02\/_0261_ ), .B2(\us02\/_0128_ ), .Y(\us02\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1361_ ( .A(\us02\/_0573_ ), .B(\us02\/_0576_ ), .C(\us02\/_0579_ ), .D(\us02\/_0580_ ), .X(\us02\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1362_ ( .A(\us02\/_0561_ ), .B(\us02\/_0563_ ), .C(\us02\/_0570_ ), .D(\us02\/_0581_ ), .X(\us02\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1363_ ( .A(\us02\/_0128_ ), .B(\us02\/_0193_ ), .X(\us02\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1364_ ( .A(\us02\/_0082_ ), .B(\us02\/_0162_ ), .X(\us02\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us02/_1365_ ( .A(\us02\/_0583_ ), .B(\us02\/_0584_ ), .C_N(\us02\/_0437_ ), .Y(\us02\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us02/_1366_ ( .A(\us02\/_0150_ ), .B(\us02\/_0118_ ), .C(\us02\/_0380_ ), .Y(\us02\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us02/_1367_ ( .A_N(\us02\/_0182_ ), .B(\us02\/_0587_ ), .C(\us02\/_0323_ ), .X(\us02\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1368_ ( .A1(\us02\/_0575_ ), .A2(\us02\/_0153_ ), .B1(\us02\/_0727_ ), .B2(\us02\/_0058_ ), .Y(\us02\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1369_ ( .A1(\us02\/_0218_ ), .A2(\us02\/_0064_ ), .B1(\us02\/_0134_ ), .B2(\us02\/_0255_ ), .Y(\us02\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1370_ ( .A(\us02\/_0585_ ), .B(\us02\/_0588_ ), .C(\us02\/_0589_ ), .D(\us02\/_0590_ ), .X(\us02\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us02/_1371_ ( .A1(\us02\/_0091_ ), .A2(\us02\/_0139_ ), .B1(\us02\/_0250_ ), .Y(\us02\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1372_ ( .A1(\us02\/_0092_ ), .A2(\us02\/_0739_ ), .B1(\us02\/_0324_ ), .B2(\us02\/_0247_ ), .Y(\us02\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1373_ ( .A1(\us02\/_0144_ ), .A2(\us02\/_0153_ ), .B1(\us02\/_0683_ ), .B2(\us02\/_0056_ ), .Y(\us02\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1374_ ( .A1(\us02\/_0091_ ), .A2(\us02\/_0218_ ), .B1(\us02\/_0330_ ), .B2(\us02\/_0056_ ), .Y(\us02\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1375_ ( .A(\us02\/_0592_ ), .B(\us02\/_0593_ ), .C(\us02\/_0594_ ), .D(\us02\/_0595_ ), .X(\us02\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1376_ ( .A(\us02\/_0218_ ), .B(\us02\/_0144_ ), .Y(\us02\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1377_ ( .A(\us02\/_0312_ ), .B(\us02\/_0598_ ), .Y(\us02\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1378_ ( .A(\us02\/_0575_ ), .B(\us02\/_0147_ ), .Y(\us02\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1379_ ( .A1(\us02\/_0293_ ), .A2(\us02\/_0137_ ), .B1(\us02\/_0093_ ), .B2(\us02\/_0739_ ), .Y(\us02\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1380_ ( .A1(\us02\/_0734_ ), .A2(\us02\/_0531_ ), .B1(\us02\/_0600_ ), .C1(\us02\/_0601_ ), .Y(\us02\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1381_ ( .A1(\us02\/_0153_ ), .A2(\us02\/_0261_ ), .B1(\us02\/_0599_ ), .C1(\us02\/_0602_ ), .Y(\us02\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1382_ ( .A(\us02\/_0591_ ), .B(\us02\/_0596_ ), .C(\us02\/_0174_ ), .D(\us02\/_0603_ ), .X(\us02\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1383_ ( .A(\us02\/_0247_ ), .B(\us02\/_0144_ ), .Y(\us02\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1384_ ( .A(\us02\/_0113_ ), .B(\us02\/_0017_ ), .Y(\us02\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1385_ ( .A(\us02\/_0381_ ), .B(\us02\/_0605_ ), .C(\us02\/_0361_ ), .D(\us02\/_0606_ ), .X(\us02\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1386_ ( .A1(\us02\/_0016_ ), .A2(\us02\/_0727_ ), .B1(\us02\/_0733_ ), .Y(\us02\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1387_ ( .A1(\us02\/_0586_ ), .A2(\us02\/_0159_ ), .B1(\us02\/_0082_ ), .B2(\us02\/_0750_ ), .Y(\us02\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1388_ ( .A1(\us02\/_0142_ ), .A2(\us02\/_0162_ ), .B1(\us02\/_0079_ ), .B2(\us02\/_0054_ ), .Y(\us02\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1389_ ( .A(\us02\/_0610_ ), .B(\us02\/_0611_ ), .C(\us02\/_0105_ ), .D(\us02\/_0106_ ), .X(\us02\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1390_ ( .A1(\us02\/_0094_ ), .A2(\us02\/_0302_ ), .B1(\us02\/_0324_ ), .B2(\us02\/_0089_ ), .Y(\us02\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1391_ ( .A(\us02\/_0607_ ), .B(\us02\/_0609_ ), .C(\us02\/_0612_ ), .D(\us02\/_0613_ ), .X(\us02\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1392_ ( .A(\us02\/_0041_ ), .B(\us02\/_0170_ ), .X(\us02\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1393_ ( .A(\us02\/_0554_ ), .B(\us02\/_0027_ ), .X(\us02\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1394_ ( .A(\us02\/_0027_ ), .B(\us02\/_0261_ ), .Y(\us02\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us02/_1395_ ( .A_N(\us02\/_0616_ ), .B(\us02\/_0617_ ), .Y(\us02\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1396_ ( .A1(\us02\/_0147_ ), .A2(\us02\/_0302_ ), .B1(\us02\/_0342_ ), .C1(\us02\/_0618_ ), .Y(\us02\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1397_ ( .A(\us02\/_0614_ ), .B(\us02\/_0272_ ), .C(\us02\/_0615_ ), .D(\us02\/_0620_ ), .X(\us02\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us02/_1398_ ( .A(\us02\/_0582_ ), .B(\us02\/_0604_ ), .C(\us02\/_0621_ ), .Y(\us02\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1399_ ( .A1(\us02\/_0084_ ), .A2(\us02\/_0134_ ), .B1(\us02\/_0089_ ), .Y(\us02\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1400_ ( .A1(\us02\/_0144_ ), .A2(\us02\/_0608_ ), .A3(\us02\/_0330_ ), .B1(\us02\/_0089_ ), .Y(\us02\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1401_ ( .A1(\us02\/_0197_ ), .A2(\us02\/_0130_ ), .A3(\us02\/_0110_ ), .B1(\us02\/_0094_ ), .Y(\us02\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1402_ ( .A(\us02\/_0432_ ), .B(\us02\/_0622_ ), .C(\us02\/_0623_ ), .D(\us02\/_0624_ ), .X(\us02\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us02/_1403_ ( .A1(\us02\/_0554_ ), .A2(\us02\/_0017_ ), .A3(\us02\/_0022_ ), .B1(\us02\/_0161_ ), .X(\us02\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us02/_1404_ ( .A_N(\us02\/_0269_ ), .B(\us02\/_0170_ ), .X(\us02\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1405_ ( .A1(\us02\/_0109_ ), .A2(\us02\/_0064_ ), .A3(\us02\/_0733_ ), .B1(\us02\/_0355_ ), .Y(\us02\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us02/_1406_ ( .A_N(\us02\/_0626_ ), .B(\us02\/_0627_ ), .C(\us02\/_0353_ ), .D(\us02\/_0628_ ), .X(\us02\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1407_ ( .A1(\us02\/_0091_ ), .A2(\us02\/_0110_ ), .A3(\us02\/_0176_ ), .B1(\us02\/_0139_ ), .Y(\us02\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1408_ ( .A1(\us02\/_0020_ ), .A2(\us02\/_0261_ ), .B1(\us02\/_0147_ ), .Y(\us02\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1409_ ( .A(\us02\/_0631_ ), .B(\us02\/_0344_ ), .C(\us02\/_0421_ ), .D(\us02\/_0632_ ), .X(\us02\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us02/_1410_ ( .A1(\us02\/_0325_ ), .A2(\us02\/_0734_ ), .B1(\us02\/_0038_ ), .C1(\us02\/_0113_ ), .X(\us02\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1411_ ( .A1(\us02\/_0134_ ), .A2(\us02\/_0114_ ), .B1(\us02\/_0221_ ), .C1(\us02\/_0634_ ), .Y(\us02\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us02/_1412_ ( .A(\us02\/_0119_ ), .B_N(\us02\/_0111_ ), .Y(\us02\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1413_ ( .A1(\us02\/_0032_ ), .A2(\us02\/_0113_ ), .B1(\us02\/_0636_ ), .C1(\us02\/_0400_ ), .Y(\us02\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1414_ ( .A1(\us02\/_0731_ ), .A2(\us02\/_0293_ ), .A3(\us02\/_0251_ ), .B1(\us02\/_0099_ ), .Y(\us02\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1415_ ( .A(\us02\/_0189_ ), .B(\us02\/_0635_ ), .C(\us02\/_0637_ ), .D(\us02\/_0638_ ), .X(\us02\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1416_ ( .A(\us02\/_0625_ ), .B(\us02\/_0630_ ), .C(\us02\/_0633_ ), .D(\us02\/_0639_ ), .X(\us02\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1417_ ( .A(\us02\/_0746_ ), .B(\us02\/_0738_ ), .X(\us02\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1418_ ( .A(\us02\/_0736_ ), .B(\us02\/_0731_ ), .X(\us02\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us02/_1419_ ( .A_N(\us02\/_0643_ ), .B(\us02\/_0577_ ), .Y(\us02\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1420_ ( .A1(\us02\/_0084_ ), .A2(\us02\/_0739_ ), .B1(\us02\/_0642_ ), .C1(\us02\/_0644_ ), .Y(\us02\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1421_ ( .A1(\us02\/_0050_ ), .A2(\us02\/_0249_ ), .B1(\us02\/_0194_ ), .C1(\us02\/_0738_ ), .Y(\us02\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1422_ ( .A(\us02\/_0646_ ), .B(\us02\/_0232_ ), .C(\us02\/_0417_ ), .D(\us02\/_0578_ ), .X(\us02\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1423_ ( .A1(\us02\/_0064_ ), .A2(\us02\/_0733_ ), .B1(\us02\/_0727_ ), .Y(\us02\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1424_ ( .A1(\us02\/_0193_ ), .A2(\us02\/_0276_ ), .B1(\us02\/_0727_ ), .Y(\us02\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1425_ ( .A(\us02\/_0645_ ), .B(\us02\/_0647_ ), .C(\us02\/_0648_ ), .D(\us02\/_0649_ ), .X(\us02\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1426_ ( .A1(\us02\/_0325_ ), .A2(\us02\/_0734_ ), .B1(\us02\/_0038_ ), .C1(\us02\/_0247_ ), .Y(\us02\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1427_ ( .A1(\us02\/_0249_ ), .A2(\us02\/_0205_ ), .B1(\us02\/_0412_ ), .C1(\us02\/_0247_ ), .Y(\us02\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1428_ ( .A(\us02\/_0652_ ), .B(\us02\/_0653_ ), .X(\us02\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1429_ ( .A1(\us02\/_0733_ ), .A2(\us02\/_0748_ ), .A3(\us02\/_0324_ ), .B1(\us02\/_0016_ ), .Y(\us02\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1430_ ( .A1(\us02\/_0640_ ), .A2(\us02\/_0193_ ), .A3(\us02\/_0091_ ), .B1(\us02\/_0016_ ), .Y(\us02\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1431_ ( .A1(\us02\/_0102_ ), .A2(\us02\/_0301_ ), .B1(\sa02\[3\] ), .C1(\us02\/_0247_ ), .Y(\us02\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1432_ ( .A(\us02\/_0654_ ), .B(\us02\/_0655_ ), .C(\us02\/_0656_ ), .D(\us02\/_0657_ ), .X(\us02\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1433_ ( .A1(\us02\/_0118_ ), .A2(\us02\/_0050_ ), .B1(\us02\/_0038_ ), .C1(\us02\/_0478_ ), .Y(\us02\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us02/_1434_ ( .A_N(\us02\/_0250_ ), .B(\us02\/_0465_ ), .C(\us02\/_0659_ ), .X(\us02\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1435_ ( .A1(\us02\/_0683_ ), .A2(\us02\/_0324_ ), .B1(\us02\/_0255_ ), .Y(\us02\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1436_ ( .A1(\us02\/_0032_ ), .A2(\us02\/_0193_ ), .A3(\us02\/_0047_ ), .B1(\us02\/_0255_ ), .Y(\us02\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1437_ ( .A1(\us02\/_0144_ ), .A2(\us02\/_0586_ ), .A3(\us02\/_0047_ ), .B1(\us02\/_0218_ ), .Y(\us02\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1438_ ( .A(\us02\/_0660_ ), .B(\us02\/_0661_ ), .C(\us02\/_0663_ ), .D(\us02\/_0664_ ), .X(\us02\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1439_ ( .A1(\us02\/_0091_ ), .A2(\us02\/_0276_ ), .B1(\us02\/_0060_ ), .Y(\us02\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1440_ ( .A1(\us02\/_0144_ ), .A2(\us02\/_0608_ ), .B1(\us02\/_0056_ ), .Y(\us02\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1441_ ( .A1(\us02\/_0412_ ), .A2(\us02\/_0038_ ), .B1(\us02\/_0102_ ), .C1(\us02\/_0060_ ), .Y(\us02\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1442_ ( .A1(\sa02\[1\] ), .A2(\us02\/_0734_ ), .B1(\us02\/_0109_ ), .C1(\us02\/_0056_ ), .Y(\us02\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1443_ ( .A(\us02\/_0666_ ), .B(\us02\/_0667_ ), .C(\us02\/_0668_ ), .D(\us02\/_0669_ ), .X(\us02\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1444_ ( .A(\us02\/_0650_ ), .B(\us02\/_0658_ ), .C(\us02\/_0665_ ), .D(\us02\/_0670_ ), .X(\us02\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us02/_1445_ ( .A(\us02\/_0641_ ), .B(\us02\/_0174_ ), .C(\us02\/_0671_ ), .Y(\us02\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us02/_1446_ ( .A(\us02\/_0049_ ), .B(\us02\/_0618_ ), .C_N(\us02\/_0052_ ), .Y(\us02\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us02/_1447_ ( .A(\us02\/_0239_ ), .Y(\us02\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1448_ ( .A(\us02\/_0705_ ), .B(\us02\/_0032_ ), .Y(\us02\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1449_ ( .A1(\us02\/_0054_ ), .A2(\us02\/_0731_ ), .B1(\us02\/_0035_ ), .B2(\us02\/_0705_ ), .Y(\us02\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1450_ ( .A1(\us02\/_0304_ ), .A2(\us02\/_0731_ ), .B1(\us02\/_0047_ ), .B2(\us02\/_0750_ ), .Y(\us02\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1451_ ( .A(\us02\/_0674_ ), .B(\us02\/_0675_ ), .C(\us02\/_0676_ ), .D(\us02\/_0677_ ), .X(\us02\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us02/_1452_ ( .A_N(\us02\/_0584_ ), .B(\us02\/_0283_ ), .X(\us02\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1453_ ( .A(\us02\/_0673_ ), .B(\us02\/_0678_ ), .C(\us02\/_0679_ ), .D(\us02\/_0508_ ), .X(\us02\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1454_ ( .A1(\us02\/_0016_ ), .A2(\us02\/_0733_ ), .B1(\us02\/_0355_ ), .B2(\us02\/_0092_ ), .Y(\us02\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1455_ ( .A(\us02\/_0681_ ), .B(\us02\/_0034_ ), .X(\us02\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us02/_1456_ ( .A1(\us02\/_0330_ ), .A2(\us02\/_0139_ ), .B1(\us02\/_0324_ ), .B2(\us02\/_0089_ ), .X(\us02\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1457_ ( .A1(\us02\/_0146_ ), .A2(\us02\/_0147_ ), .B1(\us02\/_0133_ ), .C1(\us02\/_0684_ ), .Y(\us02\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1458_ ( .A(\us02\/_0113_ ), .B(\us02\/_0251_ ), .Y(\us02\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us02/_1459_ ( .A_N(\us02\/_0463_ ), .B(\us02\/_0686_ ), .C(\us02\/_0383_ ), .D(\us02\/_0464_ ), .X(\us02\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1460_ ( .A1(\us02\/_0051_ ), .A2(\us02\/_0293_ ), .B1(\us02\/_0084_ ), .B2(\us02\/_0705_ ), .Y(\us02\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1461_ ( .A1(\us02\/_0017_ ), .A2(\us02\/_0072_ ), .B1(\us02\/_0134_ ), .B2(\us02\/_0078_ ), .Y(\us02\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1462_ ( .A(\us02\/_0687_ ), .B(\us02\/_0236_ ), .C(\us02\/_0688_ ), .D(\us02\/_0689_ ), .X(\us02\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1463_ ( .A(\us02\/_0680_ ), .B(\us02\/_0682_ ), .C(\us02\/_0685_ ), .D(\us02\/_0690_ ), .X(\us02\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us02/_1464_ ( .A1(\us02\/_0532_ ), .A2(\us02\/_0380_ ), .B1(\us02\/_0102_ ), .C1(\us02\/_0355_ ), .X(\us02\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us02/_1465_ ( .A(\us02\/_0692_ ), .B(\us02\/_0338_ ), .C(\us02\/_0644_ ), .Y(\us02\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1466_ ( .A(\us02\/_0016_ ), .B(\us02\/_0020_ ), .Y(\us02\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1467_ ( .A1(\us02\/_0032_ ), .A2(\us02\/_0137_ ), .B1(\us02\/_0279_ ), .B2(\us02\/_0094_ ), .Y(\us02\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1468_ ( .A1(\us02\/_0575_ ), .A2(\us02\/_0153_ ), .B1(\us02\/_0161_ ), .B2(\us02\/_0293_ ), .Y(\us02\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1469_ ( .A(\us02\/_0259_ ), .B(\us02\/_0695_ ), .C(\us02\/_0696_ ), .D(\us02\/_0697_ ), .X(\us02\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us02/_1470_ ( .A1(\us02\/_0255_ ), .A2(\us02\/_0640_ ), .B1(\us02\/_0016_ ), .B2(\us02\/_0193_ ), .X(\us02\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1471_ ( .A1(\us02\/_0060_ ), .A2(\us02\/_0176_ ), .B1(\us02\/_0699_ ), .C1(\us02\/_0177_ ), .Y(\us02\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1472_ ( .A1(\us02\/_0091_ ), .A2(\us02\/_0218_ ), .B1(\us02\/_0092_ ), .B2(\us02\/_0705_ ), .Y(\us02\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us02/_1473_ ( .A1(\us02\/_0705_ ), .A2(\us02\/_0683_ ), .B1(\us02\/_0093_ ), .B2(\us02\/_0114_ ), .Y(\us02\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us02/_1474_ ( .A1(\us02\/_0683_ ), .A2(\us02\/_0084_ ), .B1(\us02\/_0094_ ), .Y(\us02\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us02/_1475_ ( .A1(\us02\/_0249_ ), .A2(\us02\/_0205_ ), .B1(\us02\/_0038_ ), .C1(\us02\/_0056_ ), .Y(\us02\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1476_ ( .A(\us02\/_0701_ ), .B(\us02\/_0702_ ), .C(\us02\/_0703_ ), .D(\us02\/_0704_ ), .X(\us02\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1477_ ( .A(\us02\/_0693_ ), .B(\us02\/_0698_ ), .C(\us02\/_0700_ ), .D(\us02\/_0706_ ), .X(\us02\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us02/_1478_ ( .A1(\us02\/_0113_ ), .A2(\us02\/_0640_ ), .B1(\us02\/_0099_ ), .B2(\us02\/_0058_ ), .X(\us02\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us02/_1479_ ( .A(\us02\/_0407_ ), .B(\us02\/_0708_ ), .C(\us02\/_0529_ ), .Y(\us02\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1480_ ( .A(\us02\/_0568_ ), .B(\us02\/_0175_ ), .Y(\us02\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us02/_1481_ ( .A1(\us02\/_0247_ ), .A2(\us02\/_0114_ ), .A3(\us02\/_0051_ ), .B1(\us02\/_0130_ ), .Y(\us02\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1482_ ( .A(\us02\/_0709_ ), .B(\us02\/_0550_ ), .C(\us02\/_0710_ ), .D(\us02\/_0711_ ), .X(\us02\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us02/_1483_ ( .A1(\us02\/_0114_ ), .A2(\us02\/_0064_ ), .B1(\us02\/_0261_ ), .B2(\us02\/_0089_ ), .X(\us02\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1484_ ( .A1(\us02\/_0355_ ), .A2(\us02\/_0261_ ), .B1(\us02\/_0198_ ), .C1(\us02\/_0713_ ), .Y(\us02\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1485_ ( .A(\us02\/_0586_ ), .B(\us02\/_0478_ ), .Y(\us02\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us02/_1486_ ( .A_N(\us02\/_0541_ ), .B(\us02\/_0267_ ), .C(\us02\/_0715_ ), .D(\us02\/_0320_ ), .X(\us02\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1487_ ( .A(\us02\/_0586_ ), .B(\us02\/_0070_ ), .Y(\us02\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us02/_1488_ ( .A_N(\us02\/_0211_ ), .B(\us02\/_0155_ ), .C(\us02\/_0202_ ), .D(\us02\/_0718_ ), .X(\us02\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us02/_1489_ ( .A(\us02\/_0150_ ), .B(\us02\/_0205_ ), .C(\us02\/_0380_ ), .Y(\us02\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us02/_1490_ ( .A(\us02\/_0411_ ), .B(\us02\/_0720_ ), .X(\us02\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us02/_1491_ ( .A1(\us02\/_0017_ ), .A2(\us02\/_0022_ ), .B1(\us02\/_0078_ ), .X(\us02\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us02/_1492_ ( .A1(\us02\/_0134_ ), .A2(\us02\/_0738_ ), .B1(\us02\/_0101_ ), .C1(\us02\/_0722_ ), .Y(\us02\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1493_ ( .A(\us02\/_0717_ ), .B(\us02\/_0719_ ), .C(\us02\/_0721_ ), .D(\us02\/_0723_ ), .X(\us02\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us02/_1494_ ( .A(\us02\/_0739_ ), .B(\us02\/_0193_ ), .Y(\us02\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1495_ ( .A(\us02\/_0344_ ), .B(\us02\/_0184_ ), .C(\us02\/_0449_ ), .D(\us02\/_0725_ ), .X(\us02\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us02/_1496_ ( .A(\us02\/_0712_ ), .B(\us02\/_0714_ ), .C(\us02\/_0724_ ), .D(\us02\/_0726_ ), .X(\us02\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \us02/_1497_ ( .A(\us02\/_0691_ ), .B(\us02\/_0707_ ), .C(\us02\/_0728_ ), .Y(\us02\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \us03/_0753_ ( .A(\sa03\[2\] ), .B_N(\sa03\[3\] ), .Y(\us03\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \us03/_0755_ ( .A(\sa03\[1\] ), .B(\sa03\[0\] ), .X(\us03\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us03/_0756_ ( .A(\us03\/_0096_ ), .B(\us03\/_0118_ ), .X(\us03\/_0129_ ) );
sky130_fd_sc_hd__and2_1 \us03/_0757_ ( .A(\sa03\[7\] ), .B(\sa03\[6\] ), .X(\us03\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_0758_ ( .A(\sa03\[4\] ), .B(\sa03\[5\] ), .Y(\us03\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0759_ ( .A(\us03\/_0140_ ), .B(\us03\/_0151_ ), .X(\us03\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0761_ ( .A(\us03\/_0129_ ), .B(\us03\/_0162_ ), .X(\us03\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0762_ ( .A(\us03\/_0096_ ), .X(\us03\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \us03/_0763_ ( .A(\sa03\[1\] ), .B_N(\sa03\[0\] ), .Y(\us03\/_0205_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0764_ ( .A(\us03\/_0205_ ), .X(\us03\/_0216_ ) );
sky130_fd_sc_hd__and3_1 \us03/_0765_ ( .A(\us03\/_0162_ ), .B(\us03\/_0194_ ), .C(\us03\/_0216_ ), .X(\us03\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us03/_0766_ ( .A(\us03\/_0183_ ), .SLEEP(\us03\/_0227_ ), .X(\us03\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \us03/_0767_ ( .A(\sa03\[0\] ), .B_N(\sa03\[1\] ), .Y(\us03\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_0768_ ( .A(\sa03\[2\] ), .B(\sa03\[3\] ), .Y(\us03\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0769_ ( .A(\us03\/_0249_ ), .B(\us03\/_0260_ ), .X(\us03\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0771_ ( .A(\us03\/_0271_ ), .X(\us03\/_0293_ ) );
sky130_fd_sc_hd__buf_2 \us03/_0772_ ( .A(\us03\/_0162_ ), .X(\us03\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_0773_ ( .A(\us03\/_0293_ ), .B(\us03\/_0304_ ), .Y(\us03\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us03/_0774_ ( .A(\sa03\[1\] ), .Y(\us03\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us03/_0776_ ( .A(\sa03\[0\] ), .Y(\us03\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0777_ ( .A(\sa03\[2\] ), .B(\sa03\[3\] ), .X(\us03\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0779_ ( .A(\us03\/_0358_ ), .X(\us03\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_0780_ ( .A1(\us03\/_0325_ ), .A2(\us03\/_0347_ ), .B1(\us03\/_0380_ ), .C1(\us03\/_0304_ ), .Y(\us03\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us03/_0781_ ( .A_N(\us03\/_0238_ ), .B(\us03\/_0314_ ), .C(\us03\/_0391_ ), .X(\us03\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us03/_0782_ ( .A(\sa03\[3\] ), .B_N(\sa03\[2\] ), .Y(\us03\/_0412_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0784_ ( .A(\us03\/_0412_ ), .B(\us03\/_0205_ ), .X(\us03\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \us03/_0787_ ( .A(\sa03\[5\] ), .B_N(\sa03\[4\] ), .Y(\us03\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0788_ ( .A(\us03\/_0467_ ), .B(\us03\/_0140_ ), .X(\us03\/_0478_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0789_ ( .A(\us03\/_0478_ ), .X(\us03\/_0489_ ) );
sky130_fd_sc_hd__buf_2 \us03/_0790_ ( .A(\us03\/_0489_ ), .X(\us03\/_0499_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_0791_ ( .A(\us03\/_0134_ ), .B(\us03\/_0499_ ), .Y(\us03\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_0792_ ( .A(\us03\/_0489_ ), .B(\us03\/_0271_ ), .Y(\us03\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0793_ ( .A(\us03\/_0194_ ), .X(\us03\/_0532_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0794_ ( .A(\us03\/_0249_ ), .X(\us03\/_0543_ ) );
sky130_fd_sc_hd__and2_1 \us03/_0795_ ( .A(\us03\/_0543_ ), .B(\us03\/_0358_ ), .X(\us03\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0797_ ( .A(\us03\/_0554_ ), .X(\us03\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us03/_0798_ ( .A(\us03\/_0216_ ), .B(\us03\/_0358_ ), .X(\us03\/_0586_ ) );
sky130_fd_sc_hd__buf_2 \us03/_0800_ ( .A(\us03\/_0586_ ), .X(\us03\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_0801_ ( .A1(\us03\/_0532_ ), .A2(\us03\/_0575_ ), .A3(\us03\/_0608_ ), .B1(\us03\/_0499_ ), .Y(\us03\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us03/_0802_ ( .A(\us03\/_0401_ ), .B(\us03\/_0510_ ), .C(\us03\/_0521_ ), .D(\us03\/_0619_ ), .X(\us03\/_0629_ ) );
sky130_fd_sc_hd__and2_1 \us03/_0803_ ( .A(\us03\/_0358_ ), .B(\sa03\[1\] ), .X(\us03\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0805_ ( .A(\us03\/_0205_ ), .B(\us03\/_0260_ ), .X(\us03\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0806_ ( .A(\us03\/_0662_ ), .X(\us03\/_0672_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0807_ ( .A(\us03\/_0672_ ), .X(\us03\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us03/_0808_ ( .A(\sa03\[6\] ), .B_N(\sa03\[7\] ), .Y(\us03\/_0694_ ) );
sky130_fd_sc_hd__and2_2 \us03/_0809_ ( .A(\us03\/_0467_ ), .B(\us03\/_0694_ ), .X(\us03\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0811_ ( .A(\us03\/_0705_ ), .X(\us03\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_0812_ ( .A1(\us03\/_0640_ ), .A2(\us03\/_0293_ ), .A3(\us03\/_0683_ ), .B1(\us03\/_0727_ ), .Y(\us03\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_0813_ ( .A(\sa03\[1\] ), .B(\sa03\[0\] ), .Y(\us03\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0814_ ( .A(\us03\/_0730_ ), .B(\us03\/_0260_ ), .X(\us03\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0815_ ( .A(\us03\/_0731_ ), .X(\us03\/_0732_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0816_ ( .A(\us03\/_0732_ ), .X(\us03\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0817_ ( .A(\sa03\[0\] ), .X(\us03\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us03/_0818_ ( .A1(\us03\/_0325_ ), .A2(\us03\/_0734_ ), .B1(\us03\/_0412_ ), .X(\us03\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0819_ ( .A(\us03\/_0694_ ), .B(\us03\/_0151_ ), .X(\us03\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0821_ ( .A(\us03\/_0736_ ), .X(\us03\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0822_ ( .A(\us03\/_0738_ ), .X(\us03\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_0823_ ( .A1(\us03\/_0733_ ), .A2(\us03\/_0735_ ), .A3(\us03\/_0293_ ), .B1(\us03\/_0739_ ), .Y(\us03\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us03/_0824_ ( .A(\us03\/_0730_ ), .B_N(\us03\/_0358_ ), .Y(\us03\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_0825_ ( .A(\us03\/_0741_ ), .B(\us03\/_0739_ ), .Y(\us03\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_0827_ ( .A1(\us03\/_0118_ ), .A2(\us03\/_0216_ ), .B1(\us03\/_0532_ ), .C1(\us03\/_0739_ ), .Y(\us03\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us03/_0828_ ( .A(\us03\/_0729_ ), .B(\us03\/_0740_ ), .C(\us03\/_0742_ ), .D(\us03\/_0744_ ), .X(\us03\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0829_ ( .A(\us03\/_0412_ ), .B(\us03\/_0730_ ), .X(\us03\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0830_ ( .A(\us03\/_0746_ ), .X(\us03\/_0747_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0831_ ( .A(\us03\/_0747_ ), .X(\us03\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us03/_0832_ ( .A(\sa03\[4\] ), .B_N(\sa03\[5\] ), .Y(\us03\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0833_ ( .A(\us03\/_0749_ ), .B(\us03\/_0694_ ), .X(\us03\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0835_ ( .A(\us03\/_0750_ ), .X(\us03\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0836_ ( .A(\us03\/_0752_ ), .X(\us03\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0837_ ( .A(\us03\/_0118_ ), .B(\us03\/_0358_ ), .X(\us03\/_0017_ ) );
sky130_fd_sc_hd__buf_2 \us03/_0838_ ( .A(\us03\/_0017_ ), .X(\us03\/_0018_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0839_ ( .A(\us03\/_0752_ ), .B(\us03\/_0018_ ), .X(\us03\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0840_ ( .A(\us03\/_0358_ ), .B(\us03\/_0325_ ), .X(\us03\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0842_ ( .A(\us03\/_0096_ ), .B(\us03\/_0205_ ), .X(\us03\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \us03/_0844_ ( .A1(\us03\/_0020_ ), .A2(\us03\/_0022_ ), .B1(\us03\/_0752_ ), .X(\us03\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_0845_ ( .A1(\us03\/_0748_ ), .A2(\us03\/_0016_ ), .B1(\us03\/_0019_ ), .C1(\us03\/_0024_ ), .Y(\us03\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \us03/_0846_ ( .A(\sa03\[4\] ), .B(\sa03\[5\] ), .X(\us03\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0847_ ( .A(\us03\/_0694_ ), .B(\us03\/_0026_ ), .X(\us03\/_0027_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0848_ ( .A(\us03\/_0027_ ), .X(\us03\/_0028_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0850_ ( .A(\us03\/_0358_ ), .B(\us03\/_0730_ ), .X(\us03\/_0030_ ) );
sky130_fd_sc_hd__buf_2 \us03/_0852_ ( .A(\us03\/_0030_ ), .X(\us03\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_0853_ ( .A(\us03\/_0247_ ), .B(\us03\/_0032_ ), .Y(\us03\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_0854_ ( .A(\us03\/_0247_ ), .B(\us03\/_0735_ ), .Y(\us03\/_0034_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0855_ ( .A(\us03\/_0118_ ), .B(\us03\/_0260_ ), .X(\us03\/_0035_ ) );
sky130_fd_sc_hd__buf_2 \us03/_0856_ ( .A(\us03\/_0035_ ), .X(\us03\/_0036_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0857_ ( .A(\us03\/_0028_ ), .B(\us03\/_0036_ ), .X(\us03\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0858_ ( .A(\us03\/_0260_ ), .X(\us03\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_0859_ ( .A(\us03\/_0038_ ), .B(\us03\/_0347_ ), .Y(\us03\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us03/_0860_ ( .A_N(\us03\/_0039_ ), .B(\us03\/_0028_ ), .X(\us03\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_0861_ ( .A(\us03\/_0037_ ), .B(\us03\/_0040_ ), .Y(\us03\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us03/_0862_ ( .A(\us03\/_0025_ ), .B(\us03\/_0033_ ), .C(\us03\/_0034_ ), .D(\us03\/_0041_ ), .X(\us03\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0863_ ( .A(\us03\/_0749_ ), .B(\us03\/_0140_ ), .X(\us03\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us03/_0865_ ( .A(\sa03\[0\] ), .B(\sa03\[2\] ), .C(\sa03\[3\] ), .X(\us03\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0866_ ( .A(\us03\/_0043_ ), .B(\us03\/_0045_ ), .X(\us03\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0867_ ( .A(\us03\/_0096_ ), .B(\us03\/_0543_ ), .X(\us03\/_0047_ ) );
sky130_fd_sc_hd__buf_2 \us03/_0868_ ( .A(\us03\/_0047_ ), .X(\us03\/_0048_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0869_ ( .A(\us03\/_0048_ ), .B(\us03\/_0043_ ), .X(\us03\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0870_ ( .A(\us03\/_0730_ ), .X(\us03\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0871_ ( .A(\us03\/_0043_ ), .X(\us03\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_0872_ ( .A1(\us03\/_0118_ ), .A2(\us03\/_0050_ ), .B1(\us03\/_0194_ ), .C1(\us03\/_0051_ ), .Y(\us03\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us03/_0873_ ( .A(\us03\/_0046_ ), .B(\us03\/_0049_ ), .C_N(\us03\/_0052_ ), .Y(\us03\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0874_ ( .A(\us03\/_0026_ ), .B(\us03\/_0140_ ), .X(\us03\/_0054_ ) );
sky130_fd_sc_hd__buf_2 \us03/_0876_ ( .A(\us03\/_0054_ ), .X(\us03\/_0056_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_0877_ ( .A1(\us03\/_0532_ ), .A2(\us03\/_0575_ ), .B1(\us03\/_0056_ ), .Y(\us03\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0878_ ( .A(\us03\/_0412_ ), .B(\us03\/_0325_ ), .X(\us03\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0880_ ( .A(\us03\/_0051_ ), .X(\us03\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_0881_ ( .A1(\us03\/_0732_ ), .A2(\us03\/_0036_ ), .A3(\us03\/_0058_ ), .B1(\us03\/_0060_ ), .Y(\us03\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0882_ ( .A(\us03\/_0260_ ), .B(\sa03\[1\] ), .X(\us03\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0884_ ( .A(\us03\/_0062_ ), .X(\us03\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_0885_ ( .A1(\us03\/_0064_ ), .A2(\us03\/_0748_ ), .A3(\us03\/_0683_ ), .B1(\us03\/_0056_ ), .Y(\us03\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us03/_0886_ ( .A(\us03\/_0053_ ), .B(\us03\/_0057_ ), .C(\us03\/_0061_ ), .D(\us03\/_0065_ ), .X(\us03\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us03/_0887_ ( .A(\us03\/_0629_ ), .B(\us03\/_0745_ ), .C(\us03\/_0042_ ), .D(\us03\/_0066_ ), .X(\us03\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us03/_0889_ ( .A(\sa03\[7\] ), .B_N(\sa03\[6\] ), .Y(\us03\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0890_ ( .A(\us03\/_0069_ ), .B(\us03\/_0151_ ), .X(\us03\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0892_ ( .A(\us03\/_0070_ ), .X(\us03\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_0893_ ( .A1(\us03\/_0129_ ), .A2(\us03\/_0586_ ), .B1(\us03\/_0072_ ), .Y(\us03\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_0894_ ( .A1(\us03\/_0380_ ), .A2(\us03\/_0347_ ), .B1(\us03\/_0194_ ), .B2(\us03\/_0216_ ), .Y(\us03\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us03/_0895_ ( .A(\us03\/_0074_ ), .B_N(\us03\/_0070_ ), .Y(\us03\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us03/_0896_ ( .A(\us03\/_0073_ ), .SLEEP(\us03\/_0075_ ), .X(\us03\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us03/_0897_ ( .A(\us03\/_0467_ ), .B(\us03\/_0069_ ), .X(\us03\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0898_ ( .A(\us03\/_0077_ ), .X(\us03\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0899_ ( .A(\us03\/_0412_ ), .B(\us03\/_0118_ ), .X(\us03\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0901_ ( .A(\us03\/_0078_ ), .B(\us03\/_0079_ ), .X(\us03\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0902_ ( .A(\us03\/_0412_ ), .B(\us03\/_0249_ ), .X(\us03\/_0082_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0905_ ( .A(\us03\/_0280_ ), .B(\us03\/_0078_ ), .X(\us03\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us03/_0906_ ( .A1(\sa03\[0\] ), .A2(\us03\/_0325_ ), .B1(\us03\/_0260_ ), .Y(\us03\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us03/_0907_ ( .A_N(\us03\/_0086_ ), .B(\us03\/_0078_ ), .X(\us03\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us03/_0908_ ( .A(\us03\/_0081_ ), .B(\us03\/_0085_ ), .C(\us03\/_0087_ ), .Y(\us03\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0909_ ( .A(\us03\/_0072_ ), .X(\us03\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_0910_ ( .A1(\us03\/_0733_ ), .A2(\us03\/_0748_ ), .A3(\us03\/_0683_ ), .B1(\us03\/_0089_ ), .Y(\us03\/_0090_ ) );
sky130_fd_sc_hd__buf_2 \us03/_0911_ ( .A(\us03\/_0129_ ), .X(\us03\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0912_ ( .A(\us03\/_0018_ ), .X(\us03\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0913_ ( .A(\us03\/_0022_ ), .X(\us03\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0914_ ( .A(\us03\/_0078_ ), .X(\us03\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_0915_ ( .A1(\us03\/_0091_ ), .A2(\us03\/_0092_ ), .A3(\us03\/_0093_ ), .B1(\us03\/_0094_ ), .Y(\us03\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us03/_0916_ ( .A(\us03\/_0076_ ), .B(\us03\/_0088_ ), .C(\us03\/_0090_ ), .D(\us03\/_0095_ ), .X(\us03\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us03/_0917_ ( .A(\us03\/_0069_ ), .B(\us03\/_0026_ ), .X(\us03\/_0098_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0919_ ( .A(\us03\/_0434_ ), .B(\us03\/_0364_ ), .X(\us03\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0920_ ( .A(\us03\/_0079_ ), .B(\us03\/_0098_ ), .X(\us03\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0921_ ( .A(\us03\/_0325_ ), .X(\us03\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_0922_ ( .A1(\us03\/_0102_ ), .A2(\us03\/_0734_ ), .B1(\us03\/_0038_ ), .C1(\us03\/_0364_ ), .Y(\us03\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us03/_0923_ ( .A(\us03\/_0100_ ), .B(\us03\/_0101_ ), .C_N(\us03\/_0103_ ), .Y(\us03\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_0924_ ( .A1(\us03\/_0554_ ), .A2(\us03\/_0586_ ), .B1(\us03\/_0364_ ), .Y(\us03\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_0925_ ( .A(\us03\/_0129_ ), .B(\us03\/_0364_ ), .Y(\us03\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0926_ ( .A(\us03\/_0105_ ), .B(\us03\/_0106_ ), .X(\us03\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0927_ ( .A(\us03\/_0412_ ), .X(\us03\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us03/_0928_ ( .A(\us03\/_0260_ ), .B(\sa03\[0\] ), .X(\us03\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0929_ ( .A(\us03\/_0069_ ), .B(\us03\/_0749_ ), .X(\us03\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0931_ ( .A(\us03\/_0111_ ), .X(\us03\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0932_ ( .A(\us03\/_0113_ ), .X(\us03\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_0933_ ( .A1(\us03\/_0109_ ), .A2(\us03\/_0110_ ), .B1(\us03\/_0114_ ), .Y(\us03\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us03/_0934_ ( .A(\us03\/_0022_ ), .Y(\us03\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us03/_0935_ ( .A(\us03\/_0554_ ), .Y(\us03\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us03/_0936_ ( .A1(\us03\/_0050_ ), .A2(\us03\/_0118_ ), .B1(\us03\/_0194_ ), .Y(\us03\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us03/_0937_ ( .A(\us03\/_0113_ ), .Y(\us03\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us03/_0938_ ( .A1(\us03\/_0116_ ), .A2(\us03\/_0117_ ), .A3(\us03\/_0119_ ), .B1(\us03\/_0120_ ), .X(\us03\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us03/_0939_ ( .A(\us03\/_0104_ ), .B(\us03\/_0108_ ), .C(\us03\/_0115_ ), .D(\us03\/_0121_ ), .X(\us03\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_0940_ ( .A(\sa03\[7\] ), .B(\sa03\[6\] ), .Y(\us03\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0941_ ( .A(\us03\/_0749_ ), .B(\us03\/_0123_ ), .X(\us03\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0943_ ( .A(\us03\/_0082_ ), .B(\us03\/_0124_ ), .X(\us03\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_0944_ ( .A(\us03\/_0271_ ), .B(\us03\/_0124_ ), .Y(\us03\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0945_ ( .A(\us03\/_0124_ ), .X(\us03\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0946_ ( .A(\us03\/_0260_ ), .B(\us03\/_0325_ ), .X(\us03\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_0948_ ( .A(\us03\/_0128_ ), .B(\us03\/_0130_ ), .Y(\us03\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_0949_ ( .A(\us03\/_0127_ ), .B(\us03\/_0132_ ), .Y(\us03\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us03/_0950_ ( .A(\us03\/_0434_ ), .X(\us03\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_0951_ ( .A(\us03\/_0134_ ), .B(\us03\/_0128_ ), .Y(\us03\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us03/_0952_ ( .A(\us03\/_0126_ ), .B(\us03\/_0133_ ), .C_N(\us03\/_0135_ ), .Y(\us03\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us03/_0953_ ( .A(\us03\/_0026_ ), .B(\us03\/_0123_ ), .X(\us03\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0955_ ( .A(\us03\/_0137_ ), .X(\us03\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_0956_ ( .A1(\us03\/_0110_ ), .A2(\us03\/_0293_ ), .A3(\us03\/_0280_ ), .B1(\us03\/_0139_ ), .Y(\us03\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0957_ ( .A(\us03\/_0096_ ), .B(\us03\/_0730_ ), .X(\us03\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0959_ ( .A(\us03\/_0142_ ), .X(\us03\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_0960_ ( .A1(\us03\/_0020_ ), .A2(\us03\/_0144_ ), .A3(\us03\/_0018_ ), .B1(\us03\/_0139_ ), .Y(\us03\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \us03/_0961_ ( .A(\sa03\[2\] ), .B(\us03\/_0050_ ), .C_N(\sa03\[3\] ), .Y(\us03\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0962_ ( .A(\us03\/_0128_ ), .X(\us03\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_0963_ ( .A1(\us03\/_0146_ ), .A2(\us03\/_0032_ ), .A3(\us03\/_0640_ ), .B1(\us03\/_0147_ ), .Y(\us03\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us03/_0964_ ( .A(\us03\/_0136_ ), .B(\us03\/_0141_ ), .C(\us03\/_0145_ ), .D(\us03\/_0148_ ), .X(\us03\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0965_ ( .A(\us03\/_0123_ ), .B(\us03\/_0151_ ), .X(\us03\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_0967_ ( .A(\us03\/_0150_ ), .X(\us03\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \us03/_0968_ ( .A(\us03\/_0150_ ), .B(\us03\/_0062_ ), .X(\us03\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_0969_ ( .A(\us03\/_0079_ ), .B(\us03\/_0150_ ), .Y(\us03\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us03/_0970_ ( .A(\us03\/_0150_ ), .B(\us03\/_0412_ ), .C(\us03\/_0543_ ), .Y(\us03\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_0971_ ( .A(\us03\/_0155_ ), .B(\us03\/_0156_ ), .Y(\us03\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_0972_ ( .A1(\us03\/_0153_ ), .A2(\us03\/_0134_ ), .B1(\us03\/_0154_ ), .C1(\us03\/_0157_ ), .Y(\us03\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0973_ ( .A(\us03\/_0467_ ), .B(\us03\/_0123_ ), .X(\us03\/_0159_ ) );
sky130_fd_sc_hd__buf_2 \us03/_0975_ ( .A(\us03\/_0159_ ), .X(\us03\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us03/_0976_ ( .A_N(\us03\/_0119_ ), .B(\us03\/_0161_ ), .X(\us03\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us03/_0977_ ( .A(\us03\/_0163_ ), .Y(\us03\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_0978_ ( .A1(\us03\/_0146_ ), .A2(\us03\/_0575_ ), .A3(\us03\/_0608_ ), .B1(\us03\/_0153_ ), .Y(\us03\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_0979_ ( .A1(\us03\/_0062_ ), .A2(\us03\/_0280_ ), .A3(\us03\/_0134_ ), .B1(\us03\/_0161_ ), .Y(\us03\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us03/_0980_ ( .A(\us03\/_0158_ ), .B(\us03\/_0164_ ), .C(\us03\/_0165_ ), .D(\us03\/_0166_ ), .X(\us03\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us03/_0981_ ( .A(\us03\/_0097_ ), .B(\us03\/_0122_ ), .C(\us03\/_0149_ ), .D(\us03\/_0167_ ), .X(\us03\/_0168_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0982_ ( .A(\us03\/_0672_ ), .B(\us03\/_0150_ ), .X(\us03\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_0983_ ( .A(\us03\/_0154_ ), .B(\us03\/_0169_ ), .Y(\us03\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us03/_0984_ ( .A(\us03\/_0123_ ), .B(\us03\/_0151_ ), .C(\us03\/_0038_ ), .X(\us03\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0985_ ( .A(\us03\/_0170_ ), .B(\us03\/_0171_ ), .X(\us03\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \us03/_0986_ ( .A(\us03\/_0172_ ), .Y(\us03\/_0174_ ) );
sky130_fd_sc_hd__nand3_2 \us03/_0987_ ( .A(\us03\/_0067_ ), .B(\us03\/_0168_ ), .C(\us03\/_0174_ ), .Y(\us03\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us03/_0988_ ( .A(\sa03\[1\] ), .B(\sa03\[0\] ), .Y(\us03\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us03/_0989_ ( .A(\us03\/_0175_ ), .B(\us03\/_0358_ ), .X(\us03\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0990_ ( .A(\us03\/_0176_ ), .B(\us03\/_0489_ ), .X(\us03\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_0991_ ( .A(\us03\/_0280_ ), .B(\us03\/_0113_ ), .Y(\us03\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0992_ ( .A(\us03\/_0111_ ), .B(\us03\/_0062_ ), .X(\us03\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0993_ ( .A(\us03\/_0111_ ), .B(\us03\/_0672_ ), .X(\us03\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_0994_ ( .A(\us03\/_0179_ ), .B(\us03\/_0180_ ), .Y(\us03\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0995_ ( .A(\us03\/_0054_ ), .B(\us03\/_0058_ ), .X(\us03\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us03/_0996_ ( .A(\us03\/_0182_ ), .Y(\us03\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us03/_0997_ ( .A_N(\us03\/_0177_ ), .B(\us03\/_0178_ ), .C(\us03\/_0181_ ), .D(\us03\/_0184_ ), .X(\us03\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0998_ ( .A(\us03\/_0098_ ), .B(\us03\/_0741_ ), .X(\us03\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us03/_0999_ ( .A(\us03\/_0047_ ), .B(\us03\/_0098_ ), .X(\us03\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us03/_1000_ ( .A(\us03\/_0186_ ), .B(\us03\/_0187_ ), .X(\us03\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1001_ ( .A(\us03\/_0188_ ), .Y(\us03\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1002_ ( .A(\us03\/_0738_ ), .B(\us03\/_0735_ ), .X(\us03\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1003_ ( .A(\us03\/_0271_ ), .B(\us03\/_0736_ ), .X(\us03\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_1004_ ( .A(\us03\/_0190_ ), .B(\us03\/_0191_ ), .Y(\us03\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us03/_1005_ ( .A(\us03\/_0096_ ), .B(\us03\/_0325_ ), .X(\us03\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1006_ ( .A1(\us03\/_0193_ ), .A2(\us03\/_0176_ ), .B1(\us03\/_0043_ ), .Y(\us03\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1007_ ( .A(\us03\/_0185_ ), .B(\us03\/_0189_ ), .C(\us03\/_0192_ ), .D(\us03\/_0195_ ), .X(\us03\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us03/_1008_ ( .A_N(\sa03\[3\] ), .B(\us03\/_0734_ ), .C(\sa03\[2\] ), .X(\us03\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1009_ ( .A(\us03\/_0137_ ), .B(\us03\/_0197_ ), .X(\us03\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_1010_ ( .A(\us03\/_0198_ ), .B(\us03\/_0040_ ), .Y(\us03\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1011_ ( .A(\us03\/_0293_ ), .B(\us03\/_0137_ ), .X(\us03\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1012_ ( .A(\us03\/_0200_ ), .Y(\us03\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1013_ ( .A(\us03\/_0137_ ), .B(\us03\/_0110_ ), .Y(\us03\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1014_ ( .A(\us03\/_0139_ ), .B(\us03\/_0020_ ), .Y(\us03\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1015_ ( .A(\us03\/_0199_ ), .B(\us03\/_0201_ ), .C(\us03\/_0202_ ), .D(\us03\/_0203_ ), .X(\us03\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us03/_1016_ ( .A1(\us03\/_0532_ ), .A2(\us03\/_0109_ ), .B1(\us03\/_0102_ ), .C1(\us03\/_0727_ ), .X(\us03\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1017_ ( .A(\us03\/_0022_ ), .B(\us03\/_0078_ ), .Y(\us03\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1018_ ( .A(\us03\/_0078_ ), .B(\us03\/_0142_ ), .Y(\us03\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1019_ ( .A(\us03\/_0207_ ), .B(\us03\/_0208_ ), .Y(\us03\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1020_ ( .A1(\us03\/_0094_ ), .A2(\us03\/_0176_ ), .B1(\us03\/_0206_ ), .C1(\us03\/_0209_ ), .Y(\us03\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1021_ ( .A(\us03\/_0662_ ), .B(\us03\/_0070_ ), .X(\us03\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us03/_1022_ ( .A(\us03\/_0732_ ), .B(\us03\/_0123_ ), .C(\us03\/_0749_ ), .Y(\us03\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us03/_1023_ ( .A(\us03\/_0732_ ), .B(\us03\/_0467_ ), .C(\us03\/_0069_ ), .Y(\us03\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us03/_1024_ ( .A_N(\us03\/_0211_ ), .B(\us03\/_0127_ ), .C(\us03\/_0212_ ), .D(\us03\/_0213_ ), .X(\us03\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1025_ ( .A(\us03\/_0137_ ), .Y(\us03\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1026_ ( .A(\us03\/_0128_ ), .B(\us03\/_0036_ ), .Y(\us03\/_0217_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1028_ ( .A1(\us03\/_0159_ ), .A2(\us03\/_0747_ ), .B1(\us03\/_0434_ ), .B2(\us03\/_0499_ ), .Y(\us03\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us03/_1029_ ( .A1(\us03\/_0116_ ), .A2(\us03\/_0215_ ), .B1(\us03\/_0217_ ), .C1(\us03\/_0219_ ), .X(\us03\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1030_ ( .A(\us03\/_0113_ ), .B(\us03\/_0746_ ), .X(\us03\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us03/_1031_ ( .A1(\us03\/_0098_ ), .A2(\us03\/_0746_ ), .B1(\us03\/_0434_ ), .B2(\us03\/_0750_ ), .X(\us03\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1032_ ( .A1(\us03\/_0048_ ), .A2(\us03\/_0113_ ), .B1(\us03\/_0221_ ), .C1(\us03\/_0222_ ), .Y(\us03\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us03/_1033_ ( .A1(\us03\/_0129_ ), .A2(\us03\/_0162_ ), .B1(\us03\/_0271_ ), .B2(\us03\/_0705_ ), .X(\us03\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1034_ ( .A1(\us03\/_0093_ ), .A2(\us03\/_0738_ ), .B1(\us03\/_0081_ ), .C1(\us03\/_0224_ ), .Y(\us03\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1035_ ( .A(\us03\/_0214_ ), .B(\us03\/_0220_ ), .C(\us03\/_0223_ ), .D(\us03\/_0225_ ), .X(\us03\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1036_ ( .A(\us03\/_0196_ ), .B(\us03\/_0204_ ), .C(\us03\/_0210_ ), .D(\us03\/_0226_ ), .X(\us03\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1037_ ( .A(\us03\/_0111_ ), .B(\us03\/_0554_ ), .X(\us03\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1038_ ( .A(\us03\/_0229_ ), .Y(\us03\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1039_ ( .A(\us03\/_0111_ ), .B(\us03\/_0129_ ), .Y(\us03\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1040_ ( .A(\us03\/_0018_ ), .B(\us03\/_0738_ ), .Y(\us03\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1041_ ( .A(\us03\/_0030_ ), .B(\us03\/_0304_ ), .Y(\us03\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1042_ ( .A(\us03\/_0230_ ), .B(\us03\/_0231_ ), .C(\us03\/_0232_ ), .D(\us03\/_0233_ ), .X(\us03\/_0234_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1043_ ( .A(\us03\/_0048_ ), .B(\us03\/_0489_ ), .X(\us03\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1044_ ( .A1(\us03\/_0129_ ), .A2(\us03\/_0554_ ), .B1(\us03\/_0137_ ), .Y(\us03\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us03/_1045_ ( .A(\us03\/_0235_ ), .B(\us03\/_0049_ ), .C_N(\us03\/_0236_ ), .Y(\us03\/_0237_ ) );
sky130_fd_sc_hd__and2_1 \us03/_1046_ ( .A(\us03\/_0047_ ), .B(\us03\/_0077_ ), .X(\us03\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1047_ ( .A(\us03\/_0070_ ), .B(\us03\/_0036_ ), .X(\us03\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us03/_1048_ ( .A1(\us03\/_0048_ ), .A2(\us03\/_0736_ ), .B1(\us03\/_0022_ ), .B2(\us03\/_0364_ ), .X(\us03\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us03/_1049_ ( .A(\us03\/_0239_ ), .B(\us03\/_0240_ ), .C(\us03\/_0241_ ), .Y(\us03\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1050_ ( .A(\us03\/_0554_ ), .B(\us03\/_0072_ ), .X(\us03\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us03/_1051_ ( .A1(\us03\/_0142_ ), .A2(\us03\/_0137_ ), .B1(\us03\/_0159_ ), .B2(\us03\/_0082_ ), .X(\us03\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1052_ ( .A1(\us03\/_0608_ ), .A2(\us03\/_0072_ ), .B1(\us03\/_0243_ ), .C1(\us03\/_0244_ ), .Y(\us03\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1053_ ( .A(\us03\/_0234_ ), .B(\us03\/_0237_ ), .C(\us03\/_0242_ ), .D(\us03\/_0245_ ), .X(\us03\/_0246_ ) );
sky130_fd_sc_hd__buf_2 \us03/_1054_ ( .A(\us03\/_0028_ ), .X(\us03\/_0247_ ) );
sky130_fd_sc_hd__o21a_1 \us03/_1055_ ( .A1(\us03\/_0554_ ), .A2(\us03\/_0586_ ), .B1(\us03\/_0247_ ), .X(\us03\/_0248_ ) );
sky130_fd_sc_hd__and2_1 \us03/_1056_ ( .A(\us03\/_0082_ ), .B(\us03\/_0489_ ), .X(\us03\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_1057_ ( .A(\us03\/_0079_ ), .X(\us03\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1058_ ( .A(\us03\/_0251_ ), .B(\us03\/_0489_ ), .X(\us03\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_1059_ ( .A(\us03\/_0250_ ), .B(\us03\/_0252_ ), .Y(\us03\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1060_ ( .A(\us03\/_0016_ ), .B(\us03\/_0064_ ), .Y(\us03\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_1061_ ( .A(\us03\/_0304_ ), .X(\us03\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1062_ ( .A(\us03\/_0255_ ), .B(\us03\/_0640_ ), .Y(\us03\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us03/_1063_ ( .A_N(\us03\/_0248_ ), .B(\us03\/_0253_ ), .C(\us03\/_0254_ ), .D(\us03\/_0256_ ), .X(\us03\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1064_ ( .A(\us03\/_0364_ ), .B(\us03\/_0110_ ), .X(\us03\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us03/_1065_ ( .A1(\us03\/_0161_ ), .A2(\us03\/_0130_ ), .B1(\us03\/_0258_ ), .Y(\us03\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1066_ ( .A(\us03\/_0194_ ), .B(\sa03\[1\] ), .X(\us03\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1068_ ( .A(\us03\/_0261_ ), .B(\us03\/_0153_ ), .Y(\us03\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us03/_1069_ ( .A_N(\us03\/_0154_ ), .B(\us03\/_0259_ ), .C(\us03\/_0263_ ), .X(\us03\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1070_ ( .A(\us03\/_0246_ ), .B(\us03\/_0174_ ), .C(\us03\/_0257_ ), .D(\us03\/_0264_ ), .X(\us03\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us03/_1071_ ( .A1(\us03\/_0261_ ), .A2(\us03\/_0554_ ), .B1(\us03\/_0159_ ), .X(\us03\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1072_ ( .A(\us03\/_0747_ ), .B(\us03\/_0150_ ), .Y(\us03\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1073_ ( .A(\us03\/_0175_ ), .Y(\us03\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us03/_1074_ ( .A(\us03\/_0412_ ), .B(\us03\/_0123_ ), .C(\us03\/_0151_ ), .X(\us03\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1075_ ( .A(\us03\/_0268_ ), .B(\us03\/_0269_ ), .Y(\us03\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us03/_1076_ ( .A_N(\us03\/_0266_ ), .B(\us03\/_0267_ ), .C(\us03\/_0270_ ), .X(\us03\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1077_ ( .A(\us03\/_0554_ ), .B(\us03\/_0150_ ), .X(\us03\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1078_ ( .A(\us03\/_0273_ ), .Y(\us03\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1079_ ( .A1(\us03\/_0734_ ), .A2(\us03\/_0325_ ), .B1(\us03\/_0380_ ), .Y(\us03\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1080_ ( .A(\us03\/_0275_ ), .Y(\us03\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1081_ ( .A(\us03\/_0276_ ), .B(\us03\/_0153_ ), .Y(\us03\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us03/_1082_ ( .A(\us03\/_0272_ ), .B(\us03\/_0274_ ), .C(\us03\/_0277_ ), .X(\us03\/_0278_ ) );
sky130_fd_sc_hd__buf_2 \us03/_1083_ ( .A(\us03\/_0036_ ), .X(\us03\/_0279_ ) );
sky130_fd_sc_hd__buf_2 \us03/_1084_ ( .A(\us03\/_0082_ ), .X(\us03\/_0280_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1085_ ( .A1(\us03\/_0499_ ), .A2(\us03\/_0279_ ), .B1(\us03\/_0280_ ), .B2(\us03\/_0060_ ), .Y(\us03\/_0281_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1086_ ( .A1(\us03\/_0251_ ), .A2(\us03\/_0434_ ), .B1(\us03\/_0304_ ), .Y(\us03\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1087_ ( .A(\us03\/_0091_ ), .B(\us03\/_0056_ ), .Y(\us03\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1088_ ( .A1(\us03\/_0118_ ), .A2(\us03\/_0050_ ), .B1(\us03\/_0038_ ), .C1(\us03\/_0255_ ), .Y(\us03\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1089_ ( .A(\us03\/_0281_ ), .B(\us03\/_0283_ ), .C(\us03\/_0284_ ), .D(\us03\/_0285_ ), .X(\us03\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1090_ ( .A(\us03\/_0082_ ), .B(\us03\/_0028_ ), .X(\us03\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1091_ ( .A(\us03\/_0129_ ), .B(\us03\/_0028_ ), .X(\us03\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_1092_ ( .A(\us03\/_0287_ ), .B(\us03\/_0288_ ), .Y(\us03\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1093_ ( .A1(\us03\/_0752_ ), .A2(\us03\/_0683_ ), .B1(\us03\/_0093_ ), .B2(\us03\/_0247_ ), .Y(\us03\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1094_ ( .A1(\us03\/_0092_ ), .A2(\us03\/_0575_ ), .B1(\us03\/_0056_ ), .Y(\us03\/_0291_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1096_ ( .A1(\us03\/_0499_ ), .A2(\us03\/_0672_ ), .B1(\us03\/_0280_ ), .B2(\us03\/_0056_ ), .Y(\us03\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1097_ ( .A(\us03\/_0289_ ), .B(\us03\/_0290_ ), .C(\us03\/_0291_ ), .D(\us03\/_0294_ ), .X(\us03\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1098_ ( .A(\us03\/_0750_ ), .B(\us03\/_0193_ ), .X(\us03\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1099_ ( .A(\us03\/_0705_ ), .B(\us03\/_0380_ ), .X(\us03\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1100_ ( .A(\us03\/_0752_ ), .B(\us03\/_0129_ ), .Y(\us03\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us03/_1101_ ( .A(\us03\/_0296_ ), .B(\us03\/_0297_ ), .C_N(\us03\/_0298_ ), .Y(\us03\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1102_ ( .A(\us03\/_0089_ ), .B(\us03\/_0532_ ), .Y(\us03\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1103_ ( .A(\sa03\[2\] ), .Y(\us03\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \us03/_1104_ ( .A(\us03\/_0301_ ), .B(\sa03\[3\] ), .C(\us03\/_0118_ ), .Y(\us03\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1105_ ( .A(\us03\/_0072_ ), .B(\us03\/_0302_ ), .X(\us03\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1106_ ( .A(\us03\/_0303_ ), .Y(\us03\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1107_ ( .A(\us03\/_0147_ ), .B(\us03\/_0302_ ), .Y(\us03\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1108_ ( .A(\us03\/_0299_ ), .B(\us03\/_0300_ ), .C(\us03\/_0305_ ), .D(\us03\/_0306_ ), .X(\us03\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1109_ ( .A(\us03\/_0278_ ), .B(\us03\/_0286_ ), .C(\us03\/_0295_ ), .D(\us03\/_0307_ ), .X(\us03\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us03/_1110_ ( .A(\us03\/_0228_ ), .B(\us03\/_0265_ ), .C(\us03\/_0308_ ), .Y(\us03\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1111_ ( .A(\us03\/_0235_ ), .Y(\us03\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1112_ ( .A(\us03\/_0489_ ), .B(\us03\/_0640_ ), .X(\us03\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1113_ ( .A(\us03\/_0310_ ), .Y(\us03\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1114_ ( .A(\us03\/_0022_ ), .B(\us03\/_0499_ ), .Y(\us03\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1115_ ( .A(\us03\/_0499_ ), .B(\us03\/_0032_ ), .Y(\us03\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1116_ ( .A(\us03\/_0309_ ), .B(\us03\/_0311_ ), .C(\us03\/_0312_ ), .D(\us03\/_0313_ ), .X(\us03\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1117_ ( .A(\us03\/_0499_ ), .B(\us03\/_0064_ ), .Y(\us03\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1118_ ( .A(\us03\/_0499_ ), .B(\us03\/_0683_ ), .Y(\us03\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1119_ ( .A(\us03\/_0315_ ), .B(\us03\/_0316_ ), .C(\us03\/_0317_ ), .D(\us03\/_0253_ ), .X(\us03\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1120_ ( .A(\us03\/_0048_ ), .B(\us03\/_0304_ ), .Y(\us03\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1121_ ( .A(\us03\/_0586_ ), .B(\us03\/_0162_ ), .Y(\us03\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1122_ ( .A(\us03\/_0319_ ), .B(\us03\/_0320_ ), .Y(\us03\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_1123_ ( .A(\us03\/_0321_ ), .B(\us03\/_0238_ ), .Y(\us03\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1124_ ( .A(\us03\/_0304_ ), .B(\us03\/_0062_ ), .Y(\us03\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_1125_ ( .A(\us03\/_0251_ ), .X(\us03\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1126_ ( .A1(\us03\/_0324_ ), .A2(\us03\/_0280_ ), .B1(\us03\/_0255_ ), .Y(\us03\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1127_ ( .A1(\us03\/_0050_ ), .A2(\us03\/_0216_ ), .B1(\us03\/_0109_ ), .C1(\us03\/_0255_ ), .Y(\us03\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1128_ ( .A(\us03\/_0322_ ), .B(\us03\/_0323_ ), .C(\us03\/_0326_ ), .D(\us03\/_0327_ ), .X(\us03\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1129_ ( .A1(\us03\/_0733_ ), .A2(\us03\/_0279_ ), .A3(\us03\/_0058_ ), .B1(\us03\/_0056_ ), .Y(\us03\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_1130_ ( .A(\us03\/_0048_ ), .X(\us03\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1131_ ( .A(\us03\/_0330_ ), .B(\us03\/_0056_ ), .Y(\us03\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1132_ ( .A(\us03\/_0054_ ), .B(\us03\/_0045_ ), .Y(\us03\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1133_ ( .A(\us03\/_0329_ ), .B(\us03\/_0331_ ), .C(\us03\/_0284_ ), .D(\us03\/_0332_ ), .X(\us03\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us03/_1134_ ( .A1(\us03\/_0543_ ), .A2(\us03\/_0216_ ), .B1(\us03\/_0532_ ), .C1(\us03\/_0060_ ), .X(\us03\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1135_ ( .A(\us03\/_0280_ ), .B(\us03\/_0060_ ), .Y(\us03\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1136_ ( .A(\us03\/_0324_ ), .B(\us03\/_0060_ ), .Y(\us03\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1137_ ( .A(\us03\/_0335_ ), .B(\us03\/_0337_ ), .Y(\us03\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1138_ ( .A1(\us03\/_0276_ ), .A2(\us03\/_0060_ ), .B1(\us03\/_0334_ ), .C1(\us03\/_0338_ ), .Y(\us03\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1139_ ( .A(\us03\/_0318_ ), .B(\us03\/_0328_ ), .C(\us03\/_0333_ ), .D(\us03\/_0339_ ), .X(\us03\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us03/_1140_ ( .A1(\us03\/_0747_ ), .A2(\us03\/_0134_ ), .B1(\us03\/_0128_ ), .X(\us03\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us03/_1141_ ( .A_N(\us03\/_0086_ ), .B(\us03\/_0128_ ), .X(\us03\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1142_ ( .A(\us03\/_0079_ ), .B(\us03\/_0124_ ), .X(\us03\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_1143_ ( .A(\us03\/_0126_ ), .B(\us03\/_0343_ ), .Y(\us03\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us03/_1144_ ( .A(\us03\/_0341_ ), .B(\us03\/_0342_ ), .C_N(\us03\/_0344_ ), .Y(\us03\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1146_ ( .A1(\us03\/_0193_ ), .A2(\us03\/_0092_ ), .A3(\us03\/_0330_ ), .B1(\us03\/_0147_ ), .Y(\us03\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1147_ ( .A1(\us03\/_0130_ ), .A2(\us03\/_0280_ ), .A3(\us03\/_0134_ ), .B1(\us03\/_0139_ ), .Y(\us03\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1148_ ( .A1(\us03\/_0144_ ), .A2(\us03\/_0608_ ), .A3(\us03\/_0092_ ), .B1(\us03\/_0139_ ), .Y(\us03\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1149_ ( .A(\us03\/_0345_ ), .B(\us03\/_0348_ ), .C(\us03\/_0349_ ), .D(\us03\/_0350_ ), .X(\us03\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us03/_1150_ ( .A(\us03\/_0150_ ), .B(\us03\/_0194_ ), .C(\us03\/_0543_ ), .X(\us03\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us03/_1151_ ( .A(\us03\/_0277_ ), .SLEEP(\us03\/_0352_ ), .X(\us03\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us03/_1152_ ( .A1(\us03\/_0268_ ), .A2(\us03\/_0171_ ), .B1(\us03\/_0157_ ), .Y(\us03\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us03/_1153_ ( .A(\us03\/_0161_ ), .X(\us03\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1154_ ( .A1(\us03\/_0279_ ), .A2(\us03\/_0280_ ), .B1(\us03\/_0355_ ), .Y(\us03\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1155_ ( .A1(\us03\/_0020_ ), .A2(\us03\/_0193_ ), .A3(\us03\/_0091_ ), .B1(\us03\/_0355_ ), .Y(\us03\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1156_ ( .A(\us03\/_0353_ ), .B(\us03\/_0354_ ), .C(\us03\/_0356_ ), .D(\us03\/_0357_ ), .X(\us03\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1157_ ( .A(\us03\/_0111_ ), .B(\us03\/_0586_ ), .X(\us03\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1158_ ( .A(\us03\/_0360_ ), .Y(\us03\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us03/_1159_ ( .A1(\us03\/_0119_ ), .A2(\us03\/_0120_ ), .B1(\us03\/_0230_ ), .C1(\us03\/_0361_ ), .X(\us03\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1160_ ( .A1(\us03\/_0672_ ), .A2(\us03\/_0251_ ), .A3(\us03\/_0134_ ), .B1(\us03\/_0114_ ), .Y(\us03\/_0363_ ) );
sky130_fd_sc_hd__buf_2 \us03/_1161_ ( .A(\us03\/_0098_ ), .X(\us03\/_0364_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1162_ ( .A1(\us03\/_0036_ ), .A2(\us03\/_0251_ ), .A3(\us03\/_0134_ ), .B1(\us03\/_0364_ ), .Y(\us03\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1163_ ( .A1(\us03\/_0193_ ), .A2(\us03\/_0608_ ), .B1(\us03\/_0364_ ), .Y(\us03\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1164_ ( .A(\us03\/_0362_ ), .B(\us03\/_0363_ ), .C(\us03\/_0365_ ), .D(\us03\/_0366_ ), .X(\us03\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1165_ ( .A1(\us03\/_0575_ ), .A2(\us03\/_0092_ ), .A3(\us03\/_0330_ ), .B1(\us03\/_0089_ ), .Y(\us03\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1166_ ( .A1(\us03\/_0586_ ), .A2(\us03\/_0018_ ), .A3(\us03\/_0330_ ), .B1(\us03\/_0094_ ), .Y(\us03\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \us03/_1167_ ( .A1(\us03\/_0293_ ), .A2(\us03\/_0134_ ), .B1(\us03\/_0089_ ), .Y(\us03\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1168_ ( .A1(\us03\/_0279_ ), .A2(\us03\/_0134_ ), .B1(\us03\/_0094_ ), .Y(\us03\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1169_ ( .A(\us03\/_0368_ ), .B(\us03\/_0370_ ), .C(\us03\/_0371_ ), .D(\us03\/_0372_ ), .X(\us03\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1170_ ( .A(\us03\/_0351_ ), .B(\us03\/_0359_ ), .C(\us03\/_0367_ ), .D(\us03\/_0373_ ), .X(\us03\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1171_ ( .A1(\us03\/_0102_ ), .A2(\us03\/_0347_ ), .B1(\us03\/_0109_ ), .C1(\us03\/_0247_ ), .Y(\us03\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1172_ ( .A1(\us03\/_0102_ ), .A2(\us03\/_0347_ ), .B1(\us03\/_0532_ ), .C1(\us03\/_0247_ ), .Y(\us03\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1173_ ( .A1(\us03\/_0050_ ), .A2(\us03\/_0543_ ), .B1(\us03\/_0380_ ), .C1(\us03\/_0247_ ), .Y(\us03\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1174_ ( .A(\us03\/_0041_ ), .B(\us03\/_0375_ ), .C(\us03\/_0376_ ), .D(\us03\/_0377_ ), .X(\us03\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1175_ ( .A(\us03\/_0048_ ), .B(\us03\/_0750_ ), .X(\us03\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1176_ ( .A(\us03\/_0379_ ), .Y(\us03\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1177_ ( .A(\us03\/_0016_ ), .B(\us03\/_0608_ ), .Y(\us03\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1178_ ( .A(\us03\/_0752_ ), .B(\us03\/_0554_ ), .Y(\us03\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1179_ ( .A1(\sa03\[1\] ), .A2(\us03\/_0734_ ), .B1(\us03\/_0109_ ), .C1(\us03\/_0016_ ), .Y(\us03\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1180_ ( .A(\us03\/_0381_ ), .B(\us03\/_0382_ ), .C(\us03\/_0383_ ), .D(\us03\/_0384_ ), .X(\us03\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us03/_1181_ ( .A(\us03\/_0086_ ), .B_N(\us03\/_0736_ ), .X(\us03\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1182_ ( .A1(\us03\/_0748_ ), .A2(\us03\/_0134_ ), .B1(\us03\/_0739_ ), .Y(\us03\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1183_ ( .A1(\us03\/_0118_ ), .A2(\us03\/_0543_ ), .B1(\us03\/_0109_ ), .C1(\us03\/_0739_ ), .Y(\us03\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1184_ ( .A1(\us03\/_0102_ ), .A2(\us03\/_0301_ ), .B1(\sa03\[3\] ), .C1(\us03\/_0739_ ), .Y(\us03\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1185_ ( .A(\us03\/_0386_ ), .B(\us03\/_0387_ ), .C(\us03\/_0388_ ), .D(\us03\/_0389_ ), .X(\us03\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1186_ ( .A(\us03\/_0020_ ), .Y(\us03\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1187_ ( .A(\us03\/_0727_ ), .Y(\us03\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1188_ ( .A(\us03\/_0727_ ), .B(\us03\/_0064_ ), .Y(\us03\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1189_ ( .A1(\us03\/_0102_ ), .A2(\us03\/_0734_ ), .B1(\us03\/_0532_ ), .C1(\us03\/_0727_ ), .Y(\us03\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us03/_1190_ ( .A1(\us03\/_0392_ ), .A2(\us03\/_0393_ ), .B1(\us03\/_0394_ ), .C1(\us03\/_0395_ ), .X(\us03\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1191_ ( .A(\us03\/_0378_ ), .B(\us03\/_0385_ ), .C(\us03\/_0390_ ), .D(\us03\/_0396_ ), .X(\us03\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us03/_1192_ ( .A(\us03\/_0340_ ), .B(\us03\/_0374_ ), .C(\us03\/_0397_ ), .Y(\us03\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1193_ ( .A(\us03\/_0077_ ), .B(\us03\/_0129_ ), .X(\us03\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_1194_ ( .A(\us03\/_0398_ ), .B(\us03\/_0239_ ), .Y(\us03\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1195_ ( .A(\us03\/_0022_ ), .B(\us03\/_0111_ ), .X(\us03\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us03/_1196_ ( .A_N(\us03\/_0400_ ), .B(\us03\/_0231_ ), .Y(\us03\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us03/_1197_ ( .A(\us03\/_0399_ ), .SLEEP(\us03\/_0402_ ), .X(\us03\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_1198_ ( .A(\us03\/_0747_ ), .B(\us03\/_0251_ ), .Y(\us03\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us03/_1199_ ( .A_N(\us03\/_0404_ ), .B(\us03\/_0752_ ), .Y(\us03\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us03/_1200_ ( .A(\us03\/_0467_ ), .B(\us03\/_0194_ ), .C(\us03\/_0694_ ), .X(\us03\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us03/_1201_ ( .A_N(\us03\/_0175_ ), .B(\us03\/_0406_ ), .X(\us03\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1202_ ( .A(\us03\/_0407_ ), .Y(\us03\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1203_ ( .A1(\us03\/_0094_ ), .A2(\us03\/_0197_ ), .B1(\us03\/_0114_ ), .B2(\us03\/_0640_ ), .Y(\us03\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1204_ ( .A(\us03\/_0403_ ), .B(\us03\/_0405_ ), .C(\us03\/_0408_ ), .D(\us03\/_0409_ ), .X(\us03\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1205_ ( .A(\us03\/_0030_ ), .B(\us03\/_0150_ ), .Y(\us03\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us03/_1206_ ( .A_N(\us03\/_0169_ ), .B(\us03\/_0289_ ), .C(\us03\/_0411_ ), .X(\us03\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us03/_1207_ ( .A1(\us03\/_0467_ ), .A2(\us03\/_0151_ ), .B1(\us03\/_0140_ ), .C1(\us03\/_0129_ ), .X(\us03\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1208_ ( .A1(\us03\/_0608_ ), .A2(\us03\/_0364_ ), .B1(\us03\/_0037_ ), .C1(\us03\/_0414_ ), .Y(\us03\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1209_ ( .A(\us03\/_0738_ ), .Y(\us03\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1210_ ( .A(\us03\/_0586_ ), .B(\us03\/_0736_ ), .Y(\us03\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1211_ ( .A1(\us03\/_0194_ ), .A2(\us03\/_0038_ ), .B1(\us03\/_0118_ ), .C1(\us03\/_0153_ ), .Y(\us03\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us03/_1212_ ( .A1(\us03\/_0416_ ), .A2(\us03\/_0117_ ), .B1(\us03\/_0417_ ), .C1(\us03\/_0418_ ), .X(\us03\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1213_ ( .A(\us03\/_0077_ ), .B(\us03\/_0035_ ), .X(\us03\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1214_ ( .A(\us03\/_0672_ ), .B(\us03\/_0124_ ), .Y(\us03\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1215_ ( .A(\us03\/_0030_ ), .B(\us03\/_0137_ ), .Y(\us03\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1216_ ( .A(\us03\/_0072_ ), .B(\us03\/_0732_ ), .Y(\us03\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us03/_1217_ ( .A_N(\us03\/_0420_ ), .B(\us03\/_0421_ ), .C(\us03\/_0422_ ), .D(\us03\/_0424_ ), .X(\us03\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1218_ ( .A(\us03\/_0413_ ), .B(\us03\/_0415_ ), .C(\us03\/_0419_ ), .D(\us03\/_0425_ ), .X(\us03\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us03/_1219_ ( .A(\us03\/_0355_ ), .B(\us03\/_0102_ ), .C(\us03\/_0109_ ), .Y(\us03\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1220_ ( .A(\us03\/_0077_ ), .B(\us03\/_0018_ ), .X(\us03\/_0428_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1221_ ( .A(\us03\/_0077_ ), .B(\us03\/_0554_ ), .X(\us03\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us03/_1222_ ( .A1(\us03\/_0050_ ), .A2(\us03\/_0216_ ), .B1(\us03\/_0380_ ), .C1(\us03\/_0078_ ), .X(\us03\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us03/_1223_ ( .A(\us03\/_0428_ ), .B(\us03\/_0429_ ), .C(\us03\/_0430_ ), .Y(\us03\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us03/_1224_ ( .A_N(\us03\/_0209_ ), .B(\us03\/_0431_ ), .X(\us03\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us03/_1225_ ( .A1(\us03\/_0215_ ), .A2(\us03\/_0404_ ), .B1(\us03\/_0427_ ), .C1(\us03\/_0432_ ), .X(\us03\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1226_ ( .A(\us03\/_0043_ ), .B(\us03\/_0058_ ), .Y(\us03\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1227_ ( .A(\us03\/_0195_ ), .B(\us03\/_0233_ ), .C(\us03\/_0320_ ), .D(\us03\/_0435_ ), .X(\us03\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1228_ ( .A(\us03\/_0261_ ), .B(\us03\/_0738_ ), .Y(\us03\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1229_ ( .A1(\us03\/_0499_ ), .A2(\us03\/_0640_ ), .B1(\us03\/_0261_ ), .B2(\us03\/_0056_ ), .Y(\us03\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1230_ ( .A(\us03\/_0436_ ), .B(\us03\/_0394_ ), .C(\us03\/_0437_ ), .D(\us03\/_0438_ ), .X(\us03\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1231_ ( .A(\us03\/_0410_ ), .B(\us03\/_0426_ ), .C(\us03\/_0433_ ), .D(\us03\/_0439_ ), .X(\us03\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us03/_1232_ ( .A(\us03\/_0135_ ), .SLEEP(\us03\/_0273_ ), .X(\us03\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1233_ ( .A1(\us03\/_0279_ ), .A2(\us03\/_0134_ ), .B1(\us03\/_0364_ ), .Y(\us03\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1234_ ( .A(\us03\/_0441_ ), .B(\us03\/_0164_ ), .C(\us03\/_0270_ ), .D(\us03\/_0442_ ), .X(\us03\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1235_ ( .A(\us03\/_0051_ ), .B(\us03\/_0672_ ), .Y(\us03\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1236_ ( .A(\us03\/_0051_ ), .B(\us03\/_0271_ ), .Y(\us03\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1237_ ( .A(\us03\/_0444_ ), .B(\us03\/_0446_ ), .X(\us03\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1238_ ( .A(\us03\/_0193_ ), .B(\us03\/_0304_ ), .X(\us03\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1239_ ( .A(\us03\/_0448_ ), .Y(\us03\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1240_ ( .A(\us03\/_0162_ ), .B(\us03\/_0130_ ), .X(\us03\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1241_ ( .A(\us03\/_0450_ ), .Y(\us03\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1242_ ( .A1(\us03\/_0129_ ), .A2(\us03\/_0554_ ), .B1(\us03\/_0043_ ), .Y(\us03\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1243_ ( .A(\us03\/_0447_ ), .B(\us03\/_0449_ ), .C(\us03\/_0451_ ), .D(\us03\/_0452_ ), .X(\us03\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1244_ ( .A(\us03\/_0056_ ), .B(\us03\/_0064_ ), .Y(\us03\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us03/_1245_ ( .A_N(\us03\/_0248_ ), .B(\us03\/_0454_ ), .C(\us03\/_0254_ ), .D(\us03\/_0256_ ), .X(\us03\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1246_ ( .A1(\us03\/_0330_ ), .A2(\us03\/_0364_ ), .B1(\us03\/_0134_ ), .B2(\us03\/_0705_ ), .Y(\us03\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1247_ ( .A1(\us03\/_0748_ ), .A2(\us03\/_0738_ ), .B1(\us03\/_0092_ ), .B2(\us03\/_0752_ ), .Y(\us03\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1248_ ( .A1(\us03\/_0072_ ), .A2(\us03\/_0036_ ), .B1(\us03\/_0748_ ), .B2(\us03\/_0056_ ), .Y(\us03\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1249_ ( .A1(\us03\/_0748_ ), .A2(\us03\/_0251_ ), .B1(\us03\/_0247_ ), .Y(\us03\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1250_ ( .A(\us03\/_0457_ ), .B(\us03\/_0458_ ), .C(\us03\/_0459_ ), .D(\us03\/_0460_ ), .X(\us03\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1251_ ( .A(\us03\/_0443_ ), .B(\us03\/_0453_ ), .C(\us03\/_0455_ ), .D(\us03\/_0461_ ), .X(\us03\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1252_ ( .A(\us03\/_0705_ ), .B(\us03\/_0079_ ), .X(\us03\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1253_ ( .A(\us03\/_0586_ ), .B(\us03\/_0124_ ), .Y(\us03\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1254_ ( .A(\us03\/_0499_ ), .B(\us03\/_0747_ ), .Y(\us03\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us03/_1255_ ( .A_N(\us03\/_0463_ ), .B(\us03\/_0464_ ), .C(\us03\/_0465_ ), .X(\us03\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us03/_1256_ ( .A1(\us03\/_0271_ ), .A2(\us03\/_0072_ ), .B1(\us03\/_0142_ ), .B2(\us03\/_0028_ ), .X(\us03\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1257_ ( .A1(\us03\/_0144_ ), .A2(\us03\/_0364_ ), .B1(\us03\/_0360_ ), .C1(\us03\/_0468_ ), .Y(\us03\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us03/_1258_ ( .A1(\us03\/_0672_ ), .A2(\us03\/_0251_ ), .B1(\us03\/_0499_ ), .X(\us03\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1259_ ( .A1(\us03\/_0575_ ), .A2(\us03\/_0056_ ), .B1(\us03\/_0379_ ), .C1(\us03\/_0470_ ), .Y(\us03\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1260_ ( .A(\us03\/_0466_ ), .B(\us03\/_0469_ ), .C(\us03\/_0471_ ), .D(\us03\/_0305_ ), .X(\us03\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us03/_1261_ ( .A1(\us03\/_0247_ ), .A2(\us03\/_0683_ ), .B1(\us03\/_0324_ ), .B2(\us03\/_0056_ ), .X(\us03\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1262_ ( .A(\us03\/_0280_ ), .B(\us03\/_0364_ ), .X(\us03\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us03/_1263_ ( .A1(\us03\/_0092_ ), .A2(\us03\/_0247_ ), .B1(\us03\/_0474_ ), .X(\us03\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us03/_1264_ ( .A(\us03\/_0075_ ), .B(\us03\/_0473_ ), .C(\us03\/_0475_ ), .Y(\us03\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1265_ ( .A1(\us03\/_0279_ ), .A2(\us03\/_0255_ ), .B1(\us03\/_0280_ ), .B2(\us03\/_0060_ ), .Y(\us03\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1266_ ( .A1(\us03\/_0093_ ), .A2(\us03\/_0056_ ), .B1(\us03\/_0134_ ), .B2(\us03\/_0114_ ), .Y(\us03\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1267_ ( .A1(\us03\/_0161_ ), .A2(\us03\/_0032_ ), .B1(\us03\/_0324_ ), .B2(\us03\/_0147_ ), .Y(\us03\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1268_ ( .A1(\us03\/_0054_ ), .A2(\us03\/_0732_ ), .B1(\us03\/_0748_ ), .B2(\us03\/_0304_ ), .Y(\us03\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1269_ ( .A(\us03\/_0477_ ), .B(\us03\/_0479_ ), .C(\us03\/_0480_ ), .D(\us03\/_0481_ ), .X(\us03\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1270_ ( .A(\us03\/_0161_ ), .B(\us03\/_0064_ ), .Y(\us03\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us03/_1271_ ( .A(\us03\/_0732_ ), .B(\us03\/_0123_ ), .C(\us03\/_0467_ ), .Y(\us03\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1272_ ( .A(\us03\/_0483_ ), .B(\us03\/_0484_ ), .Y(\us03\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1273_ ( .A(\us03\/_0297_ ), .Y(\us03\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us03/_1274_ ( .A_N(\us03\/_0485_ ), .B(\us03\/_0181_ ), .C(\us03\/_0486_ ), .D(\us03\/_0386_ ), .X(\us03\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1275_ ( .A(\us03\/_0472_ ), .B(\us03\/_0476_ ), .C(\us03\/_0482_ ), .D(\us03\/_0487_ ), .X(\us03\/_0488_ ) );
sky130_fd_sc_hd__nand3_2 \us03/_1276_ ( .A(\us03\/_0440_ ), .B(\us03\/_0462_ ), .C(\us03\/_0488_ ), .Y(\us03\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1277_ ( .A(\us03\/_0403_ ), .B(\us03\/_0230_ ), .C(\us03\/_0451_ ), .D(\us03\/_0361_ ), .X(\us03\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1278_ ( .A1(\us03\/_0118_ ), .A2(\us03\/_0050_ ), .B1(\us03\/_0109_ ), .C1(\us03\/_0139_ ), .Y(\us03\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1279_ ( .A(\us03\/_0447_ ), .B(\us03\/_0437_ ), .C(\us03\/_0491_ ), .D(\us03\/_0427_ ), .X(\us03\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1280_ ( .A1(\us03\/_0280_ ), .A2(\us03\/_0255_ ), .B1(\us03\/_0608_ ), .B2(\us03\/_0247_ ), .Y(\us03\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1281_ ( .A1(\us03\/_0144_ ), .A2(\us03\/_0147_ ), .B1(\us03\/_0355_ ), .B2(\us03\/_0093_ ), .Y(\us03\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1282_ ( .A1(\us03\/_0705_ ), .A2(\us03\/_0279_ ), .B1(\us03\/_0330_ ), .B2(\us03\/_0247_ ), .Y(\us03\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1283_ ( .A1(\us03\/_0279_ ), .A2(\us03\/_0280_ ), .B1(\us03\/_0114_ ), .Y(\us03\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1284_ ( .A(\us03\/_0493_ ), .B(\us03\/_0494_ ), .C(\us03\/_0495_ ), .D(\us03\/_0496_ ), .X(\us03\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1285_ ( .A1(\us03\/_0134_ ), .A2(\us03\/_0137_ ), .B1(\us03\/_0355_ ), .B2(\us03\/_0575_ ), .Y(\us03\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1286_ ( .A1(\us03\/_0364_ ), .A2(\us03\/_0733_ ), .B1(\us03\/_0093_ ), .B2(\us03\/_0499_ ), .Y(\us03\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1287_ ( .A(\us03\/_0147_ ), .B(\us03\/_0640_ ), .Y(\us03\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1288_ ( .A1(\us03\/_0153_ ), .A2(\us03\/_0056_ ), .B1(\us03\/_0748_ ), .Y(\us03\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1289_ ( .A(\us03\/_0498_ ), .B(\us03\/_0500_ ), .C(\us03\/_0501_ ), .D(\us03\/_0502_ ), .X(\us03\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1290_ ( .A(\us03\/_0490_ ), .B(\us03\/_0492_ ), .C(\us03\/_0497_ ), .D(\us03\/_0503_ ), .X(\us03\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us03/_1291_ ( .A_N(\us03\/_0275_ ), .B(\us03\/_0705_ ), .X(\us03\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1292_ ( .A(\us03\/_0505_ ), .Y(\us03\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1293_ ( .A(\us03\/_0380_ ), .B(\us03\/_0347_ ), .X(\us03\/_0507_ ) );
sky130_fd_sc_hd__o21ai_1 \us03/_1294_ ( .A1(\us03\/_0507_ ), .A2(\us03\/_0093_ ), .B1(\us03\/_0056_ ), .Y(\us03\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1295_ ( .A(\us03\/_0322_ ), .B(\us03\/_0277_ ), .C(\us03\/_0506_ ), .D(\us03\/_0508_ ), .X(\us03\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1296_ ( .A(\us03\/_0280_ ), .B(\us03\/_0705_ ), .X(\us03\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1297_ ( .A1(\us03\/_0733_ ), .A2(\us03\/_0114_ ), .B1(\us03\/_0429_ ), .C1(\us03\/_0511_ ), .Y(\us03\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_1298_ ( .A(\us03\/_0019_ ), .B(\us03\/_0024_ ), .Y(\us03\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1299_ ( .A(\us03\/_0512_ ), .B(\us03\/_0513_ ), .C(\us03\/_0742_ ), .D(\us03\/_0306_ ), .X(\us03\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1300_ ( .A1(\us03\/_0532_ ), .A2(\us03\/_0089_ ), .B1(\us03\/_0154_ ), .C1(\us03\/_0169_ ), .Y(\us03\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us03/_1301_ ( .A1(\us03\/_0749_ ), .A2(\us03\/_0026_ ), .B1(\us03\/_0069_ ), .C1(\us03\/_0032_ ), .X(\us03\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us03/_1302_ ( .A1(\us03\/_0324_ ), .A2(\us03\/_0355_ ), .B1(\us03\/_0330_ ), .B2(\us03\/_0727_ ), .X(\us03\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us03/_1303_ ( .A(\us03\/_0133_ ), .B(\us03\/_0516_ ), .C(\us03\/_0517_ ), .Y(\us03\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1304_ ( .A(\us03\/_0509_ ), .B(\us03\/_0514_ ), .C(\us03\/_0515_ ), .D(\us03\/_0518_ ), .X(\us03\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1305_ ( .A(\us03\/_0747_ ), .B(\us03\/_0072_ ), .Y(\us03\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1306_ ( .A1(\us03\/_0082_ ), .A2(\us03\/_0070_ ), .B1(\us03\/_0043_ ), .B2(\us03\/_0193_ ), .Y(\us03\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1307_ ( .A(\us03\/_0311_ ), .B(\us03\/_0520_ ), .C(\us03\/_0332_ ), .D(\us03\/_0522_ ), .X(\us03\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1308_ ( .A(\us03\/_0129_ ), .B(\us03\/_0499_ ), .X(\us03\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_1309_ ( .A(\us03\/_0235_ ), .B(\us03\/_0524_ ), .Y(\us03\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us03/_1310_ ( .A(\us03\/_0081_ ), .B(\us03\/_0085_ ), .Y(\us03\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1311_ ( .A1(\us03\/_0051_ ), .A2(\us03\/_0045_ ), .B1(\us03\/_0130_ ), .B2(\us03\/_0094_ ), .Y(\us03\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1312_ ( .A(\us03\/_0523_ ), .B(\us03\/_0525_ ), .C(\us03\/_0526_ ), .D(\us03\/_0527_ ), .X(\us03\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us03/_1313_ ( .A_N(\us03\/_0250_ ), .B(\us03\/_0521_ ), .Y(\us03\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1314_ ( .A(\us03\/_0128_ ), .B(\us03\/_0020_ ), .X(\us03\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1315_ ( .A(\us03\/_0530_ ), .Y(\us03\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1316_ ( .A(\us03\/_0364_ ), .B(\us03\/_0058_ ), .X(\us03\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1317_ ( .A(\us03\/_0533_ ), .Y(\us03\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us03/_1318_ ( .A_N(\us03\/_0529_ ), .B(\us03\/_0531_ ), .C(\us03\/_0534_ ), .D(\us03\/_0192_ ), .X(\us03\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1319_ ( .A(\us03\/_0434_ ), .B(\us03\/_0078_ ), .X(\us03\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us03/_1320_ ( .A1(\us03\/_0750_ ), .A2(\us03\/_0079_ ), .B1(\us03\/_0129_ ), .B2(\us03\/_0705_ ), .X(\us03\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1321_ ( .A1(\us03\/_0161_ ), .A2(\us03\/_0032_ ), .B1(\us03\/_0536_ ), .C1(\us03\/_0537_ ), .Y(\us03\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us03/_1322_ ( .A1(\us03\/_0747_ ), .A2(\us03\/_0162_ ), .B1(\us03\/_0079_ ), .B2(\us03\/_0043_ ), .X(\us03\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1323_ ( .A1(\us03\/_0093_ ), .A2(\us03\/_0247_ ), .B1(\us03\/_0240_ ), .C1(\us03\/_0539_ ), .Y(\us03\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1324_ ( .A(\us03\/_0434_ ), .B(\us03\/_0043_ ), .X(\us03\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us03/_1325_ ( .A1(\us03\/_0142_ ), .A2(\us03\/_0150_ ), .B1(\us03\/_0022_ ), .B2(\us03\/_0137_ ), .X(\us03\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1326_ ( .A1(\us03\/_0279_ ), .A2(\us03\/_0051_ ), .B1(\us03\/_0541_ ), .C1(\us03\/_0542_ ), .Y(\us03\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1327_ ( .A(\us03\/_0159_ ), .B(\us03\/_0036_ ), .X(\us03\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us03/_1328_ ( .A1(\us03\/_0271_ ), .A2(\us03\/_0434_ ), .B1(\us03\/_0028_ ), .X(\us03\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1329_ ( .A1(\us03\/_0091_ ), .A2(\us03\/_0128_ ), .B1(\us03\/_0545_ ), .C1(\us03\/_0546_ ), .Y(\us03\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1330_ ( .A(\us03\/_0538_ ), .B(\us03\/_0540_ ), .C(\us03\/_0544_ ), .D(\us03\/_0547_ ), .X(\us03\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1331_ ( .A(\us03\/_0364_ ), .B(\us03\/_0193_ ), .X(\us03\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us03/_1332_ ( .A(\us03\/_0549_ ), .B(\us03\/_0186_ ), .C(\us03\/_0187_ ), .Y(\us03\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1333_ ( .A(\us03\/_0062_ ), .B(\us03\/_0347_ ), .C(\us03\/_0749_ ), .D(\us03\/_0694_ ), .X(\us03\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1334_ ( .A1(\us03\/_0130_ ), .A2(\us03\/_0499_ ), .B1(\us03\/_0551_ ), .C1(\us03\/_0101_ ), .Y(\us03\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1335_ ( .A(\us03\/_0139_ ), .B(\us03\/_0640_ ), .Y(\us03\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1336_ ( .A1(\us03\/_0752_ ), .A2(\us03\/_0672_ ), .B1(\us03\/_0280_ ), .B2(\us03\/_0364_ ), .Y(\us03\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1337_ ( .A(\us03\/_0550_ ), .B(\us03\/_0552_ ), .C(\us03\/_0553_ ), .D(\us03\/_0555_ ), .X(\us03\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1338_ ( .A(\us03\/_0528_ ), .B(\us03\/_0535_ ), .C(\us03\/_0548_ ), .D(\us03\/_0556_ ), .X(\us03\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us03/_1339_ ( .A(\us03\/_0504_ ), .B(\us03\/_0519_ ), .C(\us03\/_0557_ ), .Y(\us03\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1340_ ( .A(\us03\/_0054_ ), .B(\us03\/_0507_ ), .X(\us03\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us03/_1341_ ( .A_N(\us03\/_0558_ ), .B(\us03\/_0408_ ), .C(\us03\/_0451_ ), .D(\us03\/_0452_ ), .X(\us03\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1342_ ( .A(\us03\/_0549_ ), .Y(\us03\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1343_ ( .A(\us03\/_0559_ ), .B(\us03\/_0403_ ), .C(\us03\/_0560_ ), .D(\us03\/_0371_ ), .X(\us03\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1344_ ( .A(\us03\/_0181_ ), .B(\us03\/_0178_ ), .X(\us03\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1345_ ( .A(\us03\/_0562_ ), .B(\us03\/_0552_ ), .C(\us03\/_0553_ ), .D(\us03\/_0555_ ), .X(\us03\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1346_ ( .A(\us03\/_0247_ ), .B(\us03\/_0020_ ), .Y(\us03\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1347_ ( .A(\us03\/_0051_ ), .B(\us03\/_0130_ ), .X(\us03\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1348_ ( .A(\us03\/_0566_ ), .Y(\us03\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1349_ ( .A(\us03\/_0159_ ), .B(\us03\/_0412_ ), .X(\us03\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1350_ ( .A1(\us03\/_0752_ ), .A2(\us03\/_0640_ ), .B1(\us03\/_0568_ ), .B2(\us03\/_0175_ ), .Y(\us03\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1351_ ( .A(\us03\/_0076_ ), .B(\us03\/_0565_ ), .C(\us03\/_0567_ ), .D(\us03\/_0569_ ), .X(\us03\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us03/_1352_ ( .A1(\us03\/_0036_ ), .A2(\us03\/_0142_ ), .B1(\us03\/_0161_ ), .X(\us03\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1353_ ( .A(\us03\/_0364_ ), .B(\us03\/_0672_ ), .Y(\us03\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us03/_1354_ ( .A(\us03\/_0420_ ), .B(\us03\/_0571_ ), .C_N(\us03\/_0572_ ), .Y(\us03\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1355_ ( .A(\us03\/_0051_ ), .B(\us03\/_0747_ ), .Y(\us03\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1356_ ( .A(\us03\/_0574_ ), .B(\us03\/_0319_ ), .C(\us03\/_0320_ ), .D(\us03\/_0411_ ), .X(\us03\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1357_ ( .A(\us03\/_0736_ ), .B(\us03\/_0035_ ), .Y(\us03\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1358_ ( .A(\us03\/_0736_ ), .B(\us03\/_0030_ ), .Y(\us03\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1359_ ( .A(\us03\/_0298_ ), .B(\us03\/_0208_ ), .C(\us03\/_0577_ ), .D(\us03\/_0578_ ), .X(\us03\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1360_ ( .A1(\us03\/_0020_ ), .A2(\us03\/_0137_ ), .B1(\us03\/_0261_ ), .B2(\us03\/_0128_ ), .Y(\us03\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1361_ ( .A(\us03\/_0573_ ), .B(\us03\/_0576_ ), .C(\us03\/_0579_ ), .D(\us03\/_0580_ ), .X(\us03\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1362_ ( .A(\us03\/_0561_ ), .B(\us03\/_0563_ ), .C(\us03\/_0570_ ), .D(\us03\/_0581_ ), .X(\us03\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1363_ ( .A(\us03\/_0128_ ), .B(\us03\/_0193_ ), .X(\us03\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1364_ ( .A(\us03\/_0082_ ), .B(\us03\/_0162_ ), .X(\us03\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us03/_1365_ ( .A(\us03\/_0583_ ), .B(\us03\/_0584_ ), .C_N(\us03\/_0437_ ), .Y(\us03\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us03/_1366_ ( .A(\us03\/_0150_ ), .B(\us03\/_0118_ ), .C(\us03\/_0380_ ), .Y(\us03\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us03/_1367_ ( .A_N(\us03\/_0182_ ), .B(\us03\/_0587_ ), .C(\us03\/_0323_ ), .X(\us03\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1368_ ( .A1(\us03\/_0575_ ), .A2(\us03\/_0153_ ), .B1(\us03\/_0727_ ), .B2(\us03\/_0058_ ), .Y(\us03\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1369_ ( .A1(\us03\/_0499_ ), .A2(\us03\/_0064_ ), .B1(\us03\/_0134_ ), .B2(\us03\/_0255_ ), .Y(\us03\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1370_ ( .A(\us03\/_0585_ ), .B(\us03\/_0588_ ), .C(\us03\/_0589_ ), .D(\us03\/_0590_ ), .X(\us03\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us03/_1371_ ( .A1(\us03\/_0091_ ), .A2(\us03\/_0139_ ), .B1(\us03\/_0250_ ), .Y(\us03\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1372_ ( .A1(\us03\/_0092_ ), .A2(\us03\/_0739_ ), .B1(\us03\/_0324_ ), .B2(\us03\/_0247_ ), .Y(\us03\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1373_ ( .A1(\us03\/_0144_ ), .A2(\us03\/_0153_ ), .B1(\us03\/_0683_ ), .B2(\us03\/_0056_ ), .Y(\us03\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1374_ ( .A1(\us03\/_0091_ ), .A2(\us03\/_0499_ ), .B1(\us03\/_0330_ ), .B2(\us03\/_0056_ ), .Y(\us03\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1375_ ( .A(\us03\/_0592_ ), .B(\us03\/_0593_ ), .C(\us03\/_0594_ ), .D(\us03\/_0595_ ), .X(\us03\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1376_ ( .A(\us03\/_0499_ ), .B(\us03\/_0144_ ), .Y(\us03\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1377_ ( .A(\us03\/_0312_ ), .B(\us03\/_0598_ ), .Y(\us03\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1378_ ( .A(\us03\/_0575_ ), .B(\us03\/_0147_ ), .Y(\us03\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1379_ ( .A1(\us03\/_0293_ ), .A2(\us03\/_0137_ ), .B1(\us03\/_0093_ ), .B2(\us03\/_0739_ ), .Y(\us03\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1380_ ( .A1(\us03\/_0734_ ), .A2(\us03\/_0531_ ), .B1(\us03\/_0600_ ), .C1(\us03\/_0601_ ), .Y(\us03\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1381_ ( .A1(\us03\/_0153_ ), .A2(\us03\/_0261_ ), .B1(\us03\/_0599_ ), .C1(\us03\/_0602_ ), .Y(\us03\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1382_ ( .A(\us03\/_0591_ ), .B(\us03\/_0596_ ), .C(\us03\/_0174_ ), .D(\us03\/_0603_ ), .X(\us03\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1383_ ( .A(\us03\/_0247_ ), .B(\us03\/_0144_ ), .Y(\us03\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1384_ ( .A(\us03\/_0113_ ), .B(\us03\/_0018_ ), .Y(\us03\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1385_ ( .A(\us03\/_0381_ ), .B(\us03\/_0605_ ), .C(\us03\/_0361_ ), .D(\us03\/_0606_ ), .X(\us03\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1386_ ( .A1(\us03\/_0016_ ), .A2(\us03\/_0727_ ), .B1(\us03\/_0733_ ), .Y(\us03\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1387_ ( .A1(\us03\/_0586_ ), .A2(\us03\/_0159_ ), .B1(\us03\/_0082_ ), .B2(\us03\/_0750_ ), .Y(\us03\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1388_ ( .A1(\us03\/_0142_ ), .A2(\us03\/_0162_ ), .B1(\us03\/_0079_ ), .B2(\us03\/_0054_ ), .Y(\us03\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1389_ ( .A(\us03\/_0610_ ), .B(\us03\/_0611_ ), .C(\us03\/_0105_ ), .D(\us03\/_0106_ ), .X(\us03\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1390_ ( .A1(\us03\/_0094_ ), .A2(\us03\/_0302_ ), .B1(\us03\/_0324_ ), .B2(\us03\/_0089_ ), .Y(\us03\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1391_ ( .A(\us03\/_0607_ ), .B(\us03\/_0609_ ), .C(\us03\/_0612_ ), .D(\us03\/_0613_ ), .X(\us03\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1392_ ( .A(\us03\/_0041_ ), .B(\us03\/_0170_ ), .X(\us03\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1393_ ( .A(\us03\/_0554_ ), .B(\us03\/_0028_ ), .X(\us03\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1394_ ( .A(\us03\/_0028_ ), .B(\us03\/_0261_ ), .Y(\us03\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us03/_1395_ ( .A_N(\us03\/_0616_ ), .B(\us03\/_0617_ ), .Y(\us03\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1396_ ( .A1(\us03\/_0147_ ), .A2(\us03\/_0302_ ), .B1(\us03\/_0342_ ), .C1(\us03\/_0618_ ), .Y(\us03\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1397_ ( .A(\us03\/_0614_ ), .B(\us03\/_0272_ ), .C(\us03\/_0615_ ), .D(\us03\/_0620_ ), .X(\us03\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us03/_1398_ ( .A(\us03\/_0582_ ), .B(\us03\/_0604_ ), .C(\us03\/_0621_ ), .Y(\us03\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1399_ ( .A1(\us03\/_0280_ ), .A2(\us03\/_0134_ ), .B1(\us03\/_0089_ ), .Y(\us03\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1400_ ( .A1(\us03\/_0144_ ), .A2(\us03\/_0608_ ), .A3(\us03\/_0330_ ), .B1(\us03\/_0089_ ), .Y(\us03\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1401_ ( .A1(\us03\/_0197_ ), .A2(\us03\/_0130_ ), .A3(\us03\/_0110_ ), .B1(\us03\/_0094_ ), .Y(\us03\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1402_ ( .A(\us03\/_0432_ ), .B(\us03\/_0622_ ), .C(\us03\/_0623_ ), .D(\us03\/_0624_ ), .X(\us03\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us03/_1403_ ( .A1(\us03\/_0554_ ), .A2(\us03\/_0018_ ), .A3(\us03\/_0022_ ), .B1(\us03\/_0161_ ), .X(\us03\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us03/_1404_ ( .A_N(\us03\/_0269_ ), .B(\us03\/_0170_ ), .X(\us03\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1405_ ( .A1(\us03\/_0109_ ), .A2(\us03\/_0064_ ), .A3(\us03\/_0733_ ), .B1(\us03\/_0355_ ), .Y(\us03\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us03/_1406_ ( .A_N(\us03\/_0626_ ), .B(\us03\/_0627_ ), .C(\us03\/_0353_ ), .D(\us03\/_0628_ ), .X(\us03\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1407_ ( .A1(\us03\/_0091_ ), .A2(\us03\/_0110_ ), .A3(\us03\/_0176_ ), .B1(\us03\/_0139_ ), .Y(\us03\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1408_ ( .A1(\us03\/_0020_ ), .A2(\us03\/_0261_ ), .B1(\us03\/_0147_ ), .Y(\us03\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1409_ ( .A(\us03\/_0631_ ), .B(\us03\/_0344_ ), .C(\us03\/_0421_ ), .D(\us03\/_0632_ ), .X(\us03\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us03/_1410_ ( .A1(\us03\/_0325_ ), .A2(\us03\/_0734_ ), .B1(\us03\/_0038_ ), .C1(\us03\/_0113_ ), .X(\us03\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1411_ ( .A1(\us03\/_0134_ ), .A2(\us03\/_0114_ ), .B1(\us03\/_0221_ ), .C1(\us03\/_0634_ ), .Y(\us03\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us03/_1412_ ( .A(\us03\/_0119_ ), .B_N(\us03\/_0111_ ), .Y(\us03\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1413_ ( .A1(\us03\/_0032_ ), .A2(\us03\/_0113_ ), .B1(\us03\/_0636_ ), .C1(\us03\/_0400_ ), .Y(\us03\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1414_ ( .A1(\us03\/_0732_ ), .A2(\us03\/_0293_ ), .A3(\us03\/_0251_ ), .B1(\us03\/_0364_ ), .Y(\us03\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1415_ ( .A(\us03\/_0189_ ), .B(\us03\/_0635_ ), .C(\us03\/_0637_ ), .D(\us03\/_0638_ ), .X(\us03\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1416_ ( .A(\us03\/_0625_ ), .B(\us03\/_0630_ ), .C(\us03\/_0633_ ), .D(\us03\/_0639_ ), .X(\us03\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1417_ ( .A(\us03\/_0747_ ), .B(\us03\/_0738_ ), .X(\us03\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1418_ ( .A(\us03\/_0736_ ), .B(\us03\/_0731_ ), .X(\us03\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us03/_1419_ ( .A_N(\us03\/_0643_ ), .B(\us03\/_0577_ ), .Y(\us03\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1420_ ( .A1(\us03\/_0280_ ), .A2(\us03\/_0739_ ), .B1(\us03\/_0642_ ), .C1(\us03\/_0644_ ), .Y(\us03\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1421_ ( .A1(\us03\/_0050_ ), .A2(\us03\/_0543_ ), .B1(\us03\/_0194_ ), .C1(\us03\/_0738_ ), .Y(\us03\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1422_ ( .A(\us03\/_0646_ ), .B(\us03\/_0232_ ), .C(\us03\/_0417_ ), .D(\us03\/_0578_ ), .X(\us03\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1423_ ( .A1(\us03\/_0064_ ), .A2(\us03\/_0733_ ), .B1(\us03\/_0727_ ), .Y(\us03\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1424_ ( .A1(\us03\/_0193_ ), .A2(\us03\/_0276_ ), .B1(\us03\/_0727_ ), .Y(\us03\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1425_ ( .A(\us03\/_0645_ ), .B(\us03\/_0647_ ), .C(\us03\/_0648_ ), .D(\us03\/_0649_ ), .X(\us03\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1426_ ( .A1(\us03\/_0325_ ), .A2(\us03\/_0734_ ), .B1(\us03\/_0038_ ), .C1(\us03\/_0247_ ), .Y(\us03\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1427_ ( .A1(\us03\/_0543_ ), .A2(\us03\/_0216_ ), .B1(\us03\/_0412_ ), .C1(\us03\/_0247_ ), .Y(\us03\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1428_ ( .A(\us03\/_0652_ ), .B(\us03\/_0653_ ), .X(\us03\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1429_ ( .A1(\us03\/_0733_ ), .A2(\us03\/_0748_ ), .A3(\us03\/_0324_ ), .B1(\us03\/_0016_ ), .Y(\us03\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1430_ ( .A1(\us03\/_0640_ ), .A2(\us03\/_0193_ ), .A3(\us03\/_0091_ ), .B1(\us03\/_0016_ ), .Y(\us03\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1431_ ( .A1(\us03\/_0102_ ), .A2(\us03\/_0301_ ), .B1(\sa03\[3\] ), .C1(\us03\/_0247_ ), .Y(\us03\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1432_ ( .A(\us03\/_0654_ ), .B(\us03\/_0655_ ), .C(\us03\/_0656_ ), .D(\us03\/_0657_ ), .X(\us03\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1433_ ( .A1(\us03\/_0118_ ), .A2(\us03\/_0050_ ), .B1(\us03\/_0038_ ), .C1(\us03\/_0489_ ), .Y(\us03\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us03/_1434_ ( .A_N(\us03\/_0250_ ), .B(\us03\/_0465_ ), .C(\us03\/_0659_ ), .X(\us03\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1435_ ( .A1(\us03\/_0683_ ), .A2(\us03\/_0324_ ), .B1(\us03\/_0255_ ), .Y(\us03\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1436_ ( .A1(\us03\/_0032_ ), .A2(\us03\/_0193_ ), .A3(\us03\/_0048_ ), .B1(\us03\/_0255_ ), .Y(\us03\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1437_ ( .A1(\us03\/_0144_ ), .A2(\us03\/_0586_ ), .A3(\us03\/_0048_ ), .B1(\us03\/_0499_ ), .Y(\us03\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1438_ ( .A(\us03\/_0660_ ), .B(\us03\/_0661_ ), .C(\us03\/_0663_ ), .D(\us03\/_0664_ ), .X(\us03\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1439_ ( .A1(\us03\/_0091_ ), .A2(\us03\/_0276_ ), .B1(\us03\/_0060_ ), .Y(\us03\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1440_ ( .A1(\us03\/_0144_ ), .A2(\us03\/_0608_ ), .B1(\us03\/_0056_ ), .Y(\us03\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1441_ ( .A1(\us03\/_0412_ ), .A2(\us03\/_0038_ ), .B1(\us03\/_0102_ ), .C1(\us03\/_0060_ ), .Y(\us03\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1442_ ( .A1(\sa03\[1\] ), .A2(\us03\/_0734_ ), .B1(\us03\/_0109_ ), .C1(\us03\/_0056_ ), .Y(\us03\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1443_ ( .A(\us03\/_0666_ ), .B(\us03\/_0667_ ), .C(\us03\/_0668_ ), .D(\us03\/_0669_ ), .X(\us03\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1444_ ( .A(\us03\/_0650_ ), .B(\us03\/_0658_ ), .C(\us03\/_0665_ ), .D(\us03\/_0670_ ), .X(\us03\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us03/_1445_ ( .A(\us03\/_0641_ ), .B(\us03\/_0174_ ), .C(\us03\/_0671_ ), .Y(\us03\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us03/_1446_ ( .A(\us03\/_0049_ ), .B(\us03\/_0618_ ), .C_N(\us03\/_0052_ ), .Y(\us03\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us03/_1447_ ( .A(\us03\/_0239_ ), .Y(\us03\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1448_ ( .A(\us03\/_0705_ ), .B(\us03\/_0032_ ), .Y(\us03\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1449_ ( .A1(\us03\/_0054_ ), .A2(\us03\/_0732_ ), .B1(\us03\/_0036_ ), .B2(\us03\/_0705_ ), .Y(\us03\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1450_ ( .A1(\us03\/_0304_ ), .A2(\us03\/_0732_ ), .B1(\us03\/_0048_ ), .B2(\us03\/_0750_ ), .Y(\us03\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1451_ ( .A(\us03\/_0674_ ), .B(\us03\/_0675_ ), .C(\us03\/_0676_ ), .D(\us03\/_0677_ ), .X(\us03\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us03/_1452_ ( .A_N(\us03\/_0584_ ), .B(\us03\/_0283_ ), .X(\us03\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1453_ ( .A(\us03\/_0673_ ), .B(\us03\/_0678_ ), .C(\us03\/_0679_ ), .D(\us03\/_0508_ ), .X(\us03\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1454_ ( .A1(\us03\/_0016_ ), .A2(\us03\/_0733_ ), .B1(\us03\/_0355_ ), .B2(\us03\/_0092_ ), .Y(\us03\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1455_ ( .A(\us03\/_0681_ ), .B(\us03\/_0034_ ), .X(\us03\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us03/_1456_ ( .A1(\us03\/_0330_ ), .A2(\us03\/_0139_ ), .B1(\us03\/_0324_ ), .B2(\us03\/_0089_ ), .X(\us03\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1457_ ( .A1(\us03\/_0146_ ), .A2(\us03\/_0147_ ), .B1(\us03\/_0133_ ), .C1(\us03\/_0684_ ), .Y(\us03\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1458_ ( .A(\us03\/_0113_ ), .B(\us03\/_0251_ ), .Y(\us03\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us03/_1459_ ( .A_N(\us03\/_0463_ ), .B(\us03\/_0686_ ), .C(\us03\/_0383_ ), .D(\us03\/_0464_ ), .X(\us03\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1460_ ( .A1(\us03\/_0051_ ), .A2(\us03\/_0293_ ), .B1(\us03\/_0280_ ), .B2(\us03\/_0705_ ), .Y(\us03\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1461_ ( .A1(\us03\/_0018_ ), .A2(\us03\/_0072_ ), .B1(\us03\/_0134_ ), .B2(\us03\/_0078_ ), .Y(\us03\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1462_ ( .A(\us03\/_0687_ ), .B(\us03\/_0236_ ), .C(\us03\/_0688_ ), .D(\us03\/_0689_ ), .X(\us03\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1463_ ( .A(\us03\/_0680_ ), .B(\us03\/_0682_ ), .C(\us03\/_0685_ ), .D(\us03\/_0690_ ), .X(\us03\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us03/_1464_ ( .A1(\us03\/_0532_ ), .A2(\us03\/_0380_ ), .B1(\us03\/_0102_ ), .C1(\us03\/_0355_ ), .X(\us03\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us03/_1465_ ( .A(\us03\/_0692_ ), .B(\us03\/_0338_ ), .C(\us03\/_0644_ ), .Y(\us03\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1466_ ( .A(\us03\/_0016_ ), .B(\us03\/_0020_ ), .Y(\us03\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1467_ ( .A1(\us03\/_0032_ ), .A2(\us03\/_0137_ ), .B1(\us03\/_0279_ ), .B2(\us03\/_0094_ ), .Y(\us03\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1468_ ( .A1(\us03\/_0575_ ), .A2(\us03\/_0153_ ), .B1(\us03\/_0161_ ), .B2(\us03\/_0293_ ), .Y(\us03\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1469_ ( .A(\us03\/_0259_ ), .B(\us03\/_0695_ ), .C(\us03\/_0696_ ), .D(\us03\/_0697_ ), .X(\us03\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us03/_1470_ ( .A1(\us03\/_0255_ ), .A2(\us03\/_0640_ ), .B1(\us03\/_0016_ ), .B2(\us03\/_0193_ ), .X(\us03\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1471_ ( .A1(\us03\/_0060_ ), .A2(\us03\/_0176_ ), .B1(\us03\/_0699_ ), .C1(\us03\/_0177_ ), .Y(\us03\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1472_ ( .A1(\us03\/_0091_ ), .A2(\us03\/_0499_ ), .B1(\us03\/_0092_ ), .B2(\us03\/_0705_ ), .Y(\us03\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us03/_1473_ ( .A1(\us03\/_0705_ ), .A2(\us03\/_0683_ ), .B1(\us03\/_0093_ ), .B2(\us03\/_0114_ ), .Y(\us03\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us03/_1474_ ( .A1(\us03\/_0683_ ), .A2(\us03\/_0280_ ), .B1(\us03\/_0094_ ), .Y(\us03\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us03/_1475_ ( .A1(\us03\/_0543_ ), .A2(\us03\/_0216_ ), .B1(\us03\/_0038_ ), .C1(\us03\/_0056_ ), .Y(\us03\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1476_ ( .A(\us03\/_0701_ ), .B(\us03\/_0702_ ), .C(\us03\/_0703_ ), .D(\us03\/_0704_ ), .X(\us03\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1477_ ( .A(\us03\/_0693_ ), .B(\us03\/_0698_ ), .C(\us03\/_0700_ ), .D(\us03\/_0706_ ), .X(\us03\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us03/_1478_ ( .A1(\us03\/_0113_ ), .A2(\us03\/_0640_ ), .B1(\us03\/_0364_ ), .B2(\us03\/_0058_ ), .X(\us03\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us03/_1479_ ( .A(\us03\/_0407_ ), .B(\us03\/_0708_ ), .C(\us03\/_0529_ ), .Y(\us03\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1480_ ( .A(\us03\/_0568_ ), .B(\us03\/_0175_ ), .Y(\us03\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us03/_1481_ ( .A1(\us03\/_0247_ ), .A2(\us03\/_0114_ ), .A3(\us03\/_0051_ ), .B1(\us03\/_0130_ ), .Y(\us03\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1482_ ( .A(\us03\/_0709_ ), .B(\us03\/_0550_ ), .C(\us03\/_0710_ ), .D(\us03\/_0711_ ), .X(\us03\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us03/_1483_ ( .A1(\us03\/_0114_ ), .A2(\us03\/_0064_ ), .B1(\us03\/_0261_ ), .B2(\us03\/_0089_ ), .X(\us03\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1484_ ( .A1(\us03\/_0355_ ), .A2(\us03\/_0261_ ), .B1(\us03\/_0198_ ), .C1(\us03\/_0713_ ), .Y(\us03\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1485_ ( .A(\us03\/_0586_ ), .B(\us03\/_0489_ ), .Y(\us03\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us03/_1486_ ( .A_N(\us03\/_0541_ ), .B(\us03\/_0267_ ), .C(\us03\/_0715_ ), .D(\us03\/_0320_ ), .X(\us03\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1487_ ( .A(\us03\/_0586_ ), .B(\us03\/_0070_ ), .Y(\us03\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us03/_1488_ ( .A_N(\us03\/_0211_ ), .B(\us03\/_0155_ ), .C(\us03\/_0202_ ), .D(\us03\/_0718_ ), .X(\us03\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us03/_1489_ ( .A(\us03\/_0150_ ), .B(\us03\/_0216_ ), .C(\us03\/_0380_ ), .Y(\us03\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us03/_1490_ ( .A(\us03\/_0411_ ), .B(\us03\/_0720_ ), .X(\us03\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us03/_1491_ ( .A1(\us03\/_0018_ ), .A2(\us03\/_0022_ ), .B1(\us03\/_0078_ ), .X(\us03\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us03/_1492_ ( .A1(\us03\/_0134_ ), .A2(\us03\/_0738_ ), .B1(\us03\/_0101_ ), .C1(\us03\/_0722_ ), .Y(\us03\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1493_ ( .A(\us03\/_0717_ ), .B(\us03\/_0719_ ), .C(\us03\/_0721_ ), .D(\us03\/_0723_ ), .X(\us03\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us03/_1494_ ( .A(\us03\/_0739_ ), .B(\us03\/_0193_ ), .Y(\us03\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1495_ ( .A(\us03\/_0344_ ), .B(\us03\/_0184_ ), .C(\us03\/_0449_ ), .D(\us03\/_0725_ ), .X(\us03\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us03/_1496_ ( .A(\us03\/_0712_ ), .B(\us03\/_0714_ ), .C(\us03\/_0724_ ), .D(\us03\/_0726_ ), .X(\us03\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \us03/_1497_ ( .A(\us03\/_0691_ ), .B(\us03\/_0707_ ), .C(\us03\/_0728_ ), .Y(\us03\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \us10/_0753_ ( .A(\sa10\[2\] ), .B_N(\sa10\[3\] ), .Y(\us10\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0755_ ( .A(\sa10\[1\] ), .B(\sa10\[0\] ), .X(\us10\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0756_ ( .A(\us10\/_0096_ ), .B(\us10\/_0118_ ), .X(\us10\/_0129_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0757_ ( .A(\sa10\[7\] ), .B(\sa10\[6\] ), .X(\us10\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_0758_ ( .A(\sa10\[4\] ), .B(\sa10\[5\] ), .Y(\us10\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0759_ ( .A(\us10\/_0140_ ), .B(\us10\/_0151_ ), .X(\us10\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0761_ ( .A(\us10\/_0129_ ), .B(\us10\/_0162_ ), .X(\us10\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0762_ ( .A(\us10\/_0096_ ), .X(\us10\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \us10/_0763_ ( .A(\sa10\[1\] ), .B_N(\sa10\[0\] ), .Y(\us10\/_0205_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0764_ ( .A(\us10\/_0205_ ), .X(\us10\/_0216_ ) );
sky130_fd_sc_hd__and3_1 \us10/_0765_ ( .A(\us10\/_0162_ ), .B(\us10\/_0194_ ), .C(\us10\/_0216_ ), .X(\us10\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us10/_0766_ ( .A(\us10\/_0183_ ), .SLEEP(\us10\/_0227_ ), .X(\us10\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \us10/_0767_ ( .A(\sa10\[0\] ), .B_N(\sa10\[1\] ), .Y(\us10\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_0768_ ( .A(\sa10\[2\] ), .B(\sa10\[3\] ), .Y(\us10\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0769_ ( .A(\us10\/_0249_ ), .B(\us10\/_0260_ ), .X(\us10\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0770_ ( .A(\us10\/_0271_ ), .X(\us10\/_0282_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0771_ ( .A(\us10\/_0282_ ), .X(\us10\/_0293_ ) );
sky130_fd_sc_hd__buf_2 \us10/_0772_ ( .A(\us10\/_0162_ ), .X(\us10\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_0773_ ( .A(\us10\/_0293_ ), .B(\us10\/_0304_ ), .Y(\us10\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us10/_0774_ ( .A(\sa10\[1\] ), .Y(\us10\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us10/_0776_ ( .A(\sa10\[0\] ), .Y(\us10\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0777_ ( .A(\sa10\[2\] ), .B(\sa10\[3\] ), .X(\us10\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0779_ ( .A(\us10\/_0358_ ), .X(\us10\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_0780_ ( .A1(\us10\/_0325_ ), .A2(\us10\/_0347_ ), .B1(\us10\/_0380_ ), .C1(\us10\/_0304_ ), .Y(\us10\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us10/_0781_ ( .A_N(\us10\/_0238_ ), .B(\us10\/_0314_ ), .C(\us10\/_0391_ ), .X(\us10\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us10/_0782_ ( .A(\sa10\[3\] ), .B_N(\sa10\[2\] ), .Y(\us10\/_0412_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0783_ ( .A(\us10\/_0412_ ), .X(\us10\/_0423_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0784_ ( .A(\us10\/_0423_ ), .B(\us10\/_0205_ ), .X(\us10\/_0434_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0785_ ( .A(\us10\/_0434_ ), .X(\us10\/_0445_ ) );
sky130_fd_sc_hd__nor2b_1 \us10/_0787_ ( .A(\sa10\[5\] ), .B_N(\sa10\[4\] ), .Y(\us10\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0788_ ( .A(\us10\/_0467_ ), .B(\us10\/_0140_ ), .X(\us10\/_0478_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0789_ ( .A(\us10\/_0478_ ), .X(\us10\/_0489_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_0791_ ( .A(\us10\/_0134_ ), .B(\us10\/_0218_ ), .Y(\us10\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_0792_ ( .A(\us10\/_0489_ ), .B(\us10\/_0282_ ), .Y(\us10\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0793_ ( .A(\us10\/_0194_ ), .X(\us10\/_0532_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0794_ ( .A(\us10\/_0249_ ), .X(\us10\/_0543_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0795_ ( .A(\us10\/_0543_ ), .B(\us10\/_0358_ ), .X(\us10\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0797_ ( .A(\us10\/_0554_ ), .X(\us10\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0798_ ( .A(\us10\/_0216_ ), .B(\us10\/_0358_ ), .X(\us10\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0800_ ( .A(\us10\/_0586_ ), .X(\us10\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_0801_ ( .A1(\us10\/_0532_ ), .A2(\us10\/_0575_ ), .A3(\us10\/_0608_ ), .B1(\us10\/_0218_ ), .Y(\us10\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us10/_0802_ ( .A(\us10\/_0401_ ), .B(\us10\/_0510_ ), .C(\us10\/_0521_ ), .D(\us10\/_0619_ ), .X(\us10\/_0629_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0803_ ( .A(\us10\/_0358_ ), .B(\sa10\[1\] ), .X(\us10\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0805_ ( .A(\us10\/_0205_ ), .B(\us10\/_0260_ ), .X(\us10\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0806_ ( .A(\us10\/_0662_ ), .X(\us10\/_0672_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0807_ ( .A(\us10\/_0672_ ), .X(\us10\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us10/_0808_ ( .A(\sa10\[6\] ), .B_N(\sa10\[7\] ), .Y(\us10\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0809_ ( .A(\us10\/_0467_ ), .B(\us10\/_0694_ ), .X(\us10\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0811_ ( .A(\us10\/_0705_ ), .X(\us10\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_0812_ ( .A1(\us10\/_0640_ ), .A2(\us10\/_0293_ ), .A3(\us10\/_0683_ ), .B1(\us10\/_0727_ ), .Y(\us10\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_0813_ ( .A(\sa10\[1\] ), .B(\sa10\[0\] ), .Y(\us10\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0814_ ( .A(\us10\/_0730_ ), .B(\us10\/_0260_ ), .X(\us10\/_0731_ ) );
sky130_fd_sc_hd__buf_2 \us10/_0815_ ( .A(\us10\/_0731_ ), .X(\us10\/_0732_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0816_ ( .A(\us10\/_0732_ ), .X(\us10\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0817_ ( .A(\sa10\[0\] ), .X(\us10\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us10/_0818_ ( .A1(\us10\/_0325_ ), .A2(\us10\/_0734_ ), .B1(\us10\/_0423_ ), .X(\us10\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0819_ ( .A(\us10\/_0694_ ), .B(\us10\/_0151_ ), .X(\us10\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0821_ ( .A(\us10\/_0736_ ), .X(\us10\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0822_ ( .A(\us10\/_0738_ ), .X(\us10\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_0823_ ( .A1(\us10\/_0733_ ), .A2(\us10\/_0735_ ), .A3(\us10\/_0293_ ), .B1(\us10\/_0739_ ), .Y(\us10\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us10/_0824_ ( .A(\us10\/_0730_ ), .B_N(\us10\/_0358_ ), .Y(\us10\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_0825_ ( .A(\us10\/_0741_ ), .B(\us10\/_0739_ ), .Y(\us10\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_0827_ ( .A1(\us10\/_0118_ ), .A2(\us10\/_0216_ ), .B1(\us10\/_0532_ ), .C1(\us10\/_0739_ ), .Y(\us10\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us10/_0828_ ( .A(\us10\/_0729_ ), .B(\us10\/_0740_ ), .C(\us10\/_0742_ ), .D(\us10\/_0744_ ), .X(\us10\/_0745_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0829_ ( .A(\us10\/_0423_ ), .B(\us10\/_0730_ ), .X(\us10\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0831_ ( .A(\us10\/_0746_ ), .X(\us10\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us10/_0832_ ( .A(\sa10\[4\] ), .B_N(\sa10\[5\] ), .Y(\us10\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0833_ ( .A(\us10\/_0749_ ), .B(\us10\/_0694_ ), .X(\us10\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0835_ ( .A(\us10\/_0750_ ), .X(\us10\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0836_ ( .A(\us10\/_0752_ ), .X(\us10\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0837_ ( .A(\us10\/_0118_ ), .B(\us10\/_0358_ ), .X(\us10\/_0017_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0838_ ( .A(\us10\/_0017_ ), .X(\us10\/_0018_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0839_ ( .A(\us10\/_0752_ ), .B(\us10\/_0018_ ), .X(\us10\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0840_ ( .A(\us10\/_0358_ ), .B(\us10\/_0325_ ), .X(\us10\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0842_ ( .A(\us10\/_0096_ ), .B(\us10\/_0205_ ), .X(\us10\/_0022_ ) );
sky130_fd_sc_hd__buf_2 \us10/_0843_ ( .A(\us10\/_0022_ ), .X(\us10\/_0023_ ) );
sky130_fd_sc_hd__o21a_1 \us10/_0844_ ( .A1(\us10\/_0020_ ), .A2(\us10\/_0023_ ), .B1(\us10\/_0752_ ), .X(\us10\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_0845_ ( .A1(\us10\/_0748_ ), .A2(\us10\/_0016_ ), .B1(\us10\/_0019_ ), .C1(\us10\/_0024_ ), .Y(\us10\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0846_ ( .A(\sa10\[4\] ), .B(\sa10\[5\] ), .X(\us10\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0847_ ( .A(\us10\/_0694_ ), .B(\us10\/_0026_ ), .X(\us10\/_0027_ ) );
sky130_fd_sc_hd__buf_2 \us10/_0849_ ( .A(\us10\/_0027_ ), .X(\us10\/_0029_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0850_ ( .A(\us10\/_0358_ ), .B(\us10\/_0730_ ), .X(\us10\/_0030_ ) );
sky130_fd_sc_hd__buf_2 \us10/_0852_ ( .A(\us10\/_0030_ ), .X(\us10\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_0853_ ( .A(\us10\/_0029_ ), .B(\us10\/_0032_ ), .Y(\us10\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_0854_ ( .A(\us10\/_0029_ ), .B(\us10\/_0735_ ), .Y(\us10\/_0034_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0855_ ( .A(\us10\/_0118_ ), .B(\us10\/_0260_ ), .X(\us10\/_0035_ ) );
sky130_fd_sc_hd__buf_2 \us10/_0856_ ( .A(\us10\/_0035_ ), .X(\us10\/_0036_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0857_ ( .A(\us10\/_0027_ ), .B(\us10\/_0036_ ), .X(\us10\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0858_ ( .A(\us10\/_0260_ ), .X(\us10\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_0859_ ( .A(\us10\/_0038_ ), .B(\us10\/_0347_ ), .Y(\us10\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us10/_0860_ ( .A_N(\us10\/_0039_ ), .B(\us10\/_0027_ ), .X(\us10\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_0861_ ( .A(\us10\/_0037_ ), .B(\us10\/_0040_ ), .Y(\us10\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us10/_0862_ ( .A(\us10\/_0025_ ), .B(\us10\/_0033_ ), .C(\us10\/_0034_ ), .D(\us10\/_0041_ ), .X(\us10\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0863_ ( .A(\us10\/_0749_ ), .B(\us10\/_0140_ ), .X(\us10\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us10/_0865_ ( .A(\sa10\[0\] ), .B(\sa10\[2\] ), .C(\sa10\[3\] ), .X(\us10\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0866_ ( .A(\us10\/_0043_ ), .B(\us10\/_0045_ ), .X(\us10\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0867_ ( .A(\us10\/_0096_ ), .B(\us10\/_0543_ ), .X(\us10\/_0047_ ) );
sky130_fd_sc_hd__buf_2 \us10/_0868_ ( .A(\us10\/_0047_ ), .X(\us10\/_0048_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0869_ ( .A(\us10\/_0048_ ), .B(\us10\/_0043_ ), .X(\us10\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0870_ ( .A(\us10\/_0730_ ), .X(\us10\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0871_ ( .A(\us10\/_0043_ ), .X(\us10\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_0872_ ( .A1(\us10\/_0118_ ), .A2(\us10\/_0050_ ), .B1(\us10\/_0194_ ), .C1(\us10\/_0051_ ), .Y(\us10\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us10/_0873_ ( .A(\us10\/_0046_ ), .B(\us10\/_0049_ ), .C_N(\us10\/_0052_ ), .Y(\us10\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0874_ ( .A(\us10\/_0026_ ), .B(\us10\/_0140_ ), .X(\us10\/_0054_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0875_ ( .A(\us10\/_0054_ ), .X(\us10\/_0055_ ) );
sky130_fd_sc_hd__buf_2 \us10/_0876_ ( .A(\us10\/_0055_ ), .X(\us10\/_0056_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_0877_ ( .A1(\us10\/_0532_ ), .A2(\us10\/_0575_ ), .B1(\us10\/_0056_ ), .Y(\us10\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0878_ ( .A(\us10\/_0423_ ), .B(\us10\/_0325_ ), .X(\us10\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0880_ ( .A(\us10\/_0051_ ), .X(\us10\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_0881_ ( .A1(\us10\/_0732_ ), .A2(\us10\/_0036_ ), .A3(\us10\/_0058_ ), .B1(\us10\/_0060_ ), .Y(\us10\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0882_ ( .A(\us10\/_0260_ ), .B(\sa10\[1\] ), .X(\us10\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0884_ ( .A(\us10\/_0062_ ), .X(\us10\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_0885_ ( .A1(\us10\/_0064_ ), .A2(\us10\/_0748_ ), .A3(\us10\/_0683_ ), .B1(\us10\/_0056_ ), .Y(\us10\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us10/_0886_ ( .A(\us10\/_0053_ ), .B(\us10\/_0057_ ), .C(\us10\/_0061_ ), .D(\us10\/_0065_ ), .X(\us10\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us10/_0887_ ( .A(\us10\/_0629_ ), .B(\us10\/_0745_ ), .C(\us10\/_0042_ ), .D(\us10\/_0066_ ), .X(\us10\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us10/_0889_ ( .A(\sa10\[7\] ), .B_N(\sa10\[6\] ), .Y(\us10\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0890_ ( .A(\us10\/_0069_ ), .B(\us10\/_0151_ ), .X(\us10\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0892_ ( .A(\us10\/_0070_ ), .X(\us10\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_0893_ ( .A1(\us10\/_0129_ ), .A2(\us10\/_0586_ ), .B1(\us10\/_0072_ ), .Y(\us10\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_0894_ ( .A1(\us10\/_0380_ ), .A2(\us10\/_0347_ ), .B1(\us10\/_0194_ ), .B2(\us10\/_0216_ ), .Y(\us10\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us10/_0895_ ( .A(\us10\/_0074_ ), .B_N(\us10\/_0070_ ), .Y(\us10\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us10/_0896_ ( .A(\us10\/_0073_ ), .SLEEP(\us10\/_0075_ ), .X(\us10\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0897_ ( .A(\us10\/_0467_ ), .B(\us10\/_0069_ ), .X(\us10\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0898_ ( .A(\us10\/_0077_ ), .X(\us10\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0899_ ( .A(\us10\/_0412_ ), .B(\us10\/_0118_ ), .X(\us10\/_0079_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0901_ ( .A(\us10\/_0078_ ), .B(\us10\/_0079_ ), .X(\us10\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0902_ ( .A(\us10\/_0412_ ), .B(\us10\/_0249_ ), .X(\us10\/_0082_ ) );
sky130_fd_sc_hd__buf_2 \us10/_0903_ ( .A(\us10\/_0082_ ), .X(\us10\/_0083_ ) );
sky130_fd_sc_hd__buf_2 \us10/_0904_ ( .A(\us10\/_0083_ ), .X(\us10\/_0084_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0905_ ( .A(\us10\/_0084_ ), .B(\us10\/_0078_ ), .X(\us10\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us10/_0906_ ( .A1(\sa10\[0\] ), .A2(\us10\/_0325_ ), .B1(\us10\/_0260_ ), .Y(\us10\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us10/_0907_ ( .A_N(\us10\/_0086_ ), .B(\us10\/_0078_ ), .X(\us10\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us10/_0908_ ( .A(\us10\/_0081_ ), .B(\us10\/_0085_ ), .C(\us10\/_0087_ ), .Y(\us10\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0909_ ( .A(\us10\/_0072_ ), .X(\us10\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_0910_ ( .A1(\us10\/_0733_ ), .A2(\us10\/_0748_ ), .A3(\us10\/_0683_ ), .B1(\us10\/_0089_ ), .Y(\us10\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0911_ ( .A(\us10\/_0129_ ), .X(\us10\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0912_ ( .A(\us10\/_0018_ ), .X(\us10\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0913_ ( .A(\us10\/_0023_ ), .X(\us10\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0914_ ( .A(\us10\/_0078_ ), .X(\us10\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_0915_ ( .A1(\us10\/_0091_ ), .A2(\us10\/_0092_ ), .A3(\us10\/_0093_ ), .B1(\us10\/_0094_ ), .Y(\us10\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us10/_0916_ ( .A(\us10\/_0076_ ), .B(\us10\/_0088_ ), .C(\us10\/_0090_ ), .D(\us10\/_0095_ ), .X(\us10\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0917_ ( .A(\us10\/_0069_ ), .B(\us10\/_0026_ ), .X(\us10\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \us10/_0918_ ( .A(\us10\/_0098_ ), .X(\us10\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0919_ ( .A(\us10\/_0445_ ), .B(\us10\/_0099_ ), .X(\us10\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0920_ ( .A(\us10\/_0079_ ), .B(\us10\/_0098_ ), .X(\us10\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0921_ ( .A(\us10\/_0325_ ), .X(\us10\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_0922_ ( .A1(\us10\/_0102_ ), .A2(\us10\/_0734_ ), .B1(\us10\/_0038_ ), .C1(\us10\/_0099_ ), .Y(\us10\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us10/_0923_ ( .A(\us10\/_0100_ ), .B(\us10\/_0101_ ), .C_N(\us10\/_0103_ ), .Y(\us10\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_0924_ ( .A1(\us10\/_0554_ ), .A2(\us10\/_0586_ ), .B1(\us10\/_0099_ ), .Y(\us10\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_0925_ ( .A(\us10\/_0129_ ), .B(\us10\/_0099_ ), .Y(\us10\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0926_ ( .A(\us10\/_0105_ ), .B(\us10\/_0106_ ), .X(\us10\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0927_ ( .A(\us10\/_0423_ ), .X(\us10\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0928_ ( .A(\us10\/_0260_ ), .B(\sa10\[0\] ), .X(\us10\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0929_ ( .A(\us10\/_0069_ ), .B(\us10\/_0749_ ), .X(\us10\/_0111_ ) );
sky130_fd_sc_hd__buf_2 \us10/_0931_ ( .A(\us10\/_0111_ ), .X(\us10\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0932_ ( .A(\us10\/_0113_ ), .X(\us10\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_0933_ ( .A1(\us10\/_0109_ ), .A2(\us10\/_0110_ ), .B1(\us10\/_0114_ ), .Y(\us10\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us10/_0934_ ( .A(\us10\/_0023_ ), .Y(\us10\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us10/_0935_ ( .A(\us10\/_0554_ ), .Y(\us10\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us10/_0936_ ( .A1(\us10\/_0050_ ), .A2(\us10\/_0118_ ), .B1(\us10\/_0194_ ), .Y(\us10\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us10/_0937_ ( .A(\us10\/_0113_ ), .Y(\us10\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us10/_0938_ ( .A1(\us10\/_0116_ ), .A2(\us10\/_0117_ ), .A3(\us10\/_0119_ ), .B1(\us10\/_0120_ ), .X(\us10\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us10/_0939_ ( .A(\us10\/_0104_ ), .B(\us10\/_0108_ ), .C(\us10\/_0115_ ), .D(\us10\/_0121_ ), .X(\us10\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_0940_ ( .A(\sa10\[7\] ), .B(\sa10\[6\] ), .Y(\us10\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0941_ ( .A(\us10\/_0749_ ), .B(\us10\/_0123_ ), .X(\us10\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0943_ ( .A(\us10\/_0083_ ), .B(\us10\/_0124_ ), .X(\us10\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_0944_ ( .A(\us10\/_0282_ ), .B(\us10\/_0124_ ), .Y(\us10\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0945_ ( .A(\us10\/_0124_ ), .X(\us10\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0946_ ( .A(\us10\/_0260_ ), .B(\us10\/_0325_ ), .X(\us10\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_0948_ ( .A(\us10\/_0128_ ), .B(\us10\/_0130_ ), .Y(\us10\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_0949_ ( .A(\us10\/_0127_ ), .B(\us10\/_0132_ ), .Y(\us10\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us10/_0950_ ( .A(\us10\/_0445_ ), .X(\us10\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_0951_ ( .A(\us10\/_0134_ ), .B(\us10\/_0128_ ), .Y(\us10\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us10/_0952_ ( .A(\us10\/_0126_ ), .B(\us10\/_0133_ ), .C_N(\us10\/_0135_ ), .Y(\us10\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0953_ ( .A(\us10\/_0026_ ), .B(\us10\/_0123_ ), .X(\us10\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0955_ ( .A(\us10\/_0137_ ), .X(\us10\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_0956_ ( .A1(\us10\/_0110_ ), .A2(\us10\/_0293_ ), .A3(\us10\/_0084_ ), .B1(\us10\/_0139_ ), .Y(\us10\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0957_ ( .A(\us10\/_0096_ ), .B(\us10\/_0730_ ), .X(\us10\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0959_ ( .A(\us10\/_0142_ ), .X(\us10\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_0960_ ( .A1(\us10\/_0020_ ), .A2(\us10\/_0144_ ), .A3(\us10\/_0018_ ), .B1(\us10\/_0139_ ), .Y(\us10\/_0145_ ) );
sky130_fd_sc_hd__nor3b_2 \us10/_0961_ ( .A(\sa10\[2\] ), .B(\us10\/_0050_ ), .C_N(\sa10\[3\] ), .Y(\us10\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0962_ ( .A(\us10\/_0128_ ), .X(\us10\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_0963_ ( .A1(\us10\/_0146_ ), .A2(\us10\/_0032_ ), .A3(\us10\/_0640_ ), .B1(\us10\/_0147_ ), .Y(\us10\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us10/_0964_ ( .A(\us10\/_0136_ ), .B(\us10\/_0141_ ), .C(\us10\/_0145_ ), .D(\us10\/_0148_ ), .X(\us10\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0965_ ( .A(\us10\/_0123_ ), .B(\us10\/_0151_ ), .X(\us10\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0967_ ( .A(\us10\/_0150_ ), .X(\us10\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0968_ ( .A(\us10\/_0150_ ), .B(\us10\/_0062_ ), .X(\us10\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_0969_ ( .A(\us10\/_0079_ ), .B(\us10\/_0150_ ), .Y(\us10\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us10/_0970_ ( .A(\us10\/_0150_ ), .B(\us10\/_0423_ ), .C(\us10\/_0543_ ), .Y(\us10\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_0971_ ( .A(\us10\/_0155_ ), .B(\us10\/_0156_ ), .Y(\us10\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_0972_ ( .A1(\us10\/_0153_ ), .A2(\us10\/_0134_ ), .B1(\us10\/_0154_ ), .C1(\us10\/_0157_ ), .Y(\us10\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0973_ ( .A(\us10\/_0467_ ), .B(\us10\/_0123_ ), .X(\us10\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_0975_ ( .A(\us10\/_0159_ ), .X(\us10\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us10/_0976_ ( .A_N(\us10\/_0119_ ), .B(\us10\/_0161_ ), .X(\us10\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us10/_0977_ ( .A(\us10\/_0163_ ), .Y(\us10\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_0978_ ( .A1(\us10\/_0146_ ), .A2(\us10\/_0575_ ), .A3(\us10\/_0608_ ), .B1(\us10\/_0153_ ), .Y(\us10\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_0979_ ( .A1(\us10\/_0062_ ), .A2(\us10\/_0084_ ), .A3(\us10\/_0134_ ), .B1(\us10\/_0161_ ), .Y(\us10\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us10/_0980_ ( .A(\us10\/_0158_ ), .B(\us10\/_0164_ ), .C(\us10\/_0165_ ), .D(\us10\/_0166_ ), .X(\us10\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us10/_0981_ ( .A(\us10\/_0097_ ), .B(\us10\/_0122_ ), .C(\us10\/_0149_ ), .D(\us10\/_0167_ ), .X(\us10\/_0168_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0982_ ( .A(\us10\/_0672_ ), .B(\us10\/_0150_ ), .X(\us10\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_0983_ ( .A(\us10\/_0154_ ), .B(\us10\/_0169_ ), .Y(\us10\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us10/_0984_ ( .A(\us10\/_0123_ ), .B(\us10\/_0151_ ), .C(\us10\/_0038_ ), .X(\us10\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0985_ ( .A(\us10\/_0170_ ), .B(\us10\/_0171_ ), .X(\us10\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \us10/_0986_ ( .A(\us10\/_0172_ ), .Y(\us10\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \us10/_0987_ ( .A(\us10\/_0067_ ), .B(\us10\/_0168_ ), .C(\us10\/_0174_ ), .Y(\us10\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us10/_0988_ ( .A(\sa10\[1\] ), .B(\sa10\[0\] ), .Y(\us10\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us10/_0989_ ( .A(\us10\/_0175_ ), .B(\us10\/_0358_ ), .X(\us10\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0990_ ( .A(\us10\/_0176_ ), .B(\us10\/_0489_ ), .X(\us10\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_0991_ ( .A(\us10\/_0084_ ), .B(\us10\/_0113_ ), .Y(\us10\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0992_ ( .A(\us10\/_0111_ ), .B(\us10\/_0062_ ), .X(\us10\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0993_ ( .A(\us10\/_0111_ ), .B(\us10\/_0672_ ), .X(\us10\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_0994_ ( .A(\us10\/_0179_ ), .B(\us10\/_0180_ ), .Y(\us10\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0995_ ( .A(\us10\/_0055_ ), .B(\us10\/_0058_ ), .X(\us10\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us10/_0996_ ( .A(\us10\/_0182_ ), .Y(\us10\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us10/_0997_ ( .A_N(\us10\/_0177_ ), .B(\us10\/_0178_ ), .C(\us10\/_0181_ ), .D(\us10\/_0184_ ), .X(\us10\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0998_ ( .A(\us10\/_0098_ ), .B(\us10\/_0741_ ), .X(\us10\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us10/_0999_ ( .A(\us10\/_0047_ ), .B(\us10\/_0098_ ), .X(\us10\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us10/_1000_ ( .A(\us10\/_0186_ ), .B(\us10\/_0187_ ), .X(\us10\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1001_ ( .A(\us10\/_0188_ ), .Y(\us10\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1002_ ( .A(\us10\/_0738_ ), .B(\us10\/_0735_ ), .X(\us10\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1003_ ( .A(\us10\/_0282_ ), .B(\us10\/_0736_ ), .X(\us10\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_1004_ ( .A(\us10\/_0190_ ), .B(\us10\/_0191_ ), .Y(\us10\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us10/_1005_ ( .A(\us10\/_0096_ ), .B(\us10\/_0325_ ), .X(\us10\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1006_ ( .A1(\us10\/_0193_ ), .A2(\us10\/_0176_ ), .B1(\us10\/_0043_ ), .Y(\us10\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1007_ ( .A(\us10\/_0185_ ), .B(\us10\/_0189_ ), .C(\us10\/_0192_ ), .D(\us10\/_0195_ ), .X(\us10\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us10/_1008_ ( .A_N(\sa10\[3\] ), .B(\us10\/_0734_ ), .C(\sa10\[2\] ), .X(\us10\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1009_ ( .A(\us10\/_0137_ ), .B(\us10\/_0197_ ), .X(\us10\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_1010_ ( .A(\us10\/_0198_ ), .B(\us10\/_0040_ ), .Y(\us10\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1011_ ( .A(\us10\/_0293_ ), .B(\us10\/_0137_ ), .X(\us10\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1012_ ( .A(\us10\/_0200_ ), .Y(\us10\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1013_ ( .A(\us10\/_0137_ ), .B(\us10\/_0110_ ), .Y(\us10\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1014_ ( .A(\us10\/_0139_ ), .B(\us10\/_0020_ ), .Y(\us10\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1015_ ( .A(\us10\/_0199_ ), .B(\us10\/_0201_ ), .C(\us10\/_0202_ ), .D(\us10\/_0203_ ), .X(\us10\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us10/_1016_ ( .A1(\us10\/_0532_ ), .A2(\us10\/_0109_ ), .B1(\us10\/_0102_ ), .C1(\us10\/_0727_ ), .X(\us10\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1017_ ( .A(\us10\/_0023_ ), .B(\us10\/_0078_ ), .Y(\us10\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1018_ ( .A(\us10\/_0078_ ), .B(\us10\/_0142_ ), .Y(\us10\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1019_ ( .A(\us10\/_0207_ ), .B(\us10\/_0208_ ), .Y(\us10\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1020_ ( .A1(\us10\/_0094_ ), .A2(\us10\/_0176_ ), .B1(\us10\/_0206_ ), .C1(\us10\/_0209_ ), .Y(\us10\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1021_ ( .A(\us10\/_0662_ ), .B(\us10\/_0070_ ), .X(\us10\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us10/_1022_ ( .A(\us10\/_0732_ ), .B(\us10\/_0123_ ), .C(\us10\/_0749_ ), .Y(\us10\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us10/_1023_ ( .A(\us10\/_0732_ ), .B(\us10\/_0467_ ), .C(\us10\/_0069_ ), .Y(\us10\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us10/_1024_ ( .A_N(\us10\/_0211_ ), .B(\us10\/_0127_ ), .C(\us10\/_0212_ ), .D(\us10\/_0213_ ), .X(\us10\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1025_ ( .A(\us10\/_0137_ ), .Y(\us10\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1026_ ( .A(\us10\/_0128_ ), .B(\us10\/_0036_ ), .Y(\us10\/_0217_ ) );
sky130_fd_sc_hd__buf_2 \us10/_1027_ ( .A(\us10\/_0489_ ), .X(\us10\/_0218_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1028_ ( .A1(\us10\/_0159_ ), .A2(\us10\/_0746_ ), .B1(\us10\/_0445_ ), .B2(\us10\/_0218_ ), .Y(\us10\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us10/_1029_ ( .A1(\us10\/_0116_ ), .A2(\us10\/_0215_ ), .B1(\us10\/_0217_ ), .C1(\us10\/_0219_ ), .X(\us10\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1030_ ( .A(\us10\/_0113_ ), .B(\us10\/_0746_ ), .X(\us10\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us10/_1031_ ( .A1(\us10\/_0098_ ), .A2(\us10\/_0746_ ), .B1(\us10\/_0445_ ), .B2(\us10\/_0750_ ), .X(\us10\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1032_ ( .A1(\us10\/_0048_ ), .A2(\us10\/_0113_ ), .B1(\us10\/_0221_ ), .C1(\us10\/_0222_ ), .Y(\us10\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us10/_1033_ ( .A1(\us10\/_0129_ ), .A2(\us10\/_0162_ ), .B1(\us10\/_0282_ ), .B2(\us10\/_0705_ ), .X(\us10\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1034_ ( .A1(\us10\/_0093_ ), .A2(\us10\/_0738_ ), .B1(\us10\/_0081_ ), .C1(\us10\/_0224_ ), .Y(\us10\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1035_ ( .A(\us10\/_0214_ ), .B(\us10\/_0220_ ), .C(\us10\/_0223_ ), .D(\us10\/_0225_ ), .X(\us10\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1036_ ( .A(\us10\/_0196_ ), .B(\us10\/_0204_ ), .C(\us10\/_0210_ ), .D(\us10\/_0226_ ), .X(\us10\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1037_ ( .A(\us10\/_0111_ ), .B(\us10\/_0554_ ), .X(\us10\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1038_ ( .A(\us10\/_0229_ ), .Y(\us10\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1039_ ( .A(\us10\/_0111_ ), .B(\us10\/_0129_ ), .Y(\us10\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1040_ ( .A(\us10\/_0018_ ), .B(\us10\/_0738_ ), .Y(\us10\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1041_ ( .A(\us10\/_0030_ ), .B(\us10\/_0304_ ), .Y(\us10\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1042_ ( .A(\us10\/_0230_ ), .B(\us10\/_0231_ ), .C(\us10\/_0232_ ), .D(\us10\/_0233_ ), .X(\us10\/_0234_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1043_ ( .A(\us10\/_0048_ ), .B(\us10\/_0489_ ), .X(\us10\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1044_ ( .A1(\us10\/_0129_ ), .A2(\us10\/_0554_ ), .B1(\us10\/_0137_ ), .Y(\us10\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us10/_1045_ ( .A(\us10\/_0235_ ), .B(\us10\/_0049_ ), .C_N(\us10\/_0236_ ), .Y(\us10\/_0237_ ) );
sky130_fd_sc_hd__and2_1 \us10/_1046_ ( .A(\us10\/_0047_ ), .B(\us10\/_0077_ ), .X(\us10\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1047_ ( .A(\us10\/_0070_ ), .B(\us10\/_0036_ ), .X(\us10\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us10/_1048_ ( .A1(\us10\/_0048_ ), .A2(\us10\/_0736_ ), .B1(\us10\/_0023_ ), .B2(\us10\/_0099_ ), .X(\us10\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us10/_1049_ ( .A(\us10\/_0239_ ), .B(\us10\/_0240_ ), .C(\us10\/_0241_ ), .Y(\us10\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1050_ ( .A(\us10\/_0554_ ), .B(\us10\/_0072_ ), .X(\us10\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us10/_1051_ ( .A1(\us10\/_0142_ ), .A2(\us10\/_0137_ ), .B1(\us10\/_0159_ ), .B2(\us10\/_0083_ ), .X(\us10\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1052_ ( .A1(\us10\/_0608_ ), .A2(\us10\/_0072_ ), .B1(\us10\/_0243_ ), .C1(\us10\/_0244_ ), .Y(\us10\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1053_ ( .A(\us10\/_0234_ ), .B(\us10\/_0237_ ), .C(\us10\/_0242_ ), .D(\us10\/_0245_ ), .X(\us10\/_0246_ ) );
sky130_fd_sc_hd__o21a_1 \us10/_1055_ ( .A1(\us10\/_0554_ ), .A2(\us10\/_0586_ ), .B1(\us10\/_0029_ ), .X(\us10\/_0248_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1056_ ( .A(\us10\/_0083_ ), .B(\us10\/_0489_ ), .X(\us10\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_1057_ ( .A(\us10\/_0079_ ), .X(\us10\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1058_ ( .A(\us10\/_0251_ ), .B(\us10\/_0489_ ), .X(\us10\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_1059_ ( .A(\us10\/_0250_ ), .B(\us10\/_0252_ ), .Y(\us10\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1060_ ( .A(\us10\/_0016_ ), .B(\us10\/_0064_ ), .Y(\us10\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_1061_ ( .A(\us10\/_0304_ ), .X(\us10\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1062_ ( .A(\us10\/_0255_ ), .B(\us10\/_0640_ ), .Y(\us10\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us10/_1063_ ( .A_N(\us10\/_0248_ ), .B(\us10\/_0253_ ), .C(\us10\/_0254_ ), .D(\us10\/_0256_ ), .X(\us10\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1064_ ( .A(\us10\/_0099_ ), .B(\us10\/_0110_ ), .X(\us10\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us10/_1065_ ( .A1(\us10\/_0161_ ), .A2(\us10\/_0130_ ), .B1(\us10\/_0258_ ), .Y(\us10\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1066_ ( .A(\us10\/_0194_ ), .B(\sa10\[1\] ), .X(\us10\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1068_ ( .A(\us10\/_0261_ ), .B(\us10\/_0153_ ), .Y(\us10\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us10/_1069_ ( .A_N(\us10\/_0154_ ), .B(\us10\/_0259_ ), .C(\us10\/_0263_ ), .X(\us10\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1070_ ( .A(\us10\/_0246_ ), .B(\us10\/_0174_ ), .C(\us10\/_0257_ ), .D(\us10\/_0264_ ), .X(\us10\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us10/_1071_ ( .A1(\us10\/_0261_ ), .A2(\us10\/_0554_ ), .B1(\us10\/_0159_ ), .X(\us10\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1072_ ( .A(\us10\/_0746_ ), .B(\us10\/_0150_ ), .Y(\us10\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1073_ ( .A(\us10\/_0175_ ), .Y(\us10\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us10/_1074_ ( .A(\us10\/_0423_ ), .B(\us10\/_0123_ ), .C(\us10\/_0151_ ), .X(\us10\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1075_ ( .A(\us10\/_0268_ ), .B(\us10\/_0269_ ), .Y(\us10\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us10/_1076_ ( .A_N(\us10\/_0266_ ), .B(\us10\/_0267_ ), .C(\us10\/_0270_ ), .X(\us10\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1077_ ( .A(\us10\/_0554_ ), .B(\us10\/_0150_ ), .X(\us10\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1078_ ( .A(\us10\/_0273_ ), .Y(\us10\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1079_ ( .A1(\us10\/_0734_ ), .A2(\us10\/_0325_ ), .B1(\us10\/_0380_ ), .Y(\us10\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1080_ ( .A(\us10\/_0275_ ), .Y(\us10\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1081_ ( .A(\us10\/_0276_ ), .B(\us10\/_0153_ ), .Y(\us10\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us10/_1082_ ( .A(\us10\/_0272_ ), .B(\us10\/_0274_ ), .C(\us10\/_0277_ ), .X(\us10\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_1083_ ( .A(\us10\/_0036_ ), .X(\us10\/_0279_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1085_ ( .A1(\us10\/_0218_ ), .A2(\us10\/_0279_ ), .B1(\us10\/_0084_ ), .B2(\us10\/_0060_ ), .Y(\us10\/_0281_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1086_ ( .A1(\us10\/_0251_ ), .A2(\us10\/_0445_ ), .B1(\us10\/_0304_ ), .Y(\us10\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1087_ ( .A(\us10\/_0091_ ), .B(\us10\/_0056_ ), .Y(\us10\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1088_ ( .A1(\us10\/_0118_ ), .A2(\us10\/_0050_ ), .B1(\us10\/_0038_ ), .C1(\us10\/_0255_ ), .Y(\us10\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1089_ ( .A(\us10\/_0281_ ), .B(\us10\/_0283_ ), .C(\us10\/_0284_ ), .D(\us10\/_0285_ ), .X(\us10\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1090_ ( .A(\us10\/_0083_ ), .B(\us10\/_0027_ ), .X(\us10\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1091_ ( .A(\us10\/_0129_ ), .B(\us10\/_0027_ ), .X(\us10\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_1092_ ( .A(\us10\/_0287_ ), .B(\us10\/_0288_ ), .Y(\us10\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1093_ ( .A1(\us10\/_0752_ ), .A2(\us10\/_0683_ ), .B1(\us10\/_0093_ ), .B2(\us10\/_0029_ ), .Y(\us10\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1094_ ( .A1(\us10\/_0092_ ), .A2(\us10\/_0575_ ), .B1(\us10\/_0056_ ), .Y(\us10\/_0291_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1096_ ( .A1(\us10\/_0218_ ), .A2(\us10\/_0672_ ), .B1(\us10\/_0084_ ), .B2(\us10\/_0056_ ), .Y(\us10\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1097_ ( .A(\us10\/_0289_ ), .B(\us10\/_0290_ ), .C(\us10\/_0291_ ), .D(\us10\/_0294_ ), .X(\us10\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1098_ ( .A(\us10\/_0750_ ), .B(\us10\/_0193_ ), .X(\us10\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1099_ ( .A(\us10\/_0705_ ), .B(\us10\/_0380_ ), .X(\us10\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1100_ ( .A(\us10\/_0752_ ), .B(\us10\/_0129_ ), .Y(\us10\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us10/_1101_ ( .A(\us10\/_0296_ ), .B(\us10\/_0297_ ), .C_N(\us10\/_0298_ ), .Y(\us10\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1102_ ( .A(\us10\/_0089_ ), .B(\us10\/_0532_ ), .Y(\us10\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1103_ ( .A(\sa10\[2\] ), .Y(\us10\/_0301_ ) );
sky130_fd_sc_hd__nor3_2 \us10/_1104_ ( .A(\us10\/_0301_ ), .B(\sa10\[3\] ), .C(\us10\/_0118_ ), .Y(\us10\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1105_ ( .A(\us10\/_0072_ ), .B(\us10\/_0302_ ), .X(\us10\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1106_ ( .A(\us10\/_0303_ ), .Y(\us10\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1107_ ( .A(\us10\/_0147_ ), .B(\us10\/_0302_ ), .Y(\us10\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1108_ ( .A(\us10\/_0299_ ), .B(\us10\/_0300_ ), .C(\us10\/_0305_ ), .D(\us10\/_0306_ ), .X(\us10\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1109_ ( .A(\us10\/_0278_ ), .B(\us10\/_0286_ ), .C(\us10\/_0295_ ), .D(\us10\/_0307_ ), .X(\us10\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us10/_1110_ ( .A(\us10\/_0228_ ), .B(\us10\/_0265_ ), .C(\us10\/_0308_ ), .Y(\us10\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1111_ ( .A(\us10\/_0235_ ), .Y(\us10\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1112_ ( .A(\us10\/_0489_ ), .B(\us10\/_0640_ ), .X(\us10\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1113_ ( .A(\us10\/_0310_ ), .Y(\us10\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1114_ ( .A(\us10\/_0023_ ), .B(\us10\/_0218_ ), .Y(\us10\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1115_ ( .A(\us10\/_0218_ ), .B(\us10\/_0032_ ), .Y(\us10\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1116_ ( .A(\us10\/_0309_ ), .B(\us10\/_0311_ ), .C(\us10\/_0312_ ), .D(\us10\/_0313_ ), .X(\us10\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1117_ ( .A(\us10\/_0218_ ), .B(\us10\/_0064_ ), .Y(\us10\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1118_ ( .A(\us10\/_0218_ ), .B(\us10\/_0683_ ), .Y(\us10\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1119_ ( .A(\us10\/_0315_ ), .B(\us10\/_0316_ ), .C(\us10\/_0317_ ), .D(\us10\/_0253_ ), .X(\us10\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1120_ ( .A(\us10\/_0048_ ), .B(\us10\/_0304_ ), .Y(\us10\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1121_ ( .A(\us10\/_0586_ ), .B(\us10\/_0162_ ), .Y(\us10\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1122_ ( .A(\us10\/_0319_ ), .B(\us10\/_0320_ ), .Y(\us10\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_1123_ ( .A(\us10\/_0321_ ), .B(\us10\/_0238_ ), .Y(\us10\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1124_ ( .A(\us10\/_0304_ ), .B(\us10\/_0062_ ), .Y(\us10\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_1125_ ( .A(\us10\/_0251_ ), .X(\us10\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1126_ ( .A1(\us10\/_0324_ ), .A2(\us10\/_0084_ ), .B1(\us10\/_0255_ ), .Y(\us10\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1127_ ( .A1(\us10\/_0050_ ), .A2(\us10\/_0216_ ), .B1(\us10\/_0109_ ), .C1(\us10\/_0255_ ), .Y(\us10\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1128_ ( .A(\us10\/_0322_ ), .B(\us10\/_0323_ ), .C(\us10\/_0326_ ), .D(\us10\/_0327_ ), .X(\us10\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1129_ ( .A1(\us10\/_0733_ ), .A2(\us10\/_0279_ ), .A3(\us10\/_0058_ ), .B1(\us10\/_0056_ ), .Y(\us10\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_1130_ ( .A(\us10\/_0048_ ), .X(\us10\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1131_ ( .A(\us10\/_0330_ ), .B(\us10\/_0056_ ), .Y(\us10\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1132_ ( .A(\us10\/_0055_ ), .B(\us10\/_0045_ ), .Y(\us10\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1133_ ( .A(\us10\/_0329_ ), .B(\us10\/_0331_ ), .C(\us10\/_0284_ ), .D(\us10\/_0332_ ), .X(\us10\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us10/_1134_ ( .A1(\us10\/_0543_ ), .A2(\us10\/_0216_ ), .B1(\us10\/_0532_ ), .C1(\us10\/_0060_ ), .X(\us10\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1135_ ( .A(\us10\/_0084_ ), .B(\us10\/_0060_ ), .Y(\us10\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1136_ ( .A(\us10\/_0324_ ), .B(\us10\/_0060_ ), .Y(\us10\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1137_ ( .A(\us10\/_0335_ ), .B(\us10\/_0337_ ), .Y(\us10\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1138_ ( .A1(\us10\/_0276_ ), .A2(\us10\/_0060_ ), .B1(\us10\/_0334_ ), .C1(\us10\/_0338_ ), .Y(\us10\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1139_ ( .A(\us10\/_0318_ ), .B(\us10\/_0328_ ), .C(\us10\/_0333_ ), .D(\us10\/_0339_ ), .X(\us10\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us10/_1140_ ( .A1(\us10\/_0746_ ), .A2(\us10\/_0134_ ), .B1(\us10\/_0128_ ), .X(\us10\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us10/_1141_ ( .A_N(\us10\/_0086_ ), .B(\us10\/_0128_ ), .X(\us10\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1142_ ( .A(\us10\/_0079_ ), .B(\us10\/_0124_ ), .X(\us10\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_1143_ ( .A(\us10\/_0126_ ), .B(\us10\/_0343_ ), .Y(\us10\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us10/_1144_ ( .A(\us10\/_0341_ ), .B(\us10\/_0342_ ), .C_N(\us10\/_0344_ ), .Y(\us10\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1146_ ( .A1(\us10\/_0193_ ), .A2(\us10\/_0092_ ), .A3(\us10\/_0330_ ), .B1(\us10\/_0147_ ), .Y(\us10\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1147_ ( .A1(\us10\/_0130_ ), .A2(\us10\/_0084_ ), .A3(\us10\/_0134_ ), .B1(\us10\/_0139_ ), .Y(\us10\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1148_ ( .A1(\us10\/_0144_ ), .A2(\us10\/_0608_ ), .A3(\us10\/_0092_ ), .B1(\us10\/_0139_ ), .Y(\us10\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1149_ ( .A(\us10\/_0345_ ), .B(\us10\/_0348_ ), .C(\us10\/_0349_ ), .D(\us10\/_0350_ ), .X(\us10\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us10/_1150_ ( .A(\us10\/_0150_ ), .B(\us10\/_0194_ ), .C(\us10\/_0543_ ), .X(\us10\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us10/_1151_ ( .A(\us10\/_0277_ ), .SLEEP(\us10\/_0352_ ), .X(\us10\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us10/_1152_ ( .A1(\us10\/_0268_ ), .A2(\us10\/_0171_ ), .B1(\us10\/_0157_ ), .Y(\us10\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us10/_1153_ ( .A(\us10\/_0161_ ), .X(\us10\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1154_ ( .A1(\us10\/_0279_ ), .A2(\us10\/_0084_ ), .B1(\us10\/_0355_ ), .Y(\us10\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1155_ ( .A1(\us10\/_0020_ ), .A2(\us10\/_0193_ ), .A3(\us10\/_0091_ ), .B1(\us10\/_0355_ ), .Y(\us10\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1156_ ( .A(\us10\/_0353_ ), .B(\us10\/_0354_ ), .C(\us10\/_0356_ ), .D(\us10\/_0357_ ), .X(\us10\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1157_ ( .A(\us10\/_0111_ ), .B(\us10\/_0586_ ), .X(\us10\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1158_ ( .A(\us10\/_0360_ ), .Y(\us10\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us10/_1159_ ( .A1(\us10\/_0119_ ), .A2(\us10\/_0120_ ), .B1(\us10\/_0230_ ), .C1(\us10\/_0361_ ), .X(\us10\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1160_ ( .A1(\us10\/_0672_ ), .A2(\us10\/_0251_ ), .A3(\us10\/_0134_ ), .B1(\us10\/_0114_ ), .Y(\us10\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1162_ ( .A1(\us10\/_0036_ ), .A2(\us10\/_0251_ ), .A3(\us10\/_0134_ ), .B1(\us10\/_0099_ ), .Y(\us10\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1163_ ( .A1(\us10\/_0193_ ), .A2(\us10\/_0608_ ), .B1(\us10\/_0099_ ), .Y(\us10\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1164_ ( .A(\us10\/_0362_ ), .B(\us10\/_0363_ ), .C(\us10\/_0365_ ), .D(\us10\/_0366_ ), .X(\us10\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1165_ ( .A1(\us10\/_0575_ ), .A2(\us10\/_0092_ ), .A3(\us10\/_0330_ ), .B1(\us10\/_0089_ ), .Y(\us10\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1166_ ( .A1(\us10\/_0586_ ), .A2(\us10\/_0018_ ), .A3(\us10\/_0330_ ), .B1(\us10\/_0094_ ), .Y(\us10\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \us10/_1167_ ( .A1(\us10\/_0293_ ), .A2(\us10\/_0134_ ), .B1(\us10\/_0089_ ), .Y(\us10\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1168_ ( .A1(\us10\/_0279_ ), .A2(\us10\/_0134_ ), .B1(\us10\/_0094_ ), .Y(\us10\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1169_ ( .A(\us10\/_0368_ ), .B(\us10\/_0370_ ), .C(\us10\/_0371_ ), .D(\us10\/_0372_ ), .X(\us10\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1170_ ( .A(\us10\/_0351_ ), .B(\us10\/_0359_ ), .C(\us10\/_0367_ ), .D(\us10\/_0373_ ), .X(\us10\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1171_ ( .A1(\us10\/_0102_ ), .A2(\us10\/_0347_ ), .B1(\us10\/_0109_ ), .C1(\us10\/_0029_ ), .Y(\us10\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1172_ ( .A1(\us10\/_0102_ ), .A2(\us10\/_0347_ ), .B1(\us10\/_0532_ ), .C1(\us10\/_0029_ ), .Y(\us10\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1173_ ( .A1(\us10\/_0050_ ), .A2(\us10\/_0543_ ), .B1(\us10\/_0380_ ), .C1(\us10\/_0029_ ), .Y(\us10\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1174_ ( .A(\us10\/_0041_ ), .B(\us10\/_0375_ ), .C(\us10\/_0376_ ), .D(\us10\/_0377_ ), .X(\us10\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1175_ ( .A(\us10\/_0048_ ), .B(\us10\/_0750_ ), .X(\us10\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1176_ ( .A(\us10\/_0379_ ), .Y(\us10\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1177_ ( .A(\us10\/_0016_ ), .B(\us10\/_0608_ ), .Y(\us10\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1178_ ( .A(\us10\/_0752_ ), .B(\us10\/_0554_ ), .Y(\us10\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1179_ ( .A1(\sa10\[1\] ), .A2(\us10\/_0734_ ), .B1(\us10\/_0109_ ), .C1(\us10\/_0016_ ), .Y(\us10\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1180_ ( .A(\us10\/_0381_ ), .B(\us10\/_0382_ ), .C(\us10\/_0383_ ), .D(\us10\/_0384_ ), .X(\us10\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us10/_1181_ ( .A(\us10\/_0086_ ), .B_N(\us10\/_0736_ ), .X(\us10\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1182_ ( .A1(\us10\/_0748_ ), .A2(\us10\/_0134_ ), .B1(\us10\/_0739_ ), .Y(\us10\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1183_ ( .A1(\us10\/_0118_ ), .A2(\us10\/_0543_ ), .B1(\us10\/_0109_ ), .C1(\us10\/_0739_ ), .Y(\us10\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1184_ ( .A1(\us10\/_0102_ ), .A2(\us10\/_0301_ ), .B1(\sa10\[3\] ), .C1(\us10\/_0739_ ), .Y(\us10\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1185_ ( .A(\us10\/_0386_ ), .B(\us10\/_0387_ ), .C(\us10\/_0388_ ), .D(\us10\/_0389_ ), .X(\us10\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1186_ ( .A(\us10\/_0020_ ), .Y(\us10\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1187_ ( .A(\us10\/_0727_ ), .Y(\us10\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1188_ ( .A(\us10\/_0727_ ), .B(\us10\/_0064_ ), .Y(\us10\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1189_ ( .A1(\us10\/_0102_ ), .A2(\us10\/_0734_ ), .B1(\us10\/_0532_ ), .C1(\us10\/_0727_ ), .Y(\us10\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us10/_1190_ ( .A1(\us10\/_0392_ ), .A2(\us10\/_0393_ ), .B1(\us10\/_0394_ ), .C1(\us10\/_0395_ ), .X(\us10\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1191_ ( .A(\us10\/_0378_ ), .B(\us10\/_0385_ ), .C(\us10\/_0390_ ), .D(\us10\/_0396_ ), .X(\us10\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us10/_1192_ ( .A(\us10\/_0340_ ), .B(\us10\/_0374_ ), .C(\us10\/_0397_ ), .Y(\us10\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1193_ ( .A(\us10\/_0077_ ), .B(\us10\/_0129_ ), .X(\us10\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_1194_ ( .A(\us10\/_0398_ ), .B(\us10\/_0239_ ), .Y(\us10\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1195_ ( .A(\us10\/_0023_ ), .B(\us10\/_0111_ ), .X(\us10\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us10/_1196_ ( .A_N(\us10\/_0400_ ), .B(\us10\/_0231_ ), .Y(\us10\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us10/_1197_ ( .A(\us10\/_0399_ ), .SLEEP(\us10\/_0402_ ), .X(\us10\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_1198_ ( .A(\us10\/_0746_ ), .B(\us10\/_0251_ ), .Y(\us10\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us10/_1199_ ( .A_N(\us10\/_0404_ ), .B(\us10\/_0752_ ), .Y(\us10\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us10/_1200_ ( .A(\us10\/_0467_ ), .B(\us10\/_0194_ ), .C(\us10\/_0694_ ), .X(\us10\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us10/_1201_ ( .A_N(\us10\/_0175_ ), .B(\us10\/_0406_ ), .X(\us10\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1202_ ( .A(\us10\/_0407_ ), .Y(\us10\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1203_ ( .A1(\us10\/_0094_ ), .A2(\us10\/_0197_ ), .B1(\us10\/_0114_ ), .B2(\us10\/_0640_ ), .Y(\us10\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1204_ ( .A(\us10\/_0403_ ), .B(\us10\/_0405_ ), .C(\us10\/_0408_ ), .D(\us10\/_0409_ ), .X(\us10\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1205_ ( .A(\us10\/_0030_ ), .B(\us10\/_0150_ ), .Y(\us10\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us10/_1206_ ( .A_N(\us10\/_0169_ ), .B(\us10\/_0289_ ), .C(\us10\/_0411_ ), .X(\us10\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us10/_1207_ ( .A1(\us10\/_0467_ ), .A2(\us10\/_0151_ ), .B1(\us10\/_0140_ ), .C1(\us10\/_0129_ ), .X(\us10\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1208_ ( .A1(\us10\/_0608_ ), .A2(\us10\/_0099_ ), .B1(\us10\/_0037_ ), .C1(\us10\/_0414_ ), .Y(\us10\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1209_ ( .A(\us10\/_0738_ ), .Y(\us10\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1210_ ( .A(\us10\/_0586_ ), .B(\us10\/_0736_ ), .Y(\us10\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1211_ ( .A1(\us10\/_0194_ ), .A2(\us10\/_0038_ ), .B1(\us10\/_0118_ ), .C1(\us10\/_0153_ ), .Y(\us10\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us10/_1212_ ( .A1(\us10\/_0416_ ), .A2(\us10\/_0117_ ), .B1(\us10\/_0417_ ), .C1(\us10\/_0418_ ), .X(\us10\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1213_ ( .A(\us10\/_0077_ ), .B(\us10\/_0035_ ), .X(\us10\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1214_ ( .A(\us10\/_0672_ ), .B(\us10\/_0124_ ), .Y(\us10\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1215_ ( .A(\us10\/_0030_ ), .B(\us10\/_0137_ ), .Y(\us10\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1216_ ( .A(\us10\/_0072_ ), .B(\us10\/_0732_ ), .Y(\us10\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us10/_1217_ ( .A_N(\us10\/_0420_ ), .B(\us10\/_0421_ ), .C(\us10\/_0422_ ), .D(\us10\/_0424_ ), .X(\us10\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1218_ ( .A(\us10\/_0413_ ), .B(\us10\/_0415_ ), .C(\us10\/_0419_ ), .D(\us10\/_0425_ ), .X(\us10\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us10/_1219_ ( .A(\us10\/_0355_ ), .B(\us10\/_0102_ ), .C(\us10\/_0109_ ), .Y(\us10\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1220_ ( .A(\us10\/_0077_ ), .B(\us10\/_0018_ ), .X(\us10\/_0428_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1221_ ( .A(\us10\/_0077_ ), .B(\us10\/_0554_ ), .X(\us10\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us10/_1222_ ( .A1(\us10\/_0050_ ), .A2(\us10\/_0216_ ), .B1(\us10\/_0380_ ), .C1(\us10\/_0078_ ), .X(\us10\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us10/_1223_ ( .A(\us10\/_0428_ ), .B(\us10\/_0429_ ), .C(\us10\/_0430_ ), .Y(\us10\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us10/_1224_ ( .A_N(\us10\/_0209_ ), .B(\us10\/_0431_ ), .X(\us10\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us10/_1225_ ( .A1(\us10\/_0215_ ), .A2(\us10\/_0404_ ), .B1(\us10\/_0427_ ), .C1(\us10\/_0432_ ), .X(\us10\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1226_ ( .A(\us10\/_0043_ ), .B(\us10\/_0058_ ), .Y(\us10\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1227_ ( .A(\us10\/_0195_ ), .B(\us10\/_0233_ ), .C(\us10\/_0320_ ), .D(\us10\/_0435_ ), .X(\us10\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1228_ ( .A(\us10\/_0261_ ), .B(\us10\/_0738_ ), .Y(\us10\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1229_ ( .A1(\us10\/_0218_ ), .A2(\us10\/_0640_ ), .B1(\us10\/_0261_ ), .B2(\us10\/_0056_ ), .Y(\us10\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1230_ ( .A(\us10\/_0436_ ), .B(\us10\/_0394_ ), .C(\us10\/_0437_ ), .D(\us10\/_0438_ ), .X(\us10\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1231_ ( .A(\us10\/_0410_ ), .B(\us10\/_0426_ ), .C(\us10\/_0433_ ), .D(\us10\/_0439_ ), .X(\us10\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us10/_1232_ ( .A(\us10\/_0135_ ), .SLEEP(\us10\/_0273_ ), .X(\us10\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1233_ ( .A1(\us10\/_0279_ ), .A2(\us10\/_0134_ ), .B1(\us10\/_0099_ ), .Y(\us10\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1234_ ( .A(\us10\/_0441_ ), .B(\us10\/_0164_ ), .C(\us10\/_0270_ ), .D(\us10\/_0442_ ), .X(\us10\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1235_ ( .A(\us10\/_0051_ ), .B(\us10\/_0672_ ), .Y(\us10\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1236_ ( .A(\us10\/_0051_ ), .B(\us10\/_0282_ ), .Y(\us10\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1237_ ( .A(\us10\/_0444_ ), .B(\us10\/_0446_ ), .X(\us10\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1238_ ( .A(\us10\/_0193_ ), .B(\us10\/_0304_ ), .X(\us10\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1239_ ( .A(\us10\/_0448_ ), .Y(\us10\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1240_ ( .A(\us10\/_0162_ ), .B(\us10\/_0130_ ), .X(\us10\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1241_ ( .A(\us10\/_0450_ ), .Y(\us10\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1242_ ( .A1(\us10\/_0129_ ), .A2(\us10\/_0554_ ), .B1(\us10\/_0043_ ), .Y(\us10\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1243_ ( .A(\us10\/_0447_ ), .B(\us10\/_0449_ ), .C(\us10\/_0451_ ), .D(\us10\/_0452_ ), .X(\us10\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1244_ ( .A(\us10\/_0056_ ), .B(\us10\/_0064_ ), .Y(\us10\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us10/_1245_ ( .A_N(\us10\/_0248_ ), .B(\us10\/_0454_ ), .C(\us10\/_0254_ ), .D(\us10\/_0256_ ), .X(\us10\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1246_ ( .A1(\us10\/_0330_ ), .A2(\us10\/_0099_ ), .B1(\us10\/_0134_ ), .B2(\us10\/_0705_ ), .Y(\us10\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1247_ ( .A1(\us10\/_0748_ ), .A2(\us10\/_0738_ ), .B1(\us10\/_0092_ ), .B2(\us10\/_0752_ ), .Y(\us10\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1248_ ( .A1(\us10\/_0072_ ), .A2(\us10\/_0036_ ), .B1(\us10\/_0748_ ), .B2(\us10\/_0056_ ), .Y(\us10\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1249_ ( .A1(\us10\/_0748_ ), .A2(\us10\/_0251_ ), .B1(\us10\/_0029_ ), .Y(\us10\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1250_ ( .A(\us10\/_0457_ ), .B(\us10\/_0458_ ), .C(\us10\/_0459_ ), .D(\us10\/_0460_ ), .X(\us10\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1251_ ( .A(\us10\/_0443_ ), .B(\us10\/_0453_ ), .C(\us10\/_0455_ ), .D(\us10\/_0461_ ), .X(\us10\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1252_ ( .A(\us10\/_0705_ ), .B(\us10\/_0079_ ), .X(\us10\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1253_ ( .A(\us10\/_0586_ ), .B(\us10\/_0124_ ), .Y(\us10\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1254_ ( .A(\us10\/_0218_ ), .B(\us10\/_0746_ ), .Y(\us10\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us10/_1255_ ( .A_N(\us10\/_0463_ ), .B(\us10\/_0464_ ), .C(\us10\/_0465_ ), .X(\us10\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us10/_1256_ ( .A1(\us10\/_0282_ ), .A2(\us10\/_0072_ ), .B1(\us10\/_0142_ ), .B2(\us10\/_0027_ ), .X(\us10\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1257_ ( .A1(\us10\/_0144_ ), .A2(\us10\/_0099_ ), .B1(\us10\/_0360_ ), .C1(\us10\/_0468_ ), .Y(\us10\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us10/_1258_ ( .A1(\us10\/_0672_ ), .A2(\us10\/_0251_ ), .B1(\us10\/_0218_ ), .X(\us10\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1259_ ( .A1(\us10\/_0575_ ), .A2(\us10\/_0056_ ), .B1(\us10\/_0379_ ), .C1(\us10\/_0470_ ), .Y(\us10\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1260_ ( .A(\us10\/_0466_ ), .B(\us10\/_0469_ ), .C(\us10\/_0471_ ), .D(\us10\/_0305_ ), .X(\us10\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us10/_1261_ ( .A1(\us10\/_0029_ ), .A2(\us10\/_0683_ ), .B1(\us10\/_0324_ ), .B2(\us10\/_0056_ ), .X(\us10\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1262_ ( .A(\us10\/_0084_ ), .B(\us10\/_0099_ ), .X(\us10\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us10/_1263_ ( .A1(\us10\/_0092_ ), .A2(\us10\/_0029_ ), .B1(\us10\/_0474_ ), .X(\us10\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us10/_1264_ ( .A(\us10\/_0075_ ), .B(\us10\/_0473_ ), .C(\us10\/_0475_ ), .Y(\us10\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1265_ ( .A1(\us10\/_0279_ ), .A2(\us10\/_0255_ ), .B1(\us10\/_0084_ ), .B2(\us10\/_0060_ ), .Y(\us10\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1266_ ( .A1(\us10\/_0093_ ), .A2(\us10\/_0056_ ), .B1(\us10\/_0134_ ), .B2(\us10\/_0114_ ), .Y(\us10\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1267_ ( .A1(\us10\/_0161_ ), .A2(\us10\/_0032_ ), .B1(\us10\/_0324_ ), .B2(\us10\/_0147_ ), .Y(\us10\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1268_ ( .A1(\us10\/_0055_ ), .A2(\us10\/_0732_ ), .B1(\us10\/_0748_ ), .B2(\us10\/_0304_ ), .Y(\us10\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1269_ ( .A(\us10\/_0477_ ), .B(\us10\/_0479_ ), .C(\us10\/_0480_ ), .D(\us10\/_0481_ ), .X(\us10\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1270_ ( .A(\us10\/_0161_ ), .B(\us10\/_0064_ ), .Y(\us10\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us10/_1271_ ( .A(\us10\/_0732_ ), .B(\us10\/_0123_ ), .C(\us10\/_0467_ ), .Y(\us10\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1272_ ( .A(\us10\/_0483_ ), .B(\us10\/_0484_ ), .Y(\us10\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1273_ ( .A(\us10\/_0297_ ), .Y(\us10\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us10/_1274_ ( .A_N(\us10\/_0485_ ), .B(\us10\/_0181_ ), .C(\us10\/_0486_ ), .D(\us10\/_0386_ ), .X(\us10\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1275_ ( .A(\us10\/_0472_ ), .B(\us10\/_0476_ ), .C(\us10\/_0482_ ), .D(\us10\/_0487_ ), .X(\us10\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \us10/_1276_ ( .A(\us10\/_0440_ ), .B(\us10\/_0462_ ), .C(\us10\/_0488_ ), .Y(\us10\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1277_ ( .A(\us10\/_0403_ ), .B(\us10\/_0230_ ), .C(\us10\/_0451_ ), .D(\us10\/_0361_ ), .X(\us10\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1278_ ( .A1(\us10\/_0118_ ), .A2(\us10\/_0050_ ), .B1(\us10\/_0109_ ), .C1(\us10\/_0139_ ), .Y(\us10\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1279_ ( .A(\us10\/_0447_ ), .B(\us10\/_0437_ ), .C(\us10\/_0491_ ), .D(\us10\/_0427_ ), .X(\us10\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1280_ ( .A1(\us10\/_0084_ ), .A2(\us10\/_0255_ ), .B1(\us10\/_0608_ ), .B2(\us10\/_0029_ ), .Y(\us10\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1281_ ( .A1(\us10\/_0144_ ), .A2(\us10\/_0147_ ), .B1(\us10\/_0355_ ), .B2(\us10\/_0093_ ), .Y(\us10\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1282_ ( .A1(\us10\/_0705_ ), .A2(\us10\/_0279_ ), .B1(\us10\/_0330_ ), .B2(\us10\/_0029_ ), .Y(\us10\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1283_ ( .A1(\us10\/_0279_ ), .A2(\us10\/_0084_ ), .B1(\us10\/_0114_ ), .Y(\us10\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1284_ ( .A(\us10\/_0493_ ), .B(\us10\/_0494_ ), .C(\us10\/_0495_ ), .D(\us10\/_0496_ ), .X(\us10\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1285_ ( .A1(\us10\/_0134_ ), .A2(\us10\/_0137_ ), .B1(\us10\/_0355_ ), .B2(\us10\/_0575_ ), .Y(\us10\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1286_ ( .A1(\us10\/_0099_ ), .A2(\us10\/_0733_ ), .B1(\us10\/_0093_ ), .B2(\us10\/_0218_ ), .Y(\us10\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1287_ ( .A(\us10\/_0147_ ), .B(\us10\/_0640_ ), .Y(\us10\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1288_ ( .A1(\us10\/_0153_ ), .A2(\us10\/_0056_ ), .B1(\us10\/_0748_ ), .Y(\us10\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1289_ ( .A(\us10\/_0498_ ), .B(\us10\/_0500_ ), .C(\us10\/_0501_ ), .D(\us10\/_0502_ ), .X(\us10\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1290_ ( .A(\us10\/_0490_ ), .B(\us10\/_0492_ ), .C(\us10\/_0497_ ), .D(\us10\/_0503_ ), .X(\us10\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us10/_1291_ ( .A_N(\us10\/_0275_ ), .B(\us10\/_0705_ ), .X(\us10\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1292_ ( .A(\us10\/_0505_ ), .Y(\us10\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1293_ ( .A(\us10\/_0380_ ), .B(\us10\/_0347_ ), .X(\us10\/_0507_ ) );
sky130_fd_sc_hd__o21ai_1 \us10/_1294_ ( .A1(\us10\/_0507_ ), .A2(\us10\/_0093_ ), .B1(\us10\/_0056_ ), .Y(\us10\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1295_ ( .A(\us10\/_0322_ ), .B(\us10\/_0277_ ), .C(\us10\/_0506_ ), .D(\us10\/_0508_ ), .X(\us10\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1296_ ( .A(\us10\/_0084_ ), .B(\us10\/_0705_ ), .X(\us10\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1297_ ( .A1(\us10\/_0733_ ), .A2(\us10\/_0114_ ), .B1(\us10\/_0429_ ), .C1(\us10\/_0511_ ), .Y(\us10\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_1298_ ( .A(\us10\/_0019_ ), .B(\us10\/_0024_ ), .Y(\us10\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1299_ ( .A(\us10\/_0512_ ), .B(\us10\/_0513_ ), .C(\us10\/_0742_ ), .D(\us10\/_0306_ ), .X(\us10\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1300_ ( .A1(\us10\/_0532_ ), .A2(\us10\/_0089_ ), .B1(\us10\/_0154_ ), .C1(\us10\/_0169_ ), .Y(\us10\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us10/_1301_ ( .A1(\us10\/_0749_ ), .A2(\us10\/_0026_ ), .B1(\us10\/_0069_ ), .C1(\us10\/_0032_ ), .X(\us10\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us10/_1302_ ( .A1(\us10\/_0324_ ), .A2(\us10\/_0355_ ), .B1(\us10\/_0330_ ), .B2(\us10\/_0727_ ), .X(\us10\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us10/_1303_ ( .A(\us10\/_0133_ ), .B(\us10\/_0516_ ), .C(\us10\/_0517_ ), .Y(\us10\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1304_ ( .A(\us10\/_0509_ ), .B(\us10\/_0514_ ), .C(\us10\/_0515_ ), .D(\us10\/_0518_ ), .X(\us10\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1305_ ( .A(\us10\/_0746_ ), .B(\us10\/_0072_ ), .Y(\us10\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1306_ ( .A1(\us10\/_0083_ ), .A2(\us10\/_0070_ ), .B1(\us10\/_0043_ ), .B2(\us10\/_0193_ ), .Y(\us10\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1307_ ( .A(\us10\/_0311_ ), .B(\us10\/_0520_ ), .C(\us10\/_0332_ ), .D(\us10\/_0522_ ), .X(\us10\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1308_ ( .A(\us10\/_0129_ ), .B(\us10\/_0218_ ), .X(\us10\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_1309_ ( .A(\us10\/_0235_ ), .B(\us10\/_0524_ ), .Y(\us10\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us10/_1310_ ( .A(\us10\/_0081_ ), .B(\us10\/_0085_ ), .Y(\us10\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1311_ ( .A1(\us10\/_0051_ ), .A2(\us10\/_0045_ ), .B1(\us10\/_0130_ ), .B2(\us10\/_0094_ ), .Y(\us10\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1312_ ( .A(\us10\/_0523_ ), .B(\us10\/_0525_ ), .C(\us10\/_0526_ ), .D(\us10\/_0527_ ), .X(\us10\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us10/_1313_ ( .A_N(\us10\/_0250_ ), .B(\us10\/_0521_ ), .Y(\us10\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1314_ ( .A(\us10\/_0128_ ), .B(\us10\/_0020_ ), .X(\us10\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1315_ ( .A(\us10\/_0530_ ), .Y(\us10\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1316_ ( .A(\us10\/_0099_ ), .B(\us10\/_0058_ ), .X(\us10\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1317_ ( .A(\us10\/_0533_ ), .Y(\us10\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us10/_1318_ ( .A_N(\us10\/_0529_ ), .B(\us10\/_0531_ ), .C(\us10\/_0534_ ), .D(\us10\/_0192_ ), .X(\us10\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1319_ ( .A(\us10\/_0445_ ), .B(\us10\/_0078_ ), .X(\us10\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us10/_1320_ ( .A1(\us10\/_0750_ ), .A2(\us10\/_0079_ ), .B1(\us10\/_0129_ ), .B2(\us10\/_0705_ ), .X(\us10\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1321_ ( .A1(\us10\/_0161_ ), .A2(\us10\/_0032_ ), .B1(\us10\/_0536_ ), .C1(\us10\/_0537_ ), .Y(\us10\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us10/_1322_ ( .A1(\us10\/_0746_ ), .A2(\us10\/_0162_ ), .B1(\us10\/_0079_ ), .B2(\us10\/_0043_ ), .X(\us10\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1323_ ( .A1(\us10\/_0093_ ), .A2(\us10\/_0029_ ), .B1(\us10\/_0240_ ), .C1(\us10\/_0539_ ), .Y(\us10\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1324_ ( .A(\us10\/_0445_ ), .B(\us10\/_0043_ ), .X(\us10\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us10/_1325_ ( .A1(\us10\/_0142_ ), .A2(\us10\/_0150_ ), .B1(\us10\/_0023_ ), .B2(\us10\/_0137_ ), .X(\us10\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1326_ ( .A1(\us10\/_0279_ ), .A2(\us10\/_0051_ ), .B1(\us10\/_0541_ ), .C1(\us10\/_0542_ ), .Y(\us10\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1327_ ( .A(\us10\/_0159_ ), .B(\us10\/_0036_ ), .X(\us10\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us10/_1328_ ( .A1(\us10\/_0282_ ), .A2(\us10\/_0445_ ), .B1(\us10\/_0027_ ), .X(\us10\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1329_ ( .A1(\us10\/_0091_ ), .A2(\us10\/_0128_ ), .B1(\us10\/_0545_ ), .C1(\us10\/_0546_ ), .Y(\us10\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1330_ ( .A(\us10\/_0538_ ), .B(\us10\/_0540_ ), .C(\us10\/_0544_ ), .D(\us10\/_0547_ ), .X(\us10\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1331_ ( .A(\us10\/_0099_ ), .B(\us10\/_0193_ ), .X(\us10\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us10/_1332_ ( .A(\us10\/_0549_ ), .B(\us10\/_0186_ ), .C(\us10\/_0187_ ), .Y(\us10\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1333_ ( .A(\us10\/_0062_ ), .B(\us10\/_0347_ ), .C(\us10\/_0749_ ), .D(\us10\/_0694_ ), .X(\us10\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1334_ ( .A1(\us10\/_0130_ ), .A2(\us10\/_0218_ ), .B1(\us10\/_0551_ ), .C1(\us10\/_0101_ ), .Y(\us10\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1335_ ( .A(\us10\/_0139_ ), .B(\us10\/_0640_ ), .Y(\us10\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1336_ ( .A1(\us10\/_0752_ ), .A2(\us10\/_0672_ ), .B1(\us10\/_0084_ ), .B2(\us10\/_0099_ ), .Y(\us10\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1337_ ( .A(\us10\/_0550_ ), .B(\us10\/_0552_ ), .C(\us10\/_0553_ ), .D(\us10\/_0555_ ), .X(\us10\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1338_ ( .A(\us10\/_0528_ ), .B(\us10\/_0535_ ), .C(\us10\/_0548_ ), .D(\us10\/_0556_ ), .X(\us10\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us10/_1339_ ( .A(\us10\/_0504_ ), .B(\us10\/_0519_ ), .C(\us10\/_0557_ ), .Y(\us10\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1340_ ( .A(\us10\/_0055_ ), .B(\us10\/_0507_ ), .X(\us10\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us10/_1341_ ( .A_N(\us10\/_0558_ ), .B(\us10\/_0408_ ), .C(\us10\/_0451_ ), .D(\us10\/_0452_ ), .X(\us10\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1342_ ( .A(\us10\/_0549_ ), .Y(\us10\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1343_ ( .A(\us10\/_0559_ ), .B(\us10\/_0403_ ), .C(\us10\/_0560_ ), .D(\us10\/_0371_ ), .X(\us10\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1344_ ( .A(\us10\/_0181_ ), .B(\us10\/_0178_ ), .X(\us10\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1345_ ( .A(\us10\/_0562_ ), .B(\us10\/_0552_ ), .C(\us10\/_0553_ ), .D(\us10\/_0555_ ), .X(\us10\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1346_ ( .A(\us10\/_0029_ ), .B(\us10\/_0020_ ), .Y(\us10\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1347_ ( .A(\us10\/_0051_ ), .B(\us10\/_0130_ ), .X(\us10\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1348_ ( .A(\us10\/_0566_ ), .Y(\us10\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1349_ ( .A(\us10\/_0159_ ), .B(\us10\/_0423_ ), .X(\us10\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1350_ ( .A1(\us10\/_0752_ ), .A2(\us10\/_0640_ ), .B1(\us10\/_0568_ ), .B2(\us10\/_0175_ ), .Y(\us10\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1351_ ( .A(\us10\/_0076_ ), .B(\us10\/_0565_ ), .C(\us10\/_0567_ ), .D(\us10\/_0569_ ), .X(\us10\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us10/_1352_ ( .A1(\us10\/_0036_ ), .A2(\us10\/_0142_ ), .B1(\us10\/_0161_ ), .X(\us10\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1353_ ( .A(\us10\/_0099_ ), .B(\us10\/_0672_ ), .Y(\us10\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us10/_1354_ ( .A(\us10\/_0420_ ), .B(\us10\/_0571_ ), .C_N(\us10\/_0572_ ), .Y(\us10\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1355_ ( .A(\us10\/_0051_ ), .B(\us10\/_0746_ ), .Y(\us10\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1356_ ( .A(\us10\/_0574_ ), .B(\us10\/_0319_ ), .C(\us10\/_0320_ ), .D(\us10\/_0411_ ), .X(\us10\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1357_ ( .A(\us10\/_0736_ ), .B(\us10\/_0035_ ), .Y(\us10\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1358_ ( .A(\us10\/_0736_ ), .B(\us10\/_0030_ ), .Y(\us10\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1359_ ( .A(\us10\/_0298_ ), .B(\us10\/_0208_ ), .C(\us10\/_0577_ ), .D(\us10\/_0578_ ), .X(\us10\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1360_ ( .A1(\us10\/_0020_ ), .A2(\us10\/_0137_ ), .B1(\us10\/_0261_ ), .B2(\us10\/_0128_ ), .Y(\us10\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1361_ ( .A(\us10\/_0573_ ), .B(\us10\/_0576_ ), .C(\us10\/_0579_ ), .D(\us10\/_0580_ ), .X(\us10\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1362_ ( .A(\us10\/_0561_ ), .B(\us10\/_0563_ ), .C(\us10\/_0570_ ), .D(\us10\/_0581_ ), .X(\us10\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1363_ ( .A(\us10\/_0128_ ), .B(\us10\/_0193_ ), .X(\us10\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1364_ ( .A(\us10\/_0083_ ), .B(\us10\/_0162_ ), .X(\us10\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us10/_1365_ ( .A(\us10\/_0583_ ), .B(\us10\/_0584_ ), .C_N(\us10\/_0437_ ), .Y(\us10\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us10/_1366_ ( .A(\us10\/_0150_ ), .B(\us10\/_0118_ ), .C(\us10\/_0380_ ), .Y(\us10\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us10/_1367_ ( .A_N(\us10\/_0182_ ), .B(\us10\/_0587_ ), .C(\us10\/_0323_ ), .X(\us10\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1368_ ( .A1(\us10\/_0575_ ), .A2(\us10\/_0153_ ), .B1(\us10\/_0727_ ), .B2(\us10\/_0058_ ), .Y(\us10\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1369_ ( .A1(\us10\/_0218_ ), .A2(\us10\/_0064_ ), .B1(\us10\/_0134_ ), .B2(\us10\/_0255_ ), .Y(\us10\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1370_ ( .A(\us10\/_0585_ ), .B(\us10\/_0588_ ), .C(\us10\/_0589_ ), .D(\us10\/_0590_ ), .X(\us10\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us10/_1371_ ( .A1(\us10\/_0091_ ), .A2(\us10\/_0139_ ), .B1(\us10\/_0250_ ), .Y(\us10\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1372_ ( .A1(\us10\/_0092_ ), .A2(\us10\/_0739_ ), .B1(\us10\/_0324_ ), .B2(\us10\/_0029_ ), .Y(\us10\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1373_ ( .A1(\us10\/_0144_ ), .A2(\us10\/_0153_ ), .B1(\us10\/_0683_ ), .B2(\us10\/_0056_ ), .Y(\us10\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1374_ ( .A1(\us10\/_0091_ ), .A2(\us10\/_0218_ ), .B1(\us10\/_0330_ ), .B2(\us10\/_0056_ ), .Y(\us10\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1375_ ( .A(\us10\/_0592_ ), .B(\us10\/_0593_ ), .C(\us10\/_0594_ ), .D(\us10\/_0595_ ), .X(\us10\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1376_ ( .A(\us10\/_0218_ ), .B(\us10\/_0144_ ), .Y(\us10\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1377_ ( .A(\us10\/_0312_ ), .B(\us10\/_0598_ ), .Y(\us10\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1378_ ( .A(\us10\/_0575_ ), .B(\us10\/_0147_ ), .Y(\us10\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1379_ ( .A1(\us10\/_0293_ ), .A2(\us10\/_0137_ ), .B1(\us10\/_0093_ ), .B2(\us10\/_0739_ ), .Y(\us10\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1380_ ( .A1(\us10\/_0734_ ), .A2(\us10\/_0531_ ), .B1(\us10\/_0600_ ), .C1(\us10\/_0601_ ), .Y(\us10\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1381_ ( .A1(\us10\/_0153_ ), .A2(\us10\/_0261_ ), .B1(\us10\/_0599_ ), .C1(\us10\/_0602_ ), .Y(\us10\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1382_ ( .A(\us10\/_0591_ ), .B(\us10\/_0596_ ), .C(\us10\/_0174_ ), .D(\us10\/_0603_ ), .X(\us10\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1383_ ( .A(\us10\/_0029_ ), .B(\us10\/_0144_ ), .Y(\us10\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1384_ ( .A(\us10\/_0113_ ), .B(\us10\/_0018_ ), .Y(\us10\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1385_ ( .A(\us10\/_0381_ ), .B(\us10\/_0605_ ), .C(\us10\/_0361_ ), .D(\us10\/_0606_ ), .X(\us10\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1386_ ( .A1(\us10\/_0016_ ), .A2(\us10\/_0727_ ), .B1(\us10\/_0733_ ), .Y(\us10\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1387_ ( .A1(\us10\/_0586_ ), .A2(\us10\/_0159_ ), .B1(\us10\/_0083_ ), .B2(\us10\/_0750_ ), .Y(\us10\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1388_ ( .A1(\us10\/_0142_ ), .A2(\us10\/_0162_ ), .B1(\us10\/_0079_ ), .B2(\us10\/_0055_ ), .Y(\us10\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1389_ ( .A(\us10\/_0610_ ), .B(\us10\/_0611_ ), .C(\us10\/_0105_ ), .D(\us10\/_0106_ ), .X(\us10\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1390_ ( .A1(\us10\/_0094_ ), .A2(\us10\/_0302_ ), .B1(\us10\/_0324_ ), .B2(\us10\/_0089_ ), .Y(\us10\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1391_ ( .A(\us10\/_0607_ ), .B(\us10\/_0609_ ), .C(\us10\/_0612_ ), .D(\us10\/_0613_ ), .X(\us10\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1392_ ( .A(\us10\/_0041_ ), .B(\us10\/_0170_ ), .X(\us10\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1393_ ( .A(\us10\/_0554_ ), .B(\us10\/_0027_ ), .X(\us10\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1394_ ( .A(\us10\/_0027_ ), .B(\us10\/_0261_ ), .Y(\us10\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us10/_1395_ ( .A_N(\us10\/_0616_ ), .B(\us10\/_0617_ ), .Y(\us10\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1396_ ( .A1(\us10\/_0147_ ), .A2(\us10\/_0302_ ), .B1(\us10\/_0342_ ), .C1(\us10\/_0618_ ), .Y(\us10\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1397_ ( .A(\us10\/_0614_ ), .B(\us10\/_0272_ ), .C(\us10\/_0615_ ), .D(\us10\/_0620_ ), .X(\us10\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us10/_1398_ ( .A(\us10\/_0582_ ), .B(\us10\/_0604_ ), .C(\us10\/_0621_ ), .Y(\us10\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1399_ ( .A1(\us10\/_0084_ ), .A2(\us10\/_0134_ ), .B1(\us10\/_0089_ ), .Y(\us10\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1400_ ( .A1(\us10\/_0144_ ), .A2(\us10\/_0608_ ), .A3(\us10\/_0330_ ), .B1(\us10\/_0089_ ), .Y(\us10\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1401_ ( .A1(\us10\/_0197_ ), .A2(\us10\/_0130_ ), .A3(\us10\/_0110_ ), .B1(\us10\/_0094_ ), .Y(\us10\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1402_ ( .A(\us10\/_0432_ ), .B(\us10\/_0622_ ), .C(\us10\/_0623_ ), .D(\us10\/_0624_ ), .X(\us10\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us10/_1403_ ( .A1(\us10\/_0554_ ), .A2(\us10\/_0018_ ), .A3(\us10\/_0023_ ), .B1(\us10\/_0161_ ), .X(\us10\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us10/_1404_ ( .A_N(\us10\/_0269_ ), .B(\us10\/_0170_ ), .X(\us10\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1405_ ( .A1(\us10\/_0109_ ), .A2(\us10\/_0064_ ), .A3(\us10\/_0733_ ), .B1(\us10\/_0355_ ), .Y(\us10\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us10/_1406_ ( .A_N(\us10\/_0626_ ), .B(\us10\/_0627_ ), .C(\us10\/_0353_ ), .D(\us10\/_0628_ ), .X(\us10\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1407_ ( .A1(\us10\/_0091_ ), .A2(\us10\/_0110_ ), .A3(\us10\/_0176_ ), .B1(\us10\/_0139_ ), .Y(\us10\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1408_ ( .A1(\us10\/_0020_ ), .A2(\us10\/_0261_ ), .B1(\us10\/_0147_ ), .Y(\us10\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1409_ ( .A(\us10\/_0631_ ), .B(\us10\/_0344_ ), .C(\us10\/_0421_ ), .D(\us10\/_0632_ ), .X(\us10\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us10/_1410_ ( .A1(\us10\/_0325_ ), .A2(\us10\/_0734_ ), .B1(\us10\/_0038_ ), .C1(\us10\/_0113_ ), .X(\us10\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1411_ ( .A1(\us10\/_0134_ ), .A2(\us10\/_0114_ ), .B1(\us10\/_0221_ ), .C1(\us10\/_0634_ ), .Y(\us10\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us10/_1412_ ( .A(\us10\/_0119_ ), .B_N(\us10\/_0111_ ), .Y(\us10\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1413_ ( .A1(\us10\/_0032_ ), .A2(\us10\/_0113_ ), .B1(\us10\/_0636_ ), .C1(\us10\/_0400_ ), .Y(\us10\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1414_ ( .A1(\us10\/_0732_ ), .A2(\us10\/_0293_ ), .A3(\us10\/_0251_ ), .B1(\us10\/_0099_ ), .Y(\us10\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1415_ ( .A(\us10\/_0189_ ), .B(\us10\/_0635_ ), .C(\us10\/_0637_ ), .D(\us10\/_0638_ ), .X(\us10\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1416_ ( .A(\us10\/_0625_ ), .B(\us10\/_0630_ ), .C(\us10\/_0633_ ), .D(\us10\/_0639_ ), .X(\us10\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1417_ ( .A(\us10\/_0746_ ), .B(\us10\/_0738_ ), .X(\us10\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1418_ ( .A(\us10\/_0736_ ), .B(\us10\/_0731_ ), .X(\us10\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us10/_1419_ ( .A_N(\us10\/_0643_ ), .B(\us10\/_0577_ ), .Y(\us10\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1420_ ( .A1(\us10\/_0084_ ), .A2(\us10\/_0739_ ), .B1(\us10\/_0642_ ), .C1(\us10\/_0644_ ), .Y(\us10\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1421_ ( .A1(\us10\/_0050_ ), .A2(\us10\/_0543_ ), .B1(\us10\/_0194_ ), .C1(\us10\/_0738_ ), .Y(\us10\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1422_ ( .A(\us10\/_0646_ ), .B(\us10\/_0232_ ), .C(\us10\/_0417_ ), .D(\us10\/_0578_ ), .X(\us10\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1423_ ( .A1(\us10\/_0064_ ), .A2(\us10\/_0733_ ), .B1(\us10\/_0727_ ), .Y(\us10\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1424_ ( .A1(\us10\/_0193_ ), .A2(\us10\/_0276_ ), .B1(\us10\/_0727_ ), .Y(\us10\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1425_ ( .A(\us10\/_0645_ ), .B(\us10\/_0647_ ), .C(\us10\/_0648_ ), .D(\us10\/_0649_ ), .X(\us10\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1426_ ( .A1(\us10\/_0325_ ), .A2(\us10\/_0734_ ), .B1(\us10\/_0038_ ), .C1(\us10\/_0029_ ), .Y(\us10\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1427_ ( .A1(\us10\/_0543_ ), .A2(\us10\/_0216_ ), .B1(\us10\/_0423_ ), .C1(\us10\/_0029_ ), .Y(\us10\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1428_ ( .A(\us10\/_0652_ ), .B(\us10\/_0653_ ), .X(\us10\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1429_ ( .A1(\us10\/_0733_ ), .A2(\us10\/_0748_ ), .A3(\us10\/_0324_ ), .B1(\us10\/_0016_ ), .Y(\us10\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1430_ ( .A1(\us10\/_0640_ ), .A2(\us10\/_0193_ ), .A3(\us10\/_0091_ ), .B1(\us10\/_0016_ ), .Y(\us10\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1431_ ( .A1(\us10\/_0102_ ), .A2(\us10\/_0301_ ), .B1(\sa10\[3\] ), .C1(\us10\/_0029_ ), .Y(\us10\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1432_ ( .A(\us10\/_0654_ ), .B(\us10\/_0655_ ), .C(\us10\/_0656_ ), .D(\us10\/_0657_ ), .X(\us10\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1433_ ( .A1(\us10\/_0118_ ), .A2(\us10\/_0050_ ), .B1(\us10\/_0038_ ), .C1(\us10\/_0489_ ), .Y(\us10\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us10/_1434_ ( .A_N(\us10\/_0250_ ), .B(\us10\/_0465_ ), .C(\us10\/_0659_ ), .X(\us10\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1435_ ( .A1(\us10\/_0683_ ), .A2(\us10\/_0324_ ), .B1(\us10\/_0255_ ), .Y(\us10\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1436_ ( .A1(\us10\/_0032_ ), .A2(\us10\/_0193_ ), .A3(\us10\/_0048_ ), .B1(\us10\/_0255_ ), .Y(\us10\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1437_ ( .A1(\us10\/_0144_ ), .A2(\us10\/_0586_ ), .A3(\us10\/_0048_ ), .B1(\us10\/_0218_ ), .Y(\us10\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1438_ ( .A(\us10\/_0660_ ), .B(\us10\/_0661_ ), .C(\us10\/_0663_ ), .D(\us10\/_0664_ ), .X(\us10\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1439_ ( .A1(\us10\/_0091_ ), .A2(\us10\/_0276_ ), .B1(\us10\/_0060_ ), .Y(\us10\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1440_ ( .A1(\us10\/_0144_ ), .A2(\us10\/_0608_ ), .B1(\us10\/_0056_ ), .Y(\us10\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1441_ ( .A1(\us10\/_0423_ ), .A2(\us10\/_0038_ ), .B1(\us10\/_0102_ ), .C1(\us10\/_0060_ ), .Y(\us10\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1442_ ( .A1(\sa10\[1\] ), .A2(\us10\/_0734_ ), .B1(\us10\/_0109_ ), .C1(\us10\/_0056_ ), .Y(\us10\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1443_ ( .A(\us10\/_0666_ ), .B(\us10\/_0667_ ), .C(\us10\/_0668_ ), .D(\us10\/_0669_ ), .X(\us10\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1444_ ( .A(\us10\/_0650_ ), .B(\us10\/_0658_ ), .C(\us10\/_0665_ ), .D(\us10\/_0670_ ), .X(\us10\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us10/_1445_ ( .A(\us10\/_0641_ ), .B(\us10\/_0174_ ), .C(\us10\/_0671_ ), .Y(\us10\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us10/_1446_ ( .A(\us10\/_0049_ ), .B(\us10\/_0618_ ), .C_N(\us10\/_0052_ ), .Y(\us10\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us10/_1447_ ( .A(\us10\/_0239_ ), .Y(\us10\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1448_ ( .A(\us10\/_0705_ ), .B(\us10\/_0032_ ), .Y(\us10\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1449_ ( .A1(\us10\/_0055_ ), .A2(\us10\/_0732_ ), .B1(\us10\/_0036_ ), .B2(\us10\/_0705_ ), .Y(\us10\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1450_ ( .A1(\us10\/_0304_ ), .A2(\us10\/_0732_ ), .B1(\us10\/_0048_ ), .B2(\us10\/_0750_ ), .Y(\us10\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1451_ ( .A(\us10\/_0674_ ), .B(\us10\/_0675_ ), .C(\us10\/_0676_ ), .D(\us10\/_0677_ ), .X(\us10\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us10/_1452_ ( .A_N(\us10\/_0584_ ), .B(\us10\/_0283_ ), .X(\us10\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1453_ ( .A(\us10\/_0673_ ), .B(\us10\/_0678_ ), .C(\us10\/_0679_ ), .D(\us10\/_0508_ ), .X(\us10\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1454_ ( .A1(\us10\/_0016_ ), .A2(\us10\/_0733_ ), .B1(\us10\/_0355_ ), .B2(\us10\/_0092_ ), .Y(\us10\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1455_ ( .A(\us10\/_0681_ ), .B(\us10\/_0034_ ), .X(\us10\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us10/_1456_ ( .A1(\us10\/_0330_ ), .A2(\us10\/_0139_ ), .B1(\us10\/_0324_ ), .B2(\us10\/_0089_ ), .X(\us10\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1457_ ( .A1(\us10\/_0146_ ), .A2(\us10\/_0147_ ), .B1(\us10\/_0133_ ), .C1(\us10\/_0684_ ), .Y(\us10\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1458_ ( .A(\us10\/_0113_ ), .B(\us10\/_0251_ ), .Y(\us10\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us10/_1459_ ( .A_N(\us10\/_0463_ ), .B(\us10\/_0686_ ), .C(\us10\/_0383_ ), .D(\us10\/_0464_ ), .X(\us10\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1460_ ( .A1(\us10\/_0051_ ), .A2(\us10\/_0293_ ), .B1(\us10\/_0084_ ), .B2(\us10\/_0705_ ), .Y(\us10\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1461_ ( .A1(\us10\/_0018_ ), .A2(\us10\/_0072_ ), .B1(\us10\/_0134_ ), .B2(\us10\/_0078_ ), .Y(\us10\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1462_ ( .A(\us10\/_0687_ ), .B(\us10\/_0236_ ), .C(\us10\/_0688_ ), .D(\us10\/_0689_ ), .X(\us10\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1463_ ( .A(\us10\/_0680_ ), .B(\us10\/_0682_ ), .C(\us10\/_0685_ ), .D(\us10\/_0690_ ), .X(\us10\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us10/_1464_ ( .A1(\us10\/_0532_ ), .A2(\us10\/_0380_ ), .B1(\us10\/_0102_ ), .C1(\us10\/_0355_ ), .X(\us10\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us10/_1465_ ( .A(\us10\/_0692_ ), .B(\us10\/_0338_ ), .C(\us10\/_0644_ ), .Y(\us10\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1466_ ( .A(\us10\/_0016_ ), .B(\us10\/_0020_ ), .Y(\us10\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1467_ ( .A1(\us10\/_0032_ ), .A2(\us10\/_0137_ ), .B1(\us10\/_0279_ ), .B2(\us10\/_0094_ ), .Y(\us10\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1468_ ( .A1(\us10\/_0575_ ), .A2(\us10\/_0153_ ), .B1(\us10\/_0161_ ), .B2(\us10\/_0293_ ), .Y(\us10\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1469_ ( .A(\us10\/_0259_ ), .B(\us10\/_0695_ ), .C(\us10\/_0696_ ), .D(\us10\/_0697_ ), .X(\us10\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us10/_1470_ ( .A1(\us10\/_0255_ ), .A2(\us10\/_0640_ ), .B1(\us10\/_0016_ ), .B2(\us10\/_0193_ ), .X(\us10\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1471_ ( .A1(\us10\/_0060_ ), .A2(\us10\/_0176_ ), .B1(\us10\/_0699_ ), .C1(\us10\/_0177_ ), .Y(\us10\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1472_ ( .A1(\us10\/_0091_ ), .A2(\us10\/_0218_ ), .B1(\us10\/_0092_ ), .B2(\us10\/_0705_ ), .Y(\us10\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us10/_1473_ ( .A1(\us10\/_0705_ ), .A2(\us10\/_0683_ ), .B1(\us10\/_0093_ ), .B2(\us10\/_0114_ ), .Y(\us10\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us10/_1474_ ( .A1(\us10\/_0683_ ), .A2(\us10\/_0084_ ), .B1(\us10\/_0094_ ), .Y(\us10\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us10/_1475_ ( .A1(\us10\/_0543_ ), .A2(\us10\/_0216_ ), .B1(\us10\/_0038_ ), .C1(\us10\/_0056_ ), .Y(\us10\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1476_ ( .A(\us10\/_0701_ ), .B(\us10\/_0702_ ), .C(\us10\/_0703_ ), .D(\us10\/_0704_ ), .X(\us10\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1477_ ( .A(\us10\/_0693_ ), .B(\us10\/_0698_ ), .C(\us10\/_0700_ ), .D(\us10\/_0706_ ), .X(\us10\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us10/_1478_ ( .A1(\us10\/_0113_ ), .A2(\us10\/_0640_ ), .B1(\us10\/_0099_ ), .B2(\us10\/_0058_ ), .X(\us10\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us10/_1479_ ( .A(\us10\/_0407_ ), .B(\us10\/_0708_ ), .C(\us10\/_0529_ ), .Y(\us10\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1480_ ( .A(\us10\/_0568_ ), .B(\us10\/_0175_ ), .Y(\us10\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us10/_1481_ ( .A1(\us10\/_0029_ ), .A2(\us10\/_0114_ ), .A3(\us10\/_0051_ ), .B1(\us10\/_0130_ ), .Y(\us10\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1482_ ( .A(\us10\/_0709_ ), .B(\us10\/_0550_ ), .C(\us10\/_0710_ ), .D(\us10\/_0711_ ), .X(\us10\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us10/_1483_ ( .A1(\us10\/_0114_ ), .A2(\us10\/_0064_ ), .B1(\us10\/_0261_ ), .B2(\us10\/_0089_ ), .X(\us10\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1484_ ( .A1(\us10\/_0355_ ), .A2(\us10\/_0261_ ), .B1(\us10\/_0198_ ), .C1(\us10\/_0713_ ), .Y(\us10\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1485_ ( .A(\us10\/_0586_ ), .B(\us10\/_0489_ ), .Y(\us10\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us10/_1486_ ( .A_N(\us10\/_0541_ ), .B(\us10\/_0267_ ), .C(\us10\/_0715_ ), .D(\us10\/_0320_ ), .X(\us10\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1487_ ( .A(\us10\/_0586_ ), .B(\us10\/_0070_ ), .Y(\us10\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us10/_1488_ ( .A_N(\us10\/_0211_ ), .B(\us10\/_0155_ ), .C(\us10\/_0202_ ), .D(\us10\/_0718_ ), .X(\us10\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us10/_1489_ ( .A(\us10\/_0150_ ), .B(\us10\/_0216_ ), .C(\us10\/_0380_ ), .Y(\us10\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us10/_1490_ ( .A(\us10\/_0411_ ), .B(\us10\/_0720_ ), .X(\us10\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us10/_1491_ ( .A1(\us10\/_0018_ ), .A2(\us10\/_0023_ ), .B1(\us10\/_0078_ ), .X(\us10\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us10/_1492_ ( .A1(\us10\/_0134_ ), .A2(\us10\/_0738_ ), .B1(\us10\/_0101_ ), .C1(\us10\/_0722_ ), .Y(\us10\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1493_ ( .A(\us10\/_0717_ ), .B(\us10\/_0719_ ), .C(\us10\/_0721_ ), .D(\us10\/_0723_ ), .X(\us10\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us10/_1494_ ( .A(\us10\/_0739_ ), .B(\us10\/_0193_ ), .Y(\us10\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1495_ ( .A(\us10\/_0344_ ), .B(\us10\/_0184_ ), .C(\us10\/_0449_ ), .D(\us10\/_0725_ ), .X(\us10\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us10/_1496_ ( .A(\us10\/_0712_ ), .B(\us10\/_0714_ ), .C(\us10\/_0724_ ), .D(\us10\/_0726_ ), .X(\us10\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \us10/_1497_ ( .A(\us10\/_0691_ ), .B(\us10\/_0707_ ), .C(\us10\/_0728_ ), .Y(\us10\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \us11/_0753_ ( .A(\sa11\[2\] ), .B_N(\sa11\[3\] ), .Y(\us11\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \us11/_0755_ ( .A(\sa11\[1\] ), .B(\sa11\[0\] ), .X(\us11\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us11/_0756_ ( .A(\us11\/_0096_ ), .B(\us11\/_0118_ ), .X(\us11\/_0129_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0757_ ( .A(\sa11\[7\] ), .B(\sa11\[6\] ), .X(\us11\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_0758_ ( .A(\sa11\[4\] ), .B(\sa11\[5\] ), .Y(\us11\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0759_ ( .A(\us11\/_0140_ ), .B(\us11\/_0151_ ), .X(\us11\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0761_ ( .A(\us11\/_0129_ ), .B(\us11\/_0162_ ), .X(\us11\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0762_ ( .A(\us11\/_0096_ ), .X(\us11\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \us11/_0763_ ( .A(\sa11\[1\] ), .B_N(\sa11\[0\] ), .Y(\us11\/_0205_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0764_ ( .A(\us11\/_0205_ ), .X(\us11\/_0216_ ) );
sky130_fd_sc_hd__and3_1 \us11/_0765_ ( .A(\us11\/_0162_ ), .B(\us11\/_0194_ ), .C(\us11\/_0216_ ), .X(\us11\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us11/_0766_ ( .A(\us11\/_0183_ ), .SLEEP(\us11\/_0227_ ), .X(\us11\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \us11/_0767_ ( .A(\sa11\[0\] ), .B_N(\sa11\[1\] ), .Y(\us11\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_0768_ ( .A(\sa11\[2\] ), .B(\sa11\[3\] ), .Y(\us11\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0769_ ( .A(\us11\/_0249_ ), .B(\us11\/_0260_ ), .X(\us11\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0771_ ( .A(\us11\/_0271_ ), .X(\us11\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0772_ ( .A(\us11\/_0162_ ), .X(\us11\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_0773_ ( .A(\us11\/_0293_ ), .B(\us11\/_0304_ ), .Y(\us11\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us11/_0774_ ( .A(\sa11\[1\] ), .Y(\us11\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us11/_0776_ ( .A(\sa11\[0\] ), .Y(\us11\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0777_ ( .A(\sa11\[2\] ), .B(\sa11\[3\] ), .X(\us11\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0779_ ( .A(\us11\/_0358_ ), .X(\us11\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_0780_ ( .A1(\us11\/_0325_ ), .A2(\us11\/_0347_ ), .B1(\us11\/_0380_ ), .C1(\us11\/_0304_ ), .Y(\us11\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us11/_0781_ ( .A_N(\us11\/_0238_ ), .B(\us11\/_0314_ ), .C(\us11\/_0391_ ), .X(\us11\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us11/_0782_ ( .A(\sa11\[3\] ), .B_N(\sa11\[2\] ), .Y(\us11\/_0412_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0783_ ( .A(\us11\/_0412_ ), .X(\us11\/_0423_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0784_ ( .A(\us11\/_0423_ ), .B(\us11\/_0205_ ), .X(\us11\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \us11/_0787_ ( .A(\sa11\[5\] ), .B_N(\sa11\[4\] ), .Y(\us11\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0788_ ( .A(\us11\/_0467_ ), .B(\us11\/_0140_ ), .X(\us11\/_0478_ ) );
sky130_fd_sc_hd__buf_2 \us11/_0790_ ( .A(\us11\/_0478_ ), .X(\us11\/_0499_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_0791_ ( .A(\us11\/_0134_ ), .B(\us11\/_0499_ ), .Y(\us11\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_0792_ ( .A(\us11\/_0478_ ), .B(\us11\/_0271_ ), .Y(\us11\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0793_ ( .A(\us11\/_0194_ ), .X(\us11\/_0532_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0794_ ( .A(\us11\/_0249_ ), .X(\us11\/_0543_ ) );
sky130_fd_sc_hd__and2_1 \us11/_0795_ ( .A(\us11\/_0543_ ), .B(\us11\/_0358_ ), .X(\us11\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0797_ ( .A(\us11\/_0554_ ), .X(\us11\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us11/_0798_ ( .A(\us11\/_0216_ ), .B(\us11\/_0358_ ), .X(\us11\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0800_ ( .A(\us11\/_0586_ ), .X(\us11\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_0801_ ( .A1(\us11\/_0532_ ), .A2(\us11\/_0575_ ), .A3(\us11\/_0608_ ), .B1(\us11\/_0499_ ), .Y(\us11\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us11/_0802_ ( .A(\us11\/_0401_ ), .B(\us11\/_0510_ ), .C(\us11\/_0521_ ), .D(\us11\/_0619_ ), .X(\us11\/_0629_ ) );
sky130_fd_sc_hd__and2_1 \us11/_0803_ ( .A(\us11\/_0358_ ), .B(\sa11\[1\] ), .X(\us11\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0805_ ( .A(\us11\/_0205_ ), .B(\us11\/_0260_ ), .X(\us11\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0807_ ( .A(\us11\/_0662_ ), .X(\us11\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us11/_0808_ ( .A(\sa11\[6\] ), .B_N(\sa11\[7\] ), .Y(\us11\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \us11/_0809_ ( .A(\us11\/_0467_ ), .B(\us11\/_0694_ ), .X(\us11\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0811_ ( .A(\us11\/_0705_ ), .X(\us11\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_0812_ ( .A1(\us11\/_0640_ ), .A2(\us11\/_0293_ ), .A3(\us11\/_0683_ ), .B1(\us11\/_0727_ ), .Y(\us11\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_0813_ ( .A(\sa11\[1\] ), .B(\sa11\[0\] ), .Y(\us11\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0814_ ( .A(\us11\/_0730_ ), .B(\us11\/_0260_ ), .X(\us11\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0815_ ( .A(\us11\/_0731_ ), .X(\us11\/_0732_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0816_ ( .A(\us11\/_0732_ ), .X(\us11\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0817_ ( .A(\sa11\[0\] ), .X(\us11\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us11/_0818_ ( .A1(\us11\/_0325_ ), .A2(\us11\/_0734_ ), .B1(\us11\/_0423_ ), .X(\us11\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0819_ ( .A(\us11\/_0694_ ), .B(\us11\/_0151_ ), .X(\us11\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0821_ ( .A(\us11\/_0736_ ), .X(\us11\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0822_ ( .A(\us11\/_0738_ ), .X(\us11\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_0823_ ( .A1(\us11\/_0733_ ), .A2(\us11\/_0735_ ), .A3(\us11\/_0293_ ), .B1(\us11\/_0739_ ), .Y(\us11\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us11/_0824_ ( .A(\us11\/_0730_ ), .B_N(\us11\/_0358_ ), .Y(\us11\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_0825_ ( .A(\us11\/_0741_ ), .B(\us11\/_0739_ ), .Y(\us11\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_0827_ ( .A1(\us11\/_0118_ ), .A2(\us11\/_0216_ ), .B1(\us11\/_0532_ ), .C1(\us11\/_0739_ ), .Y(\us11\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us11/_0828_ ( .A(\us11\/_0729_ ), .B(\us11\/_0740_ ), .C(\us11\/_0742_ ), .D(\us11\/_0744_ ), .X(\us11\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0829_ ( .A(\us11\/_0423_ ), .B(\us11\/_0730_ ), .X(\us11\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0831_ ( .A(\us11\/_0746_ ), .X(\us11\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us11/_0832_ ( .A(\sa11\[4\] ), .B_N(\sa11\[5\] ), .Y(\us11\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0833_ ( .A(\us11\/_0749_ ), .B(\us11\/_0694_ ), .X(\us11\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0835_ ( .A(\us11\/_0750_ ), .X(\us11\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0836_ ( .A(\us11\/_0752_ ), .X(\us11\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0837_ ( .A(\us11\/_0118_ ), .B(\us11\/_0358_ ), .X(\us11\/_0017_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0839_ ( .A(\us11\/_0752_ ), .B(\us11\/_0017_ ), .X(\us11\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0840_ ( .A(\us11\/_0358_ ), .B(\us11\/_0325_ ), .X(\us11\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0842_ ( .A(\us11\/_0096_ ), .B(\us11\/_0205_ ), .X(\us11\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \us11/_0844_ ( .A1(\us11\/_0020_ ), .A2(\us11\/_0022_ ), .B1(\us11\/_0752_ ), .X(\us11\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_0845_ ( .A1(\us11\/_0748_ ), .A2(\us11\/_0016_ ), .B1(\us11\/_0019_ ), .C1(\us11\/_0024_ ), .Y(\us11\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \us11/_0846_ ( .A(\sa11\[4\] ), .B(\sa11\[5\] ), .X(\us11\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0847_ ( .A(\us11\/_0694_ ), .B(\us11\/_0026_ ), .X(\us11\/_0027_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0850_ ( .A(\us11\/_0358_ ), .B(\us11\/_0730_ ), .X(\us11\/_0030_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0852_ ( .A(\us11\/_0030_ ), .X(\us11\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_0853_ ( .A(\us11\/_0247_ ), .B(\us11\/_0032_ ), .Y(\us11\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_0854_ ( .A(\us11\/_0247_ ), .B(\us11\/_0735_ ), .Y(\us11\/_0034_ ) );
sky130_fd_sc_hd__and2_1 \us11/_0855_ ( .A(\us11\/_0118_ ), .B(\us11\/_0260_ ), .X(\us11\/_0035_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0857_ ( .A(\us11\/_0027_ ), .B(\us11\/_0035_ ), .X(\us11\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0858_ ( .A(\us11\/_0260_ ), .X(\us11\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_0859_ ( .A(\us11\/_0038_ ), .B(\us11\/_0347_ ), .Y(\us11\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us11/_0860_ ( .A_N(\us11\/_0039_ ), .B(\us11\/_0027_ ), .X(\us11\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_0861_ ( .A(\us11\/_0037_ ), .B(\us11\/_0040_ ), .Y(\us11\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us11/_0862_ ( .A(\us11\/_0025_ ), .B(\us11\/_0033_ ), .C(\us11\/_0034_ ), .D(\us11\/_0041_ ), .X(\us11\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0863_ ( .A(\us11\/_0749_ ), .B(\us11\/_0140_ ), .X(\us11\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us11/_0865_ ( .A(\sa11\[0\] ), .B(\sa11\[2\] ), .C(\sa11\[3\] ), .X(\us11\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0866_ ( .A(\us11\/_0043_ ), .B(\us11\/_0045_ ), .X(\us11\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0867_ ( .A(\us11\/_0096_ ), .B(\us11\/_0543_ ), .X(\us11\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0869_ ( .A(\us11\/_0047_ ), .B(\us11\/_0043_ ), .X(\us11\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0870_ ( .A(\us11\/_0730_ ), .X(\us11\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0871_ ( .A(\us11\/_0043_ ), .X(\us11\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_0872_ ( .A1(\us11\/_0118_ ), .A2(\us11\/_0050_ ), .B1(\us11\/_0194_ ), .C1(\us11\/_0051_ ), .Y(\us11\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us11/_0873_ ( .A(\us11\/_0046_ ), .B(\us11\/_0049_ ), .C_N(\us11\/_0052_ ), .Y(\us11\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0874_ ( .A(\us11\/_0026_ ), .B(\us11\/_0140_ ), .X(\us11\/_0054_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_0877_ ( .A1(\us11\/_0532_ ), .A2(\us11\/_0575_ ), .B1(\us11\/_0292_ ), .Y(\us11\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0878_ ( .A(\us11\/_0423_ ), .B(\us11\/_0325_ ), .X(\us11\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0880_ ( .A(\us11\/_0051_ ), .X(\us11\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_0881_ ( .A1(\us11\/_0732_ ), .A2(\us11\/_0035_ ), .A3(\us11\/_0058_ ), .B1(\us11\/_0060_ ), .Y(\us11\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0882_ ( .A(\us11\/_0260_ ), .B(\sa11\[1\] ), .X(\us11\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0884_ ( .A(\us11\/_0062_ ), .X(\us11\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_0885_ ( .A1(\us11\/_0064_ ), .A2(\us11\/_0748_ ), .A3(\us11\/_0683_ ), .B1(\us11\/_0292_ ), .Y(\us11\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us11/_0886_ ( .A(\us11\/_0053_ ), .B(\us11\/_0057_ ), .C(\us11\/_0061_ ), .D(\us11\/_0065_ ), .X(\us11\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us11/_0887_ ( .A(\us11\/_0629_ ), .B(\us11\/_0745_ ), .C(\us11\/_0042_ ), .D(\us11\/_0066_ ), .X(\us11\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us11/_0889_ ( .A(\sa11\[7\] ), .B_N(\sa11\[6\] ), .Y(\us11\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0890_ ( .A(\us11\/_0069_ ), .B(\us11\/_0151_ ), .X(\us11\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0892_ ( .A(\us11\/_0070_ ), .X(\us11\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_0893_ ( .A1(\us11\/_0129_ ), .A2(\us11\/_0586_ ), .B1(\us11\/_0072_ ), .Y(\us11\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_0894_ ( .A1(\us11\/_0380_ ), .A2(\us11\/_0347_ ), .B1(\us11\/_0194_ ), .B2(\us11\/_0216_ ), .Y(\us11\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us11/_0895_ ( .A(\us11\/_0074_ ), .B_N(\us11\/_0070_ ), .Y(\us11\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us11/_0896_ ( .A(\us11\/_0073_ ), .SLEEP(\us11\/_0075_ ), .X(\us11\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us11/_0897_ ( .A(\us11\/_0467_ ), .B(\us11\/_0069_ ), .X(\us11\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0898_ ( .A(\us11\/_0077_ ), .X(\us11\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0899_ ( .A(\us11\/_0412_ ), .B(\us11\/_0118_ ), .X(\us11\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0901_ ( .A(\us11\/_0078_ ), .B(\us11\/_0079_ ), .X(\us11\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0902_ ( .A(\us11\/_0412_ ), .B(\us11\/_0249_ ), .X(\us11\/_0082_ ) );
sky130_fd_sc_hd__buf_2 \us11/_0904_ ( .A(\us11\/_0082_ ), .X(\us11\/_0084_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0905_ ( .A(\us11\/_0084_ ), .B(\us11\/_0078_ ), .X(\us11\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us11/_0906_ ( .A1(\sa11\[0\] ), .A2(\us11\/_0325_ ), .B1(\us11\/_0260_ ), .Y(\us11\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us11/_0907_ ( .A_N(\us11\/_0086_ ), .B(\us11\/_0078_ ), .X(\us11\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us11/_0908_ ( .A(\us11\/_0081_ ), .B(\us11\/_0085_ ), .C(\us11\/_0087_ ), .Y(\us11\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0909_ ( .A(\us11\/_0072_ ), .X(\us11\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_0910_ ( .A1(\us11\/_0733_ ), .A2(\us11\/_0748_ ), .A3(\us11\/_0683_ ), .B1(\us11\/_0089_ ), .Y(\us11\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0911_ ( .A(\us11\/_0129_ ), .X(\us11\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0912_ ( .A(\us11\/_0017_ ), .X(\us11\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0913_ ( .A(\us11\/_0022_ ), .X(\us11\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0914_ ( .A(\us11\/_0078_ ), .X(\us11\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_0915_ ( .A1(\us11\/_0091_ ), .A2(\us11\/_0092_ ), .A3(\us11\/_0093_ ), .B1(\us11\/_0094_ ), .Y(\us11\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us11/_0916_ ( .A(\us11\/_0076_ ), .B(\us11\/_0088_ ), .C(\us11\/_0090_ ), .D(\us11\/_0095_ ), .X(\us11\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us11/_0917_ ( .A(\us11\/_0069_ ), .B(\us11\/_0026_ ), .X(\us11\/_0098_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0919_ ( .A(\us11\/_0434_ ), .B(\us11\/_0364_ ), .X(\us11\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0920_ ( .A(\us11\/_0079_ ), .B(\us11\/_0098_ ), .X(\us11\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0921_ ( .A(\us11\/_0325_ ), .X(\us11\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_0922_ ( .A1(\us11\/_0102_ ), .A2(\us11\/_0734_ ), .B1(\us11\/_0038_ ), .C1(\us11\/_0364_ ), .Y(\us11\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us11/_0923_ ( .A(\us11\/_0100_ ), .B(\us11\/_0101_ ), .C_N(\us11\/_0103_ ), .Y(\us11\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_0924_ ( .A1(\us11\/_0554_ ), .A2(\us11\/_0586_ ), .B1(\us11\/_0364_ ), .Y(\us11\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_0925_ ( .A(\us11\/_0129_ ), .B(\us11\/_0364_ ), .Y(\us11\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0926_ ( .A(\us11\/_0105_ ), .B(\us11\/_0106_ ), .X(\us11\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0927_ ( .A(\us11\/_0423_ ), .X(\us11\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us11/_0928_ ( .A(\us11\/_0260_ ), .B(\sa11\[0\] ), .X(\us11\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0929_ ( .A(\us11\/_0069_ ), .B(\us11\/_0749_ ), .X(\us11\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0931_ ( .A(\us11\/_0111_ ), .X(\us11\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0932_ ( .A(\us11\/_0113_ ), .X(\us11\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_0933_ ( .A1(\us11\/_0109_ ), .A2(\us11\/_0110_ ), .B1(\us11\/_0114_ ), .Y(\us11\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us11/_0934_ ( .A(\us11\/_0022_ ), .Y(\us11\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us11/_0935_ ( .A(\us11\/_0554_ ), .Y(\us11\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us11/_0936_ ( .A1(\us11\/_0050_ ), .A2(\us11\/_0118_ ), .B1(\us11\/_0194_ ), .Y(\us11\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us11/_0937_ ( .A(\us11\/_0113_ ), .Y(\us11\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us11/_0938_ ( .A1(\us11\/_0116_ ), .A2(\us11\/_0117_ ), .A3(\us11\/_0119_ ), .B1(\us11\/_0120_ ), .X(\us11\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us11/_0939_ ( .A(\us11\/_0104_ ), .B(\us11\/_0108_ ), .C(\us11\/_0115_ ), .D(\us11\/_0121_ ), .X(\us11\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_0940_ ( .A(\sa11\[7\] ), .B(\sa11\[6\] ), .Y(\us11\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0941_ ( .A(\us11\/_0749_ ), .B(\us11\/_0123_ ), .X(\us11\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0943_ ( .A(\us11\/_0082_ ), .B(\us11\/_0124_ ), .X(\us11\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_0944_ ( .A(\us11\/_0271_ ), .B(\us11\/_0124_ ), .Y(\us11\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0945_ ( .A(\us11\/_0124_ ), .X(\us11\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0946_ ( .A(\us11\/_0260_ ), .B(\us11\/_0325_ ), .X(\us11\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_0948_ ( .A(\us11\/_0128_ ), .B(\us11\/_0130_ ), .Y(\us11\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_0949_ ( .A(\us11\/_0127_ ), .B(\us11\/_0132_ ), .Y(\us11\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us11/_0950_ ( .A(\us11\/_0434_ ), .X(\us11\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_0951_ ( .A(\us11\/_0134_ ), .B(\us11\/_0128_ ), .Y(\us11\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us11/_0952_ ( .A(\us11\/_0126_ ), .B(\us11\/_0133_ ), .C_N(\us11\/_0135_ ), .Y(\us11\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us11/_0953_ ( .A(\us11\/_0026_ ), .B(\us11\/_0123_ ), .X(\us11\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0955_ ( .A(\us11\/_0137_ ), .X(\us11\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_0956_ ( .A1(\us11\/_0110_ ), .A2(\us11\/_0293_ ), .A3(\us11\/_0084_ ), .B1(\us11\/_0139_ ), .Y(\us11\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0957_ ( .A(\us11\/_0096_ ), .B(\us11\/_0730_ ), .X(\us11\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0959_ ( .A(\us11\/_0142_ ), .X(\us11\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_0960_ ( .A1(\us11\/_0020_ ), .A2(\us11\/_0144_ ), .A3(\us11\/_0017_ ), .B1(\us11\/_0139_ ), .Y(\us11\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \us11/_0961_ ( .A(\sa11\[2\] ), .B(\us11\/_0050_ ), .C_N(\sa11\[3\] ), .Y(\us11\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0962_ ( .A(\us11\/_0128_ ), .X(\us11\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_0963_ ( .A1(\us11\/_0146_ ), .A2(\us11\/_0032_ ), .A3(\us11\/_0640_ ), .B1(\us11\/_0147_ ), .Y(\us11\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us11/_0964_ ( .A(\us11\/_0136_ ), .B(\us11\/_0141_ ), .C(\us11\/_0145_ ), .D(\us11\/_0148_ ), .X(\us11\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0965_ ( .A(\us11\/_0123_ ), .B(\us11\/_0151_ ), .X(\us11\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0967_ ( .A(\us11\/_0150_ ), .X(\us11\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \us11/_0968_ ( .A(\us11\/_0150_ ), .B(\us11\/_0062_ ), .X(\us11\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_0969_ ( .A(\us11\/_0079_ ), .B(\us11\/_0150_ ), .Y(\us11\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us11/_0970_ ( .A(\us11\/_0150_ ), .B(\us11\/_0423_ ), .C(\us11\/_0543_ ), .Y(\us11\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_0971_ ( .A(\us11\/_0155_ ), .B(\us11\/_0156_ ), .Y(\us11\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_0972_ ( .A1(\us11\/_0153_ ), .A2(\us11\/_0134_ ), .B1(\us11\/_0154_ ), .C1(\us11\/_0157_ ), .Y(\us11\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0973_ ( .A(\us11\/_0467_ ), .B(\us11\/_0123_ ), .X(\us11\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_0975_ ( .A(\us11\/_0159_ ), .X(\us11\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us11/_0976_ ( .A_N(\us11\/_0119_ ), .B(\us11\/_0161_ ), .X(\us11\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us11/_0977_ ( .A(\us11\/_0163_ ), .Y(\us11\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_0978_ ( .A1(\us11\/_0146_ ), .A2(\us11\/_0575_ ), .A3(\us11\/_0608_ ), .B1(\us11\/_0153_ ), .Y(\us11\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_0979_ ( .A1(\us11\/_0062_ ), .A2(\us11\/_0084_ ), .A3(\us11\/_0134_ ), .B1(\us11\/_0161_ ), .Y(\us11\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us11/_0980_ ( .A(\us11\/_0158_ ), .B(\us11\/_0164_ ), .C(\us11\/_0165_ ), .D(\us11\/_0166_ ), .X(\us11\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us11/_0981_ ( .A(\us11\/_0097_ ), .B(\us11\/_0122_ ), .C(\us11\/_0149_ ), .D(\us11\/_0167_ ), .X(\us11\/_0168_ ) );
sky130_fd_sc_hd__and2_1 \us11/_0982_ ( .A(\us11\/_0662_ ), .B(\us11\/_0150_ ), .X(\us11\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_0983_ ( .A(\us11\/_0154_ ), .B(\us11\/_0169_ ), .Y(\us11\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us11/_0984_ ( .A(\us11\/_0123_ ), .B(\us11\/_0151_ ), .C(\us11\/_0038_ ), .X(\us11\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0985_ ( .A(\us11\/_0170_ ), .B(\us11\/_0171_ ), .X(\us11\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \us11/_0986_ ( .A(\us11\/_0172_ ), .Y(\us11\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \us11/_0987_ ( .A(\us11\/_0067_ ), .B(\us11\/_0168_ ), .C(\us11\/_0174_ ), .Y(\us11\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us11/_0988_ ( .A(\sa11\[1\] ), .B(\sa11\[0\] ), .Y(\us11\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us11/_0989_ ( .A(\us11\/_0175_ ), .B(\us11\/_0358_ ), .X(\us11\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0990_ ( .A(\us11\/_0176_ ), .B(\us11\/_0478_ ), .X(\us11\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_0991_ ( .A(\us11\/_0084_ ), .B(\us11\/_0113_ ), .Y(\us11\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0992_ ( .A(\us11\/_0111_ ), .B(\us11\/_0062_ ), .X(\us11\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0993_ ( .A(\us11\/_0111_ ), .B(\us11\/_0662_ ), .X(\us11\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_0994_ ( .A(\us11\/_0179_ ), .B(\us11\/_0180_ ), .Y(\us11\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0995_ ( .A(\us11\/_0054_ ), .B(\us11\/_0058_ ), .X(\us11\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us11/_0996_ ( .A(\us11\/_0182_ ), .Y(\us11\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us11/_0997_ ( .A_N(\us11\/_0177_ ), .B(\us11\/_0178_ ), .C(\us11\/_0181_ ), .D(\us11\/_0184_ ), .X(\us11\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0998_ ( .A(\us11\/_0098_ ), .B(\us11\/_0741_ ), .X(\us11\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us11/_0999_ ( .A(\us11\/_0047_ ), .B(\us11\/_0098_ ), .X(\us11\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us11/_1000_ ( .A(\us11\/_0186_ ), .B(\us11\/_0187_ ), .X(\us11\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1001_ ( .A(\us11\/_0188_ ), .Y(\us11\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1002_ ( .A(\us11\/_0738_ ), .B(\us11\/_0735_ ), .X(\us11\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1003_ ( .A(\us11\/_0271_ ), .B(\us11\/_0736_ ), .X(\us11\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_1004_ ( .A(\us11\/_0190_ ), .B(\us11\/_0191_ ), .Y(\us11\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us11/_1005_ ( .A(\us11\/_0096_ ), .B(\us11\/_0325_ ), .X(\us11\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1006_ ( .A1(\us11\/_0193_ ), .A2(\us11\/_0176_ ), .B1(\us11\/_0043_ ), .Y(\us11\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1007_ ( .A(\us11\/_0185_ ), .B(\us11\/_0189_ ), .C(\us11\/_0192_ ), .D(\us11\/_0195_ ), .X(\us11\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us11/_1008_ ( .A_N(\sa11\[3\] ), .B(\us11\/_0734_ ), .C(\sa11\[2\] ), .X(\us11\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1009_ ( .A(\us11\/_0137_ ), .B(\us11\/_0197_ ), .X(\us11\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_1010_ ( .A(\us11\/_0198_ ), .B(\us11\/_0040_ ), .Y(\us11\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1011_ ( .A(\us11\/_0293_ ), .B(\us11\/_0137_ ), .X(\us11\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1012_ ( .A(\us11\/_0200_ ), .Y(\us11\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1013_ ( .A(\us11\/_0137_ ), .B(\us11\/_0110_ ), .Y(\us11\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1014_ ( .A(\us11\/_0139_ ), .B(\us11\/_0020_ ), .Y(\us11\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1015_ ( .A(\us11\/_0199_ ), .B(\us11\/_0201_ ), .C(\us11\/_0202_ ), .D(\us11\/_0203_ ), .X(\us11\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us11/_1016_ ( .A1(\us11\/_0532_ ), .A2(\us11\/_0109_ ), .B1(\us11\/_0102_ ), .C1(\us11\/_0727_ ), .X(\us11\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1017_ ( .A(\us11\/_0022_ ), .B(\us11\/_0078_ ), .Y(\us11\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1018_ ( .A(\us11\/_0078_ ), .B(\us11\/_0142_ ), .Y(\us11\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1019_ ( .A(\us11\/_0207_ ), .B(\us11\/_0208_ ), .Y(\us11\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1020_ ( .A1(\us11\/_0094_ ), .A2(\us11\/_0176_ ), .B1(\us11\/_0206_ ), .C1(\us11\/_0209_ ), .Y(\us11\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1021_ ( .A(\us11\/_0662_ ), .B(\us11\/_0070_ ), .X(\us11\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us11/_1022_ ( .A(\us11\/_0732_ ), .B(\us11\/_0123_ ), .C(\us11\/_0749_ ), .Y(\us11\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us11/_1023_ ( .A(\us11\/_0732_ ), .B(\us11\/_0467_ ), .C(\us11\/_0069_ ), .Y(\us11\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us11/_1024_ ( .A_N(\us11\/_0211_ ), .B(\us11\/_0127_ ), .C(\us11\/_0212_ ), .D(\us11\/_0213_ ), .X(\us11\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1025_ ( .A(\us11\/_0137_ ), .Y(\us11\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1026_ ( .A(\us11\/_0128_ ), .B(\us11\/_0035_ ), .Y(\us11\/_0217_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1028_ ( .A1(\us11\/_0159_ ), .A2(\us11\/_0746_ ), .B1(\us11\/_0434_ ), .B2(\us11\/_0499_ ), .Y(\us11\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us11/_1029_ ( .A1(\us11\/_0116_ ), .A2(\us11\/_0215_ ), .B1(\us11\/_0217_ ), .C1(\us11\/_0219_ ), .X(\us11\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1030_ ( .A(\us11\/_0113_ ), .B(\us11\/_0746_ ), .X(\us11\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us11/_1031_ ( .A1(\us11\/_0098_ ), .A2(\us11\/_0746_ ), .B1(\us11\/_0434_ ), .B2(\us11\/_0750_ ), .X(\us11\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1032_ ( .A1(\us11\/_0047_ ), .A2(\us11\/_0113_ ), .B1(\us11\/_0221_ ), .C1(\us11\/_0222_ ), .Y(\us11\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us11/_1033_ ( .A1(\us11\/_0129_ ), .A2(\us11\/_0162_ ), .B1(\us11\/_0271_ ), .B2(\us11\/_0705_ ), .X(\us11\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1034_ ( .A1(\us11\/_0093_ ), .A2(\us11\/_0738_ ), .B1(\us11\/_0081_ ), .C1(\us11\/_0224_ ), .Y(\us11\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1035_ ( .A(\us11\/_0214_ ), .B(\us11\/_0220_ ), .C(\us11\/_0223_ ), .D(\us11\/_0225_ ), .X(\us11\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1036_ ( .A(\us11\/_0196_ ), .B(\us11\/_0204_ ), .C(\us11\/_0210_ ), .D(\us11\/_0226_ ), .X(\us11\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1037_ ( .A(\us11\/_0111_ ), .B(\us11\/_0554_ ), .X(\us11\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1038_ ( .A(\us11\/_0229_ ), .Y(\us11\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1039_ ( .A(\us11\/_0111_ ), .B(\us11\/_0129_ ), .Y(\us11\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1040_ ( .A(\us11\/_0017_ ), .B(\us11\/_0738_ ), .Y(\us11\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1041_ ( .A(\us11\/_0030_ ), .B(\us11\/_0304_ ), .Y(\us11\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1042_ ( .A(\us11\/_0230_ ), .B(\us11\/_0231_ ), .C(\us11\/_0232_ ), .D(\us11\/_0233_ ), .X(\us11\/_0234_ ) );
sky130_fd_sc_hd__and2_1 \us11/_1043_ ( .A(\us11\/_0047_ ), .B(\us11\/_0478_ ), .X(\us11\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1044_ ( .A1(\us11\/_0129_ ), .A2(\us11\/_0554_ ), .B1(\us11\/_0137_ ), .Y(\us11\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us11/_1045_ ( .A(\us11\/_0235_ ), .B(\us11\/_0049_ ), .C_N(\us11\/_0236_ ), .Y(\us11\/_0237_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1046_ ( .A(\us11\/_0047_ ), .B(\us11\/_0077_ ), .X(\us11\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1047_ ( .A(\us11\/_0070_ ), .B(\us11\/_0035_ ), .X(\us11\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us11/_1048_ ( .A1(\us11\/_0047_ ), .A2(\us11\/_0736_ ), .B1(\us11\/_0022_ ), .B2(\us11\/_0364_ ), .X(\us11\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us11/_1049_ ( .A(\us11\/_0239_ ), .B(\us11\/_0240_ ), .C(\us11\/_0241_ ), .Y(\us11\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1050_ ( .A(\us11\/_0554_ ), .B(\us11\/_0072_ ), .X(\us11\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us11/_1051_ ( .A1(\us11\/_0142_ ), .A2(\us11\/_0137_ ), .B1(\us11\/_0159_ ), .B2(\us11\/_0082_ ), .X(\us11\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1052_ ( .A1(\us11\/_0608_ ), .A2(\us11\/_0072_ ), .B1(\us11\/_0243_ ), .C1(\us11\/_0244_ ), .Y(\us11\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1053_ ( .A(\us11\/_0234_ ), .B(\us11\/_0237_ ), .C(\us11\/_0242_ ), .D(\us11\/_0245_ ), .X(\us11\/_0246_ ) );
sky130_fd_sc_hd__buf_2 \us11/_1054_ ( .A(\us11\/_0027_ ), .X(\us11\/_0247_ ) );
sky130_fd_sc_hd__o21a_1 \us11/_1055_ ( .A1(\us11\/_0554_ ), .A2(\us11\/_0586_ ), .B1(\us11\/_0247_ ), .X(\us11\/_0248_ ) );
sky130_fd_sc_hd__and2_1 \us11/_1056_ ( .A(\us11\/_0082_ ), .B(\us11\/_0478_ ), .X(\us11\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_1057_ ( .A(\us11\/_0079_ ), .X(\us11\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1058_ ( .A(\us11\/_0251_ ), .B(\us11\/_0478_ ), .X(\us11\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_1059_ ( .A(\us11\/_0250_ ), .B(\us11\/_0252_ ), .Y(\us11\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1060_ ( .A(\us11\/_0016_ ), .B(\us11\/_0064_ ), .Y(\us11\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_1061_ ( .A(\us11\/_0304_ ), .X(\us11\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1062_ ( .A(\us11\/_0255_ ), .B(\us11\/_0640_ ), .Y(\us11\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us11/_1063_ ( .A_N(\us11\/_0248_ ), .B(\us11\/_0253_ ), .C(\us11\/_0254_ ), .D(\us11\/_0256_ ), .X(\us11\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1064_ ( .A(\us11\/_0364_ ), .B(\us11\/_0110_ ), .X(\us11\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us11/_1065_ ( .A1(\us11\/_0161_ ), .A2(\us11\/_0130_ ), .B1(\us11\/_0258_ ), .Y(\us11\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1066_ ( .A(\us11\/_0194_ ), .B(\sa11\[1\] ), .X(\us11\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1068_ ( .A(\us11\/_0261_ ), .B(\us11\/_0153_ ), .Y(\us11\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us11/_1069_ ( .A_N(\us11\/_0154_ ), .B(\us11\/_0259_ ), .C(\us11\/_0263_ ), .X(\us11\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1070_ ( .A(\us11\/_0246_ ), .B(\us11\/_0174_ ), .C(\us11\/_0257_ ), .D(\us11\/_0264_ ), .X(\us11\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us11/_1071_ ( .A1(\us11\/_0261_ ), .A2(\us11\/_0554_ ), .B1(\us11\/_0159_ ), .X(\us11\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1072_ ( .A(\us11\/_0746_ ), .B(\us11\/_0150_ ), .Y(\us11\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1073_ ( .A(\us11\/_0175_ ), .Y(\us11\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us11/_1074_ ( .A(\us11\/_0423_ ), .B(\us11\/_0123_ ), .C(\us11\/_0151_ ), .X(\us11\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1075_ ( .A(\us11\/_0268_ ), .B(\us11\/_0269_ ), .Y(\us11\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us11/_1076_ ( .A_N(\us11\/_0266_ ), .B(\us11\/_0267_ ), .C(\us11\/_0270_ ), .X(\us11\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1077_ ( .A(\us11\/_0554_ ), .B(\us11\/_0150_ ), .X(\us11\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1078_ ( .A(\us11\/_0273_ ), .Y(\us11\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1079_ ( .A1(\us11\/_0734_ ), .A2(\us11\/_0325_ ), .B1(\us11\/_0380_ ), .Y(\us11\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1080_ ( .A(\us11\/_0275_ ), .Y(\us11\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1081_ ( .A(\us11\/_0276_ ), .B(\us11\/_0153_ ), .Y(\us11\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us11/_1082_ ( .A(\us11\/_0272_ ), .B(\us11\/_0274_ ), .C(\us11\/_0277_ ), .X(\us11\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_1083_ ( .A(\us11\/_0035_ ), .X(\us11\/_0279_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1085_ ( .A1(\us11\/_0499_ ), .A2(\us11\/_0279_ ), .B1(\us11\/_0084_ ), .B2(\us11\/_0060_ ), .Y(\us11\/_0281_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1086_ ( .A1(\us11\/_0251_ ), .A2(\us11\/_0434_ ), .B1(\us11\/_0304_ ), .Y(\us11\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1087_ ( .A(\us11\/_0091_ ), .B(\us11\/_0292_ ), .Y(\us11\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1088_ ( .A1(\us11\/_0118_ ), .A2(\us11\/_0050_ ), .B1(\us11\/_0038_ ), .C1(\us11\/_0255_ ), .Y(\us11\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1089_ ( .A(\us11\/_0281_ ), .B(\us11\/_0283_ ), .C(\us11\/_0284_ ), .D(\us11\/_0285_ ), .X(\us11\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1090_ ( .A(\us11\/_0082_ ), .B(\us11\/_0027_ ), .X(\us11\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1091_ ( .A(\us11\/_0129_ ), .B(\us11\/_0027_ ), .X(\us11\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_1092_ ( .A(\us11\/_0287_ ), .B(\us11\/_0288_ ), .Y(\us11\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1093_ ( .A1(\us11\/_0752_ ), .A2(\us11\/_0683_ ), .B1(\us11\/_0093_ ), .B2(\us11\/_0247_ ), .Y(\us11\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1094_ ( .A1(\us11\/_0092_ ), .A2(\us11\/_0575_ ), .B1(\us11\/_0292_ ), .Y(\us11\/_0291_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_1095_ ( .A(\us11\/_0054_ ), .X(\us11\/_0292_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1096_ ( .A1(\us11\/_0499_ ), .A2(\us11\/_0662_ ), .B1(\us11\/_0084_ ), .B2(\us11\/_0292_ ), .Y(\us11\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1097_ ( .A(\us11\/_0289_ ), .B(\us11\/_0290_ ), .C(\us11\/_0291_ ), .D(\us11\/_0294_ ), .X(\us11\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1098_ ( .A(\us11\/_0750_ ), .B(\us11\/_0193_ ), .X(\us11\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1099_ ( .A(\us11\/_0705_ ), .B(\us11\/_0380_ ), .X(\us11\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1100_ ( .A(\us11\/_0752_ ), .B(\us11\/_0129_ ), .Y(\us11\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us11/_1101_ ( .A(\us11\/_0296_ ), .B(\us11\/_0297_ ), .C_N(\us11\/_0298_ ), .Y(\us11\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1102_ ( .A(\us11\/_0089_ ), .B(\us11\/_0532_ ), .Y(\us11\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1103_ ( .A(\sa11\[2\] ), .Y(\us11\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \us11/_1104_ ( .A(\us11\/_0301_ ), .B(\sa11\[3\] ), .C(\us11\/_0118_ ), .Y(\us11\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1105_ ( .A(\us11\/_0072_ ), .B(\us11\/_0302_ ), .X(\us11\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1106_ ( .A(\us11\/_0303_ ), .Y(\us11\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1107_ ( .A(\us11\/_0147_ ), .B(\us11\/_0302_ ), .Y(\us11\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1108_ ( .A(\us11\/_0299_ ), .B(\us11\/_0300_ ), .C(\us11\/_0305_ ), .D(\us11\/_0306_ ), .X(\us11\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1109_ ( .A(\us11\/_0278_ ), .B(\us11\/_0286_ ), .C(\us11\/_0295_ ), .D(\us11\/_0307_ ), .X(\us11\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us11/_1110_ ( .A(\us11\/_0228_ ), .B(\us11\/_0265_ ), .C(\us11\/_0308_ ), .Y(\us11\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1111_ ( .A(\us11\/_0235_ ), .Y(\us11\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1112_ ( .A(\us11\/_0478_ ), .B(\us11\/_0640_ ), .X(\us11\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1113_ ( .A(\us11\/_0310_ ), .Y(\us11\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1114_ ( .A(\us11\/_0022_ ), .B(\us11\/_0499_ ), .Y(\us11\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1115_ ( .A(\us11\/_0499_ ), .B(\us11\/_0032_ ), .Y(\us11\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1116_ ( .A(\us11\/_0309_ ), .B(\us11\/_0311_ ), .C(\us11\/_0312_ ), .D(\us11\/_0313_ ), .X(\us11\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1117_ ( .A(\us11\/_0499_ ), .B(\us11\/_0064_ ), .Y(\us11\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1118_ ( .A(\us11\/_0499_ ), .B(\us11\/_0683_ ), .Y(\us11\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1119_ ( .A(\us11\/_0315_ ), .B(\us11\/_0316_ ), .C(\us11\/_0317_ ), .D(\us11\/_0253_ ), .X(\us11\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1120_ ( .A(\us11\/_0047_ ), .B(\us11\/_0304_ ), .Y(\us11\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1121_ ( .A(\us11\/_0586_ ), .B(\us11\/_0162_ ), .Y(\us11\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1122_ ( .A(\us11\/_0319_ ), .B(\us11\/_0320_ ), .Y(\us11\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_1123_ ( .A(\us11\/_0321_ ), .B(\us11\/_0238_ ), .Y(\us11\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1124_ ( .A(\us11\/_0304_ ), .B(\us11\/_0062_ ), .Y(\us11\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_1125_ ( .A(\us11\/_0251_ ), .X(\us11\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1126_ ( .A1(\us11\/_0324_ ), .A2(\us11\/_0084_ ), .B1(\us11\/_0255_ ), .Y(\us11\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1127_ ( .A1(\us11\/_0050_ ), .A2(\us11\/_0216_ ), .B1(\us11\/_0109_ ), .C1(\us11\/_0255_ ), .Y(\us11\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1128_ ( .A(\us11\/_0322_ ), .B(\us11\/_0323_ ), .C(\us11\/_0326_ ), .D(\us11\/_0327_ ), .X(\us11\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1129_ ( .A1(\us11\/_0733_ ), .A2(\us11\/_0279_ ), .A3(\us11\/_0058_ ), .B1(\us11\/_0292_ ), .Y(\us11\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_1130_ ( .A(\us11\/_0047_ ), .X(\us11\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1131_ ( .A(\us11\/_0330_ ), .B(\us11\/_0292_ ), .Y(\us11\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1132_ ( .A(\us11\/_0054_ ), .B(\us11\/_0045_ ), .Y(\us11\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1133_ ( .A(\us11\/_0329_ ), .B(\us11\/_0331_ ), .C(\us11\/_0284_ ), .D(\us11\/_0332_ ), .X(\us11\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us11/_1134_ ( .A1(\us11\/_0543_ ), .A2(\us11\/_0216_ ), .B1(\us11\/_0532_ ), .C1(\us11\/_0060_ ), .X(\us11\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1135_ ( .A(\us11\/_0084_ ), .B(\us11\/_0060_ ), .Y(\us11\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1136_ ( .A(\us11\/_0324_ ), .B(\us11\/_0060_ ), .Y(\us11\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1137_ ( .A(\us11\/_0335_ ), .B(\us11\/_0337_ ), .Y(\us11\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1138_ ( .A1(\us11\/_0276_ ), .A2(\us11\/_0060_ ), .B1(\us11\/_0334_ ), .C1(\us11\/_0338_ ), .Y(\us11\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1139_ ( .A(\us11\/_0318_ ), .B(\us11\/_0328_ ), .C(\us11\/_0333_ ), .D(\us11\/_0339_ ), .X(\us11\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us11/_1140_ ( .A1(\us11\/_0746_ ), .A2(\us11\/_0134_ ), .B1(\us11\/_0128_ ), .X(\us11\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us11/_1141_ ( .A_N(\us11\/_0086_ ), .B(\us11\/_0128_ ), .X(\us11\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1142_ ( .A(\us11\/_0079_ ), .B(\us11\/_0124_ ), .X(\us11\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_1143_ ( .A(\us11\/_0126_ ), .B(\us11\/_0343_ ), .Y(\us11\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us11/_1144_ ( .A(\us11\/_0341_ ), .B(\us11\/_0342_ ), .C_N(\us11\/_0344_ ), .Y(\us11\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1146_ ( .A1(\us11\/_0193_ ), .A2(\us11\/_0092_ ), .A3(\us11\/_0330_ ), .B1(\us11\/_0147_ ), .Y(\us11\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1147_ ( .A1(\us11\/_0130_ ), .A2(\us11\/_0084_ ), .A3(\us11\/_0134_ ), .B1(\us11\/_0139_ ), .Y(\us11\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1148_ ( .A1(\us11\/_0144_ ), .A2(\us11\/_0608_ ), .A3(\us11\/_0092_ ), .B1(\us11\/_0139_ ), .Y(\us11\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1149_ ( .A(\us11\/_0345_ ), .B(\us11\/_0348_ ), .C(\us11\/_0349_ ), .D(\us11\/_0350_ ), .X(\us11\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us11/_1150_ ( .A(\us11\/_0150_ ), .B(\us11\/_0194_ ), .C(\us11\/_0543_ ), .X(\us11\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us11/_1151_ ( .A(\us11\/_0277_ ), .SLEEP(\us11\/_0352_ ), .X(\us11\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us11/_1152_ ( .A1(\us11\/_0268_ ), .A2(\us11\/_0171_ ), .B1(\us11\/_0157_ ), .Y(\us11\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us11/_1153_ ( .A(\us11\/_0161_ ), .X(\us11\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1154_ ( .A1(\us11\/_0279_ ), .A2(\us11\/_0084_ ), .B1(\us11\/_0355_ ), .Y(\us11\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1155_ ( .A1(\us11\/_0020_ ), .A2(\us11\/_0193_ ), .A3(\us11\/_0091_ ), .B1(\us11\/_0355_ ), .Y(\us11\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1156_ ( .A(\us11\/_0353_ ), .B(\us11\/_0354_ ), .C(\us11\/_0356_ ), .D(\us11\/_0357_ ), .X(\us11\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1157_ ( .A(\us11\/_0111_ ), .B(\us11\/_0586_ ), .X(\us11\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1158_ ( .A(\us11\/_0360_ ), .Y(\us11\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us11/_1159_ ( .A1(\us11\/_0119_ ), .A2(\us11\/_0120_ ), .B1(\us11\/_0230_ ), .C1(\us11\/_0361_ ), .X(\us11\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1160_ ( .A1(\us11\/_0662_ ), .A2(\us11\/_0251_ ), .A3(\us11\/_0134_ ), .B1(\us11\/_0114_ ), .Y(\us11\/_0363_ ) );
sky130_fd_sc_hd__buf_2 \us11/_1161_ ( .A(\us11\/_0098_ ), .X(\us11\/_0364_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1162_ ( .A1(\us11\/_0035_ ), .A2(\us11\/_0251_ ), .A3(\us11\/_0134_ ), .B1(\us11\/_0364_ ), .Y(\us11\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1163_ ( .A1(\us11\/_0193_ ), .A2(\us11\/_0608_ ), .B1(\us11\/_0364_ ), .Y(\us11\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1164_ ( .A(\us11\/_0362_ ), .B(\us11\/_0363_ ), .C(\us11\/_0365_ ), .D(\us11\/_0366_ ), .X(\us11\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1165_ ( .A1(\us11\/_0575_ ), .A2(\us11\/_0092_ ), .A3(\us11\/_0330_ ), .B1(\us11\/_0089_ ), .Y(\us11\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1166_ ( .A1(\us11\/_0586_ ), .A2(\us11\/_0017_ ), .A3(\us11\/_0330_ ), .B1(\us11\/_0094_ ), .Y(\us11\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \us11/_1167_ ( .A1(\us11\/_0293_ ), .A2(\us11\/_0134_ ), .B1(\us11\/_0089_ ), .Y(\us11\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1168_ ( .A1(\us11\/_0279_ ), .A2(\us11\/_0134_ ), .B1(\us11\/_0094_ ), .Y(\us11\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1169_ ( .A(\us11\/_0368_ ), .B(\us11\/_0370_ ), .C(\us11\/_0371_ ), .D(\us11\/_0372_ ), .X(\us11\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1170_ ( .A(\us11\/_0351_ ), .B(\us11\/_0359_ ), .C(\us11\/_0367_ ), .D(\us11\/_0373_ ), .X(\us11\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1171_ ( .A1(\us11\/_0102_ ), .A2(\us11\/_0347_ ), .B1(\us11\/_0109_ ), .C1(\us11\/_0247_ ), .Y(\us11\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1172_ ( .A1(\us11\/_0102_ ), .A2(\us11\/_0347_ ), .B1(\us11\/_0532_ ), .C1(\us11\/_0247_ ), .Y(\us11\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1173_ ( .A1(\us11\/_0050_ ), .A2(\us11\/_0543_ ), .B1(\us11\/_0380_ ), .C1(\us11\/_0247_ ), .Y(\us11\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1174_ ( .A(\us11\/_0041_ ), .B(\us11\/_0375_ ), .C(\us11\/_0376_ ), .D(\us11\/_0377_ ), .X(\us11\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1175_ ( .A(\us11\/_0047_ ), .B(\us11\/_0750_ ), .X(\us11\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1176_ ( .A(\us11\/_0379_ ), .Y(\us11\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1177_ ( .A(\us11\/_0016_ ), .B(\us11\/_0608_ ), .Y(\us11\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1178_ ( .A(\us11\/_0752_ ), .B(\us11\/_0554_ ), .Y(\us11\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1179_ ( .A1(\sa11\[1\] ), .A2(\us11\/_0734_ ), .B1(\us11\/_0109_ ), .C1(\us11\/_0016_ ), .Y(\us11\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1180_ ( .A(\us11\/_0381_ ), .B(\us11\/_0382_ ), .C(\us11\/_0383_ ), .D(\us11\/_0384_ ), .X(\us11\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us11/_1181_ ( .A(\us11\/_0086_ ), .B_N(\us11\/_0736_ ), .X(\us11\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1182_ ( .A1(\us11\/_0748_ ), .A2(\us11\/_0134_ ), .B1(\us11\/_0739_ ), .Y(\us11\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1183_ ( .A1(\us11\/_0118_ ), .A2(\us11\/_0543_ ), .B1(\us11\/_0109_ ), .C1(\us11\/_0739_ ), .Y(\us11\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1184_ ( .A1(\us11\/_0102_ ), .A2(\us11\/_0301_ ), .B1(\sa11\[3\] ), .C1(\us11\/_0739_ ), .Y(\us11\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1185_ ( .A(\us11\/_0386_ ), .B(\us11\/_0387_ ), .C(\us11\/_0388_ ), .D(\us11\/_0389_ ), .X(\us11\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1186_ ( .A(\us11\/_0020_ ), .Y(\us11\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1187_ ( .A(\us11\/_0727_ ), .Y(\us11\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1188_ ( .A(\us11\/_0727_ ), .B(\us11\/_0064_ ), .Y(\us11\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1189_ ( .A1(\us11\/_0102_ ), .A2(\us11\/_0734_ ), .B1(\us11\/_0532_ ), .C1(\us11\/_0727_ ), .Y(\us11\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us11/_1190_ ( .A1(\us11\/_0392_ ), .A2(\us11\/_0393_ ), .B1(\us11\/_0394_ ), .C1(\us11\/_0395_ ), .X(\us11\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1191_ ( .A(\us11\/_0378_ ), .B(\us11\/_0385_ ), .C(\us11\/_0390_ ), .D(\us11\/_0396_ ), .X(\us11\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us11/_1192_ ( .A(\us11\/_0340_ ), .B(\us11\/_0374_ ), .C(\us11\/_0397_ ), .Y(\us11\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1193_ ( .A(\us11\/_0077_ ), .B(\us11\/_0129_ ), .X(\us11\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_1194_ ( .A(\us11\/_0398_ ), .B(\us11\/_0239_ ), .Y(\us11\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1195_ ( .A(\us11\/_0022_ ), .B(\us11\/_0111_ ), .X(\us11\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us11/_1196_ ( .A_N(\us11\/_0400_ ), .B(\us11\/_0231_ ), .Y(\us11\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us11/_1197_ ( .A(\us11\/_0399_ ), .SLEEP(\us11\/_0402_ ), .X(\us11\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_1198_ ( .A(\us11\/_0746_ ), .B(\us11\/_0251_ ), .Y(\us11\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us11/_1199_ ( .A_N(\us11\/_0404_ ), .B(\us11\/_0752_ ), .Y(\us11\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us11/_1200_ ( .A(\us11\/_0467_ ), .B(\us11\/_0194_ ), .C(\us11\/_0694_ ), .X(\us11\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us11/_1201_ ( .A_N(\us11\/_0175_ ), .B(\us11\/_0406_ ), .X(\us11\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1202_ ( .A(\us11\/_0407_ ), .Y(\us11\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1203_ ( .A1(\us11\/_0094_ ), .A2(\us11\/_0197_ ), .B1(\us11\/_0114_ ), .B2(\us11\/_0640_ ), .Y(\us11\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1204_ ( .A(\us11\/_0403_ ), .B(\us11\/_0405_ ), .C(\us11\/_0408_ ), .D(\us11\/_0409_ ), .X(\us11\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1205_ ( .A(\us11\/_0030_ ), .B(\us11\/_0150_ ), .Y(\us11\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us11/_1206_ ( .A_N(\us11\/_0169_ ), .B(\us11\/_0289_ ), .C(\us11\/_0411_ ), .X(\us11\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us11/_1207_ ( .A1(\us11\/_0467_ ), .A2(\us11\/_0151_ ), .B1(\us11\/_0140_ ), .C1(\us11\/_0129_ ), .X(\us11\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1208_ ( .A1(\us11\/_0608_ ), .A2(\us11\/_0364_ ), .B1(\us11\/_0037_ ), .C1(\us11\/_0414_ ), .Y(\us11\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1209_ ( .A(\us11\/_0738_ ), .Y(\us11\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1210_ ( .A(\us11\/_0586_ ), .B(\us11\/_0736_ ), .Y(\us11\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1211_ ( .A1(\us11\/_0194_ ), .A2(\us11\/_0038_ ), .B1(\us11\/_0118_ ), .C1(\us11\/_0153_ ), .Y(\us11\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us11/_1212_ ( .A1(\us11\/_0416_ ), .A2(\us11\/_0117_ ), .B1(\us11\/_0417_ ), .C1(\us11\/_0418_ ), .X(\us11\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1213_ ( .A(\us11\/_0077_ ), .B(\us11\/_0035_ ), .X(\us11\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1214_ ( .A(\us11\/_0662_ ), .B(\us11\/_0124_ ), .Y(\us11\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1215_ ( .A(\us11\/_0030_ ), .B(\us11\/_0137_ ), .Y(\us11\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1216_ ( .A(\us11\/_0072_ ), .B(\us11\/_0732_ ), .Y(\us11\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us11/_1217_ ( .A_N(\us11\/_0420_ ), .B(\us11\/_0421_ ), .C(\us11\/_0422_ ), .D(\us11\/_0424_ ), .X(\us11\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1218_ ( .A(\us11\/_0413_ ), .B(\us11\/_0415_ ), .C(\us11\/_0419_ ), .D(\us11\/_0425_ ), .X(\us11\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us11/_1219_ ( .A(\us11\/_0355_ ), .B(\us11\/_0102_ ), .C(\us11\/_0109_ ), .Y(\us11\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1220_ ( .A(\us11\/_0077_ ), .B(\us11\/_0017_ ), .X(\us11\/_0428_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1221_ ( .A(\us11\/_0077_ ), .B(\us11\/_0554_ ), .X(\us11\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us11/_1222_ ( .A1(\us11\/_0050_ ), .A2(\us11\/_0216_ ), .B1(\us11\/_0380_ ), .C1(\us11\/_0078_ ), .X(\us11\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us11/_1223_ ( .A(\us11\/_0428_ ), .B(\us11\/_0429_ ), .C(\us11\/_0430_ ), .Y(\us11\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us11/_1224_ ( .A_N(\us11\/_0209_ ), .B(\us11\/_0431_ ), .X(\us11\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us11/_1225_ ( .A1(\us11\/_0215_ ), .A2(\us11\/_0404_ ), .B1(\us11\/_0427_ ), .C1(\us11\/_0432_ ), .X(\us11\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1226_ ( .A(\us11\/_0043_ ), .B(\us11\/_0058_ ), .Y(\us11\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1227_ ( .A(\us11\/_0195_ ), .B(\us11\/_0233_ ), .C(\us11\/_0320_ ), .D(\us11\/_0435_ ), .X(\us11\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1228_ ( .A(\us11\/_0261_ ), .B(\us11\/_0738_ ), .Y(\us11\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1229_ ( .A1(\us11\/_0499_ ), .A2(\us11\/_0640_ ), .B1(\us11\/_0261_ ), .B2(\us11\/_0292_ ), .Y(\us11\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1230_ ( .A(\us11\/_0436_ ), .B(\us11\/_0394_ ), .C(\us11\/_0437_ ), .D(\us11\/_0438_ ), .X(\us11\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1231_ ( .A(\us11\/_0410_ ), .B(\us11\/_0426_ ), .C(\us11\/_0433_ ), .D(\us11\/_0439_ ), .X(\us11\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us11/_1232_ ( .A(\us11\/_0135_ ), .SLEEP(\us11\/_0273_ ), .X(\us11\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1233_ ( .A1(\us11\/_0279_ ), .A2(\us11\/_0134_ ), .B1(\us11\/_0364_ ), .Y(\us11\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1234_ ( .A(\us11\/_0441_ ), .B(\us11\/_0164_ ), .C(\us11\/_0270_ ), .D(\us11\/_0442_ ), .X(\us11\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1235_ ( .A(\us11\/_0051_ ), .B(\us11\/_0662_ ), .Y(\us11\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1236_ ( .A(\us11\/_0051_ ), .B(\us11\/_0271_ ), .Y(\us11\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1237_ ( .A(\us11\/_0444_ ), .B(\us11\/_0446_ ), .X(\us11\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1238_ ( .A(\us11\/_0193_ ), .B(\us11\/_0304_ ), .X(\us11\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1239_ ( .A(\us11\/_0448_ ), .Y(\us11\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1240_ ( .A(\us11\/_0162_ ), .B(\us11\/_0130_ ), .X(\us11\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1241_ ( .A(\us11\/_0450_ ), .Y(\us11\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1242_ ( .A1(\us11\/_0129_ ), .A2(\us11\/_0554_ ), .B1(\us11\/_0043_ ), .Y(\us11\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1243_ ( .A(\us11\/_0447_ ), .B(\us11\/_0449_ ), .C(\us11\/_0451_ ), .D(\us11\/_0452_ ), .X(\us11\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1244_ ( .A(\us11\/_0292_ ), .B(\us11\/_0064_ ), .Y(\us11\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us11/_1245_ ( .A_N(\us11\/_0248_ ), .B(\us11\/_0454_ ), .C(\us11\/_0254_ ), .D(\us11\/_0256_ ), .X(\us11\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1246_ ( .A1(\us11\/_0330_ ), .A2(\us11\/_0364_ ), .B1(\us11\/_0134_ ), .B2(\us11\/_0705_ ), .Y(\us11\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1247_ ( .A1(\us11\/_0748_ ), .A2(\us11\/_0738_ ), .B1(\us11\/_0092_ ), .B2(\us11\/_0752_ ), .Y(\us11\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1248_ ( .A1(\us11\/_0072_ ), .A2(\us11\/_0035_ ), .B1(\us11\/_0748_ ), .B2(\us11\/_0292_ ), .Y(\us11\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1249_ ( .A1(\us11\/_0748_ ), .A2(\us11\/_0251_ ), .B1(\us11\/_0247_ ), .Y(\us11\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1250_ ( .A(\us11\/_0457_ ), .B(\us11\/_0458_ ), .C(\us11\/_0459_ ), .D(\us11\/_0460_ ), .X(\us11\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1251_ ( .A(\us11\/_0443_ ), .B(\us11\/_0453_ ), .C(\us11\/_0455_ ), .D(\us11\/_0461_ ), .X(\us11\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1252_ ( .A(\us11\/_0705_ ), .B(\us11\/_0079_ ), .X(\us11\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1253_ ( .A(\us11\/_0586_ ), .B(\us11\/_0124_ ), .Y(\us11\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1254_ ( .A(\us11\/_0499_ ), .B(\us11\/_0746_ ), .Y(\us11\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us11/_1255_ ( .A_N(\us11\/_0463_ ), .B(\us11\/_0464_ ), .C(\us11\/_0465_ ), .X(\us11\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us11/_1256_ ( .A1(\us11\/_0271_ ), .A2(\us11\/_0072_ ), .B1(\us11\/_0142_ ), .B2(\us11\/_0027_ ), .X(\us11\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1257_ ( .A1(\us11\/_0144_ ), .A2(\us11\/_0364_ ), .B1(\us11\/_0360_ ), .C1(\us11\/_0468_ ), .Y(\us11\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us11/_1258_ ( .A1(\us11\/_0662_ ), .A2(\us11\/_0251_ ), .B1(\us11\/_0499_ ), .X(\us11\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1259_ ( .A1(\us11\/_0575_ ), .A2(\us11\/_0292_ ), .B1(\us11\/_0379_ ), .C1(\us11\/_0470_ ), .Y(\us11\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1260_ ( .A(\us11\/_0466_ ), .B(\us11\/_0469_ ), .C(\us11\/_0471_ ), .D(\us11\/_0305_ ), .X(\us11\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us11/_1261_ ( .A1(\us11\/_0247_ ), .A2(\us11\/_0683_ ), .B1(\us11\/_0324_ ), .B2(\us11\/_0292_ ), .X(\us11\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1262_ ( .A(\us11\/_0084_ ), .B(\us11\/_0364_ ), .X(\us11\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us11/_1263_ ( .A1(\us11\/_0092_ ), .A2(\us11\/_0247_ ), .B1(\us11\/_0474_ ), .X(\us11\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us11/_1264_ ( .A(\us11\/_0075_ ), .B(\us11\/_0473_ ), .C(\us11\/_0475_ ), .Y(\us11\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1265_ ( .A1(\us11\/_0279_ ), .A2(\us11\/_0255_ ), .B1(\us11\/_0084_ ), .B2(\us11\/_0060_ ), .Y(\us11\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1266_ ( .A1(\us11\/_0093_ ), .A2(\us11\/_0292_ ), .B1(\us11\/_0134_ ), .B2(\us11\/_0114_ ), .Y(\us11\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1267_ ( .A1(\us11\/_0161_ ), .A2(\us11\/_0032_ ), .B1(\us11\/_0324_ ), .B2(\us11\/_0147_ ), .Y(\us11\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1268_ ( .A1(\us11\/_0054_ ), .A2(\us11\/_0732_ ), .B1(\us11\/_0748_ ), .B2(\us11\/_0304_ ), .Y(\us11\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1269_ ( .A(\us11\/_0477_ ), .B(\us11\/_0479_ ), .C(\us11\/_0480_ ), .D(\us11\/_0481_ ), .X(\us11\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1270_ ( .A(\us11\/_0161_ ), .B(\us11\/_0064_ ), .Y(\us11\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us11/_1271_ ( .A(\us11\/_0732_ ), .B(\us11\/_0123_ ), .C(\us11\/_0467_ ), .Y(\us11\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1272_ ( .A(\us11\/_0483_ ), .B(\us11\/_0484_ ), .Y(\us11\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1273_ ( .A(\us11\/_0297_ ), .Y(\us11\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us11/_1274_ ( .A_N(\us11\/_0485_ ), .B(\us11\/_0181_ ), .C(\us11\/_0486_ ), .D(\us11\/_0386_ ), .X(\us11\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1275_ ( .A(\us11\/_0472_ ), .B(\us11\/_0476_ ), .C(\us11\/_0482_ ), .D(\us11\/_0487_ ), .X(\us11\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \us11/_1276_ ( .A(\us11\/_0440_ ), .B(\us11\/_0462_ ), .C(\us11\/_0488_ ), .Y(\us11\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1277_ ( .A(\us11\/_0403_ ), .B(\us11\/_0230_ ), .C(\us11\/_0451_ ), .D(\us11\/_0361_ ), .X(\us11\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1278_ ( .A1(\us11\/_0118_ ), .A2(\us11\/_0050_ ), .B1(\us11\/_0109_ ), .C1(\us11\/_0139_ ), .Y(\us11\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1279_ ( .A(\us11\/_0447_ ), .B(\us11\/_0437_ ), .C(\us11\/_0491_ ), .D(\us11\/_0427_ ), .X(\us11\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1280_ ( .A1(\us11\/_0084_ ), .A2(\us11\/_0255_ ), .B1(\us11\/_0608_ ), .B2(\us11\/_0247_ ), .Y(\us11\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1281_ ( .A1(\us11\/_0144_ ), .A2(\us11\/_0147_ ), .B1(\us11\/_0355_ ), .B2(\us11\/_0093_ ), .Y(\us11\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1282_ ( .A1(\us11\/_0705_ ), .A2(\us11\/_0279_ ), .B1(\us11\/_0330_ ), .B2(\us11\/_0247_ ), .Y(\us11\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1283_ ( .A1(\us11\/_0279_ ), .A2(\us11\/_0084_ ), .B1(\us11\/_0114_ ), .Y(\us11\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1284_ ( .A(\us11\/_0493_ ), .B(\us11\/_0494_ ), .C(\us11\/_0495_ ), .D(\us11\/_0496_ ), .X(\us11\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1285_ ( .A1(\us11\/_0134_ ), .A2(\us11\/_0137_ ), .B1(\us11\/_0355_ ), .B2(\us11\/_0575_ ), .Y(\us11\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1286_ ( .A1(\us11\/_0364_ ), .A2(\us11\/_0733_ ), .B1(\us11\/_0093_ ), .B2(\us11\/_0499_ ), .Y(\us11\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1287_ ( .A(\us11\/_0147_ ), .B(\us11\/_0640_ ), .Y(\us11\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1288_ ( .A1(\us11\/_0153_ ), .A2(\us11\/_0292_ ), .B1(\us11\/_0748_ ), .Y(\us11\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1289_ ( .A(\us11\/_0498_ ), .B(\us11\/_0500_ ), .C(\us11\/_0501_ ), .D(\us11\/_0502_ ), .X(\us11\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1290_ ( .A(\us11\/_0490_ ), .B(\us11\/_0492_ ), .C(\us11\/_0497_ ), .D(\us11\/_0503_ ), .X(\us11\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us11/_1291_ ( .A_N(\us11\/_0275_ ), .B(\us11\/_0705_ ), .X(\us11\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1292_ ( .A(\us11\/_0505_ ), .Y(\us11\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1293_ ( .A(\us11\/_0380_ ), .B(\us11\/_0347_ ), .X(\us11\/_0507_ ) );
sky130_fd_sc_hd__o21ai_1 \us11/_1294_ ( .A1(\us11\/_0507_ ), .A2(\us11\/_0093_ ), .B1(\us11\/_0292_ ), .Y(\us11\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1295_ ( .A(\us11\/_0322_ ), .B(\us11\/_0277_ ), .C(\us11\/_0506_ ), .D(\us11\/_0508_ ), .X(\us11\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1296_ ( .A(\us11\/_0084_ ), .B(\us11\/_0705_ ), .X(\us11\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1297_ ( .A1(\us11\/_0733_ ), .A2(\us11\/_0114_ ), .B1(\us11\/_0429_ ), .C1(\us11\/_0511_ ), .Y(\us11\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_1298_ ( .A(\us11\/_0019_ ), .B(\us11\/_0024_ ), .Y(\us11\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1299_ ( .A(\us11\/_0512_ ), .B(\us11\/_0513_ ), .C(\us11\/_0742_ ), .D(\us11\/_0306_ ), .X(\us11\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1300_ ( .A1(\us11\/_0532_ ), .A2(\us11\/_0089_ ), .B1(\us11\/_0154_ ), .C1(\us11\/_0169_ ), .Y(\us11\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us11/_1301_ ( .A1(\us11\/_0749_ ), .A2(\us11\/_0026_ ), .B1(\us11\/_0069_ ), .C1(\us11\/_0032_ ), .X(\us11\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us11/_1302_ ( .A1(\us11\/_0324_ ), .A2(\us11\/_0355_ ), .B1(\us11\/_0330_ ), .B2(\us11\/_0727_ ), .X(\us11\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us11/_1303_ ( .A(\us11\/_0133_ ), .B(\us11\/_0516_ ), .C(\us11\/_0517_ ), .Y(\us11\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1304_ ( .A(\us11\/_0509_ ), .B(\us11\/_0514_ ), .C(\us11\/_0515_ ), .D(\us11\/_0518_ ), .X(\us11\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1305_ ( .A(\us11\/_0746_ ), .B(\us11\/_0072_ ), .Y(\us11\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1306_ ( .A1(\us11\/_0082_ ), .A2(\us11\/_0070_ ), .B1(\us11\/_0043_ ), .B2(\us11\/_0193_ ), .Y(\us11\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1307_ ( .A(\us11\/_0311_ ), .B(\us11\/_0520_ ), .C(\us11\/_0332_ ), .D(\us11\/_0522_ ), .X(\us11\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1308_ ( .A(\us11\/_0129_ ), .B(\us11\/_0499_ ), .X(\us11\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_1309_ ( .A(\us11\/_0235_ ), .B(\us11\/_0524_ ), .Y(\us11\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us11/_1310_ ( .A(\us11\/_0081_ ), .B(\us11\/_0085_ ), .Y(\us11\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1311_ ( .A1(\us11\/_0051_ ), .A2(\us11\/_0045_ ), .B1(\us11\/_0130_ ), .B2(\us11\/_0094_ ), .Y(\us11\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1312_ ( .A(\us11\/_0523_ ), .B(\us11\/_0525_ ), .C(\us11\/_0526_ ), .D(\us11\/_0527_ ), .X(\us11\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us11/_1313_ ( .A_N(\us11\/_0250_ ), .B(\us11\/_0521_ ), .Y(\us11\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1314_ ( .A(\us11\/_0128_ ), .B(\us11\/_0020_ ), .X(\us11\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1315_ ( .A(\us11\/_0530_ ), .Y(\us11\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1316_ ( .A(\us11\/_0364_ ), .B(\us11\/_0058_ ), .X(\us11\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1317_ ( .A(\us11\/_0533_ ), .Y(\us11\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us11/_1318_ ( .A_N(\us11\/_0529_ ), .B(\us11\/_0531_ ), .C(\us11\/_0534_ ), .D(\us11\/_0192_ ), .X(\us11\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1319_ ( .A(\us11\/_0434_ ), .B(\us11\/_0078_ ), .X(\us11\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us11/_1320_ ( .A1(\us11\/_0750_ ), .A2(\us11\/_0079_ ), .B1(\us11\/_0129_ ), .B2(\us11\/_0705_ ), .X(\us11\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1321_ ( .A1(\us11\/_0161_ ), .A2(\us11\/_0032_ ), .B1(\us11\/_0536_ ), .C1(\us11\/_0537_ ), .Y(\us11\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us11/_1322_ ( .A1(\us11\/_0746_ ), .A2(\us11\/_0162_ ), .B1(\us11\/_0079_ ), .B2(\us11\/_0043_ ), .X(\us11\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1323_ ( .A1(\us11\/_0093_ ), .A2(\us11\/_0247_ ), .B1(\us11\/_0240_ ), .C1(\us11\/_0539_ ), .Y(\us11\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1324_ ( .A(\us11\/_0434_ ), .B(\us11\/_0043_ ), .X(\us11\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us11/_1325_ ( .A1(\us11\/_0142_ ), .A2(\us11\/_0150_ ), .B1(\us11\/_0022_ ), .B2(\us11\/_0137_ ), .X(\us11\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1326_ ( .A1(\us11\/_0279_ ), .A2(\us11\/_0051_ ), .B1(\us11\/_0541_ ), .C1(\us11\/_0542_ ), .Y(\us11\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1327_ ( .A(\us11\/_0159_ ), .B(\us11\/_0035_ ), .X(\us11\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us11/_1328_ ( .A1(\us11\/_0271_ ), .A2(\us11\/_0434_ ), .B1(\us11\/_0027_ ), .X(\us11\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1329_ ( .A1(\us11\/_0091_ ), .A2(\us11\/_0128_ ), .B1(\us11\/_0545_ ), .C1(\us11\/_0546_ ), .Y(\us11\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1330_ ( .A(\us11\/_0538_ ), .B(\us11\/_0540_ ), .C(\us11\/_0544_ ), .D(\us11\/_0547_ ), .X(\us11\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1331_ ( .A(\us11\/_0364_ ), .B(\us11\/_0193_ ), .X(\us11\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us11/_1332_ ( .A(\us11\/_0549_ ), .B(\us11\/_0186_ ), .C(\us11\/_0187_ ), .Y(\us11\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1333_ ( .A(\us11\/_0062_ ), .B(\us11\/_0347_ ), .C(\us11\/_0749_ ), .D(\us11\/_0694_ ), .X(\us11\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1334_ ( .A1(\us11\/_0130_ ), .A2(\us11\/_0499_ ), .B1(\us11\/_0551_ ), .C1(\us11\/_0101_ ), .Y(\us11\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1335_ ( .A(\us11\/_0139_ ), .B(\us11\/_0640_ ), .Y(\us11\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1336_ ( .A1(\us11\/_0752_ ), .A2(\us11\/_0662_ ), .B1(\us11\/_0084_ ), .B2(\us11\/_0364_ ), .Y(\us11\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1337_ ( .A(\us11\/_0550_ ), .B(\us11\/_0552_ ), .C(\us11\/_0553_ ), .D(\us11\/_0555_ ), .X(\us11\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1338_ ( .A(\us11\/_0528_ ), .B(\us11\/_0535_ ), .C(\us11\/_0548_ ), .D(\us11\/_0556_ ), .X(\us11\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us11/_1339_ ( .A(\us11\/_0504_ ), .B(\us11\/_0519_ ), .C(\us11\/_0557_ ), .Y(\us11\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1340_ ( .A(\us11\/_0054_ ), .B(\us11\/_0507_ ), .X(\us11\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us11/_1341_ ( .A_N(\us11\/_0558_ ), .B(\us11\/_0408_ ), .C(\us11\/_0451_ ), .D(\us11\/_0452_ ), .X(\us11\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1342_ ( .A(\us11\/_0549_ ), .Y(\us11\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1343_ ( .A(\us11\/_0559_ ), .B(\us11\/_0403_ ), .C(\us11\/_0560_ ), .D(\us11\/_0371_ ), .X(\us11\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1344_ ( .A(\us11\/_0181_ ), .B(\us11\/_0178_ ), .X(\us11\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1345_ ( .A(\us11\/_0562_ ), .B(\us11\/_0552_ ), .C(\us11\/_0553_ ), .D(\us11\/_0555_ ), .X(\us11\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1346_ ( .A(\us11\/_0247_ ), .B(\us11\/_0020_ ), .Y(\us11\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1347_ ( .A(\us11\/_0051_ ), .B(\us11\/_0130_ ), .X(\us11\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1348_ ( .A(\us11\/_0566_ ), .Y(\us11\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1349_ ( .A(\us11\/_0159_ ), .B(\us11\/_0423_ ), .X(\us11\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1350_ ( .A1(\us11\/_0752_ ), .A2(\us11\/_0640_ ), .B1(\us11\/_0568_ ), .B2(\us11\/_0175_ ), .Y(\us11\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1351_ ( .A(\us11\/_0076_ ), .B(\us11\/_0565_ ), .C(\us11\/_0567_ ), .D(\us11\/_0569_ ), .X(\us11\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us11/_1352_ ( .A1(\us11\/_0035_ ), .A2(\us11\/_0142_ ), .B1(\us11\/_0161_ ), .X(\us11\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1353_ ( .A(\us11\/_0364_ ), .B(\us11\/_0662_ ), .Y(\us11\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us11/_1354_ ( .A(\us11\/_0420_ ), .B(\us11\/_0571_ ), .C_N(\us11\/_0572_ ), .Y(\us11\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1355_ ( .A(\us11\/_0051_ ), .B(\us11\/_0746_ ), .Y(\us11\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1356_ ( .A(\us11\/_0574_ ), .B(\us11\/_0319_ ), .C(\us11\/_0320_ ), .D(\us11\/_0411_ ), .X(\us11\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1357_ ( .A(\us11\/_0736_ ), .B(\us11\/_0035_ ), .Y(\us11\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1358_ ( .A(\us11\/_0736_ ), .B(\us11\/_0030_ ), .Y(\us11\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1359_ ( .A(\us11\/_0298_ ), .B(\us11\/_0208_ ), .C(\us11\/_0577_ ), .D(\us11\/_0578_ ), .X(\us11\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1360_ ( .A1(\us11\/_0020_ ), .A2(\us11\/_0137_ ), .B1(\us11\/_0261_ ), .B2(\us11\/_0128_ ), .Y(\us11\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1361_ ( .A(\us11\/_0573_ ), .B(\us11\/_0576_ ), .C(\us11\/_0579_ ), .D(\us11\/_0580_ ), .X(\us11\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1362_ ( .A(\us11\/_0561_ ), .B(\us11\/_0563_ ), .C(\us11\/_0570_ ), .D(\us11\/_0581_ ), .X(\us11\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1363_ ( .A(\us11\/_0128_ ), .B(\us11\/_0193_ ), .X(\us11\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1364_ ( .A(\us11\/_0082_ ), .B(\us11\/_0162_ ), .X(\us11\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us11/_1365_ ( .A(\us11\/_0583_ ), .B(\us11\/_0584_ ), .C_N(\us11\/_0437_ ), .Y(\us11\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us11/_1366_ ( .A(\us11\/_0150_ ), .B(\us11\/_0118_ ), .C(\us11\/_0380_ ), .Y(\us11\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us11/_1367_ ( .A_N(\us11\/_0182_ ), .B(\us11\/_0587_ ), .C(\us11\/_0323_ ), .X(\us11\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1368_ ( .A1(\us11\/_0575_ ), .A2(\us11\/_0153_ ), .B1(\us11\/_0727_ ), .B2(\us11\/_0058_ ), .Y(\us11\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1369_ ( .A1(\us11\/_0499_ ), .A2(\us11\/_0064_ ), .B1(\us11\/_0134_ ), .B2(\us11\/_0255_ ), .Y(\us11\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1370_ ( .A(\us11\/_0585_ ), .B(\us11\/_0588_ ), .C(\us11\/_0589_ ), .D(\us11\/_0590_ ), .X(\us11\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us11/_1371_ ( .A1(\us11\/_0091_ ), .A2(\us11\/_0139_ ), .B1(\us11\/_0250_ ), .Y(\us11\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1372_ ( .A1(\us11\/_0092_ ), .A2(\us11\/_0739_ ), .B1(\us11\/_0324_ ), .B2(\us11\/_0247_ ), .Y(\us11\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1373_ ( .A1(\us11\/_0144_ ), .A2(\us11\/_0153_ ), .B1(\us11\/_0683_ ), .B2(\us11\/_0292_ ), .Y(\us11\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1374_ ( .A1(\us11\/_0091_ ), .A2(\us11\/_0499_ ), .B1(\us11\/_0330_ ), .B2(\us11\/_0292_ ), .Y(\us11\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1375_ ( .A(\us11\/_0592_ ), .B(\us11\/_0593_ ), .C(\us11\/_0594_ ), .D(\us11\/_0595_ ), .X(\us11\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1376_ ( .A(\us11\/_0499_ ), .B(\us11\/_0144_ ), .Y(\us11\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1377_ ( .A(\us11\/_0312_ ), .B(\us11\/_0598_ ), .Y(\us11\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1378_ ( .A(\us11\/_0575_ ), .B(\us11\/_0147_ ), .Y(\us11\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1379_ ( .A1(\us11\/_0293_ ), .A2(\us11\/_0137_ ), .B1(\us11\/_0093_ ), .B2(\us11\/_0739_ ), .Y(\us11\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1380_ ( .A1(\us11\/_0734_ ), .A2(\us11\/_0531_ ), .B1(\us11\/_0600_ ), .C1(\us11\/_0601_ ), .Y(\us11\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1381_ ( .A1(\us11\/_0153_ ), .A2(\us11\/_0261_ ), .B1(\us11\/_0599_ ), .C1(\us11\/_0602_ ), .Y(\us11\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1382_ ( .A(\us11\/_0591_ ), .B(\us11\/_0596_ ), .C(\us11\/_0174_ ), .D(\us11\/_0603_ ), .X(\us11\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1383_ ( .A(\us11\/_0247_ ), .B(\us11\/_0144_ ), .Y(\us11\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1384_ ( .A(\us11\/_0113_ ), .B(\us11\/_0017_ ), .Y(\us11\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1385_ ( .A(\us11\/_0381_ ), .B(\us11\/_0605_ ), .C(\us11\/_0361_ ), .D(\us11\/_0606_ ), .X(\us11\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1386_ ( .A1(\us11\/_0016_ ), .A2(\us11\/_0727_ ), .B1(\us11\/_0733_ ), .Y(\us11\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1387_ ( .A1(\us11\/_0586_ ), .A2(\us11\/_0159_ ), .B1(\us11\/_0082_ ), .B2(\us11\/_0750_ ), .Y(\us11\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1388_ ( .A1(\us11\/_0142_ ), .A2(\us11\/_0162_ ), .B1(\us11\/_0079_ ), .B2(\us11\/_0054_ ), .Y(\us11\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1389_ ( .A(\us11\/_0610_ ), .B(\us11\/_0611_ ), .C(\us11\/_0105_ ), .D(\us11\/_0106_ ), .X(\us11\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1390_ ( .A1(\us11\/_0094_ ), .A2(\us11\/_0302_ ), .B1(\us11\/_0324_ ), .B2(\us11\/_0089_ ), .Y(\us11\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1391_ ( .A(\us11\/_0607_ ), .B(\us11\/_0609_ ), .C(\us11\/_0612_ ), .D(\us11\/_0613_ ), .X(\us11\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1392_ ( .A(\us11\/_0041_ ), .B(\us11\/_0170_ ), .X(\us11\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1393_ ( .A(\us11\/_0554_ ), .B(\us11\/_0027_ ), .X(\us11\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1394_ ( .A(\us11\/_0027_ ), .B(\us11\/_0261_ ), .Y(\us11\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us11/_1395_ ( .A_N(\us11\/_0616_ ), .B(\us11\/_0617_ ), .Y(\us11\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1396_ ( .A1(\us11\/_0147_ ), .A2(\us11\/_0302_ ), .B1(\us11\/_0342_ ), .C1(\us11\/_0618_ ), .Y(\us11\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1397_ ( .A(\us11\/_0614_ ), .B(\us11\/_0272_ ), .C(\us11\/_0615_ ), .D(\us11\/_0620_ ), .X(\us11\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us11/_1398_ ( .A(\us11\/_0582_ ), .B(\us11\/_0604_ ), .C(\us11\/_0621_ ), .Y(\us11\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1399_ ( .A1(\us11\/_0084_ ), .A2(\us11\/_0134_ ), .B1(\us11\/_0089_ ), .Y(\us11\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1400_ ( .A1(\us11\/_0144_ ), .A2(\us11\/_0608_ ), .A3(\us11\/_0330_ ), .B1(\us11\/_0089_ ), .Y(\us11\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1401_ ( .A1(\us11\/_0197_ ), .A2(\us11\/_0130_ ), .A3(\us11\/_0110_ ), .B1(\us11\/_0094_ ), .Y(\us11\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1402_ ( .A(\us11\/_0432_ ), .B(\us11\/_0622_ ), .C(\us11\/_0623_ ), .D(\us11\/_0624_ ), .X(\us11\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us11/_1403_ ( .A1(\us11\/_0554_ ), .A2(\us11\/_0017_ ), .A3(\us11\/_0022_ ), .B1(\us11\/_0161_ ), .X(\us11\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us11/_1404_ ( .A_N(\us11\/_0269_ ), .B(\us11\/_0170_ ), .X(\us11\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1405_ ( .A1(\us11\/_0109_ ), .A2(\us11\/_0064_ ), .A3(\us11\/_0733_ ), .B1(\us11\/_0355_ ), .Y(\us11\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us11/_1406_ ( .A_N(\us11\/_0626_ ), .B(\us11\/_0627_ ), .C(\us11\/_0353_ ), .D(\us11\/_0628_ ), .X(\us11\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1407_ ( .A1(\us11\/_0091_ ), .A2(\us11\/_0110_ ), .A3(\us11\/_0176_ ), .B1(\us11\/_0139_ ), .Y(\us11\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1408_ ( .A1(\us11\/_0020_ ), .A2(\us11\/_0261_ ), .B1(\us11\/_0147_ ), .Y(\us11\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1409_ ( .A(\us11\/_0631_ ), .B(\us11\/_0344_ ), .C(\us11\/_0421_ ), .D(\us11\/_0632_ ), .X(\us11\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us11/_1410_ ( .A1(\us11\/_0325_ ), .A2(\us11\/_0734_ ), .B1(\us11\/_0038_ ), .C1(\us11\/_0113_ ), .X(\us11\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1411_ ( .A1(\us11\/_0134_ ), .A2(\us11\/_0114_ ), .B1(\us11\/_0221_ ), .C1(\us11\/_0634_ ), .Y(\us11\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us11/_1412_ ( .A(\us11\/_0119_ ), .B_N(\us11\/_0111_ ), .Y(\us11\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1413_ ( .A1(\us11\/_0032_ ), .A2(\us11\/_0113_ ), .B1(\us11\/_0636_ ), .C1(\us11\/_0400_ ), .Y(\us11\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1414_ ( .A1(\us11\/_0732_ ), .A2(\us11\/_0293_ ), .A3(\us11\/_0251_ ), .B1(\us11\/_0364_ ), .Y(\us11\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1415_ ( .A(\us11\/_0189_ ), .B(\us11\/_0635_ ), .C(\us11\/_0637_ ), .D(\us11\/_0638_ ), .X(\us11\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1416_ ( .A(\us11\/_0625_ ), .B(\us11\/_0630_ ), .C(\us11\/_0633_ ), .D(\us11\/_0639_ ), .X(\us11\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1417_ ( .A(\us11\/_0746_ ), .B(\us11\/_0738_ ), .X(\us11\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1418_ ( .A(\us11\/_0736_ ), .B(\us11\/_0731_ ), .X(\us11\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us11/_1419_ ( .A_N(\us11\/_0643_ ), .B(\us11\/_0577_ ), .Y(\us11\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1420_ ( .A1(\us11\/_0084_ ), .A2(\us11\/_0739_ ), .B1(\us11\/_0642_ ), .C1(\us11\/_0644_ ), .Y(\us11\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1421_ ( .A1(\us11\/_0050_ ), .A2(\us11\/_0543_ ), .B1(\us11\/_0194_ ), .C1(\us11\/_0738_ ), .Y(\us11\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1422_ ( .A(\us11\/_0646_ ), .B(\us11\/_0232_ ), .C(\us11\/_0417_ ), .D(\us11\/_0578_ ), .X(\us11\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1423_ ( .A1(\us11\/_0064_ ), .A2(\us11\/_0733_ ), .B1(\us11\/_0727_ ), .Y(\us11\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1424_ ( .A1(\us11\/_0193_ ), .A2(\us11\/_0276_ ), .B1(\us11\/_0727_ ), .Y(\us11\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1425_ ( .A(\us11\/_0645_ ), .B(\us11\/_0647_ ), .C(\us11\/_0648_ ), .D(\us11\/_0649_ ), .X(\us11\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1426_ ( .A1(\us11\/_0325_ ), .A2(\us11\/_0734_ ), .B1(\us11\/_0038_ ), .C1(\us11\/_0247_ ), .Y(\us11\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1427_ ( .A1(\us11\/_0543_ ), .A2(\us11\/_0216_ ), .B1(\us11\/_0423_ ), .C1(\us11\/_0247_ ), .Y(\us11\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1428_ ( .A(\us11\/_0652_ ), .B(\us11\/_0653_ ), .X(\us11\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1429_ ( .A1(\us11\/_0733_ ), .A2(\us11\/_0748_ ), .A3(\us11\/_0324_ ), .B1(\us11\/_0016_ ), .Y(\us11\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1430_ ( .A1(\us11\/_0640_ ), .A2(\us11\/_0193_ ), .A3(\us11\/_0091_ ), .B1(\us11\/_0016_ ), .Y(\us11\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1431_ ( .A1(\us11\/_0102_ ), .A2(\us11\/_0301_ ), .B1(\sa11\[3\] ), .C1(\us11\/_0247_ ), .Y(\us11\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1432_ ( .A(\us11\/_0654_ ), .B(\us11\/_0655_ ), .C(\us11\/_0656_ ), .D(\us11\/_0657_ ), .X(\us11\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1433_ ( .A1(\us11\/_0118_ ), .A2(\us11\/_0050_ ), .B1(\us11\/_0038_ ), .C1(\us11\/_0478_ ), .Y(\us11\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us11/_1434_ ( .A_N(\us11\/_0250_ ), .B(\us11\/_0465_ ), .C(\us11\/_0659_ ), .X(\us11\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1435_ ( .A1(\us11\/_0683_ ), .A2(\us11\/_0324_ ), .B1(\us11\/_0255_ ), .Y(\us11\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1436_ ( .A1(\us11\/_0032_ ), .A2(\us11\/_0193_ ), .A3(\us11\/_0047_ ), .B1(\us11\/_0255_ ), .Y(\us11\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1437_ ( .A1(\us11\/_0144_ ), .A2(\us11\/_0586_ ), .A3(\us11\/_0047_ ), .B1(\us11\/_0499_ ), .Y(\us11\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1438_ ( .A(\us11\/_0660_ ), .B(\us11\/_0661_ ), .C(\us11\/_0663_ ), .D(\us11\/_0664_ ), .X(\us11\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1439_ ( .A1(\us11\/_0091_ ), .A2(\us11\/_0276_ ), .B1(\us11\/_0060_ ), .Y(\us11\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1440_ ( .A1(\us11\/_0144_ ), .A2(\us11\/_0608_ ), .B1(\us11\/_0292_ ), .Y(\us11\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1441_ ( .A1(\us11\/_0423_ ), .A2(\us11\/_0038_ ), .B1(\us11\/_0102_ ), .C1(\us11\/_0060_ ), .Y(\us11\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1442_ ( .A1(\sa11\[1\] ), .A2(\us11\/_0734_ ), .B1(\us11\/_0109_ ), .C1(\us11\/_0292_ ), .Y(\us11\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1443_ ( .A(\us11\/_0666_ ), .B(\us11\/_0667_ ), .C(\us11\/_0668_ ), .D(\us11\/_0669_ ), .X(\us11\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1444_ ( .A(\us11\/_0650_ ), .B(\us11\/_0658_ ), .C(\us11\/_0665_ ), .D(\us11\/_0670_ ), .X(\us11\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us11/_1445_ ( .A(\us11\/_0641_ ), .B(\us11\/_0174_ ), .C(\us11\/_0671_ ), .Y(\us11\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us11/_1446_ ( .A(\us11\/_0049_ ), .B(\us11\/_0618_ ), .C_N(\us11\/_0052_ ), .Y(\us11\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us11/_1447_ ( .A(\us11\/_0239_ ), .Y(\us11\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1448_ ( .A(\us11\/_0705_ ), .B(\us11\/_0032_ ), .Y(\us11\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1449_ ( .A1(\us11\/_0054_ ), .A2(\us11\/_0732_ ), .B1(\us11\/_0035_ ), .B2(\us11\/_0705_ ), .Y(\us11\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1450_ ( .A1(\us11\/_0304_ ), .A2(\us11\/_0732_ ), .B1(\us11\/_0047_ ), .B2(\us11\/_0750_ ), .Y(\us11\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1451_ ( .A(\us11\/_0674_ ), .B(\us11\/_0675_ ), .C(\us11\/_0676_ ), .D(\us11\/_0677_ ), .X(\us11\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us11/_1452_ ( .A_N(\us11\/_0584_ ), .B(\us11\/_0283_ ), .X(\us11\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1453_ ( .A(\us11\/_0673_ ), .B(\us11\/_0678_ ), .C(\us11\/_0679_ ), .D(\us11\/_0508_ ), .X(\us11\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1454_ ( .A1(\us11\/_0016_ ), .A2(\us11\/_0733_ ), .B1(\us11\/_0355_ ), .B2(\us11\/_0092_ ), .Y(\us11\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1455_ ( .A(\us11\/_0681_ ), .B(\us11\/_0034_ ), .X(\us11\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us11/_1456_ ( .A1(\us11\/_0330_ ), .A2(\us11\/_0139_ ), .B1(\us11\/_0324_ ), .B2(\us11\/_0089_ ), .X(\us11\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1457_ ( .A1(\us11\/_0146_ ), .A2(\us11\/_0147_ ), .B1(\us11\/_0133_ ), .C1(\us11\/_0684_ ), .Y(\us11\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1458_ ( .A(\us11\/_0113_ ), .B(\us11\/_0251_ ), .Y(\us11\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us11/_1459_ ( .A_N(\us11\/_0463_ ), .B(\us11\/_0686_ ), .C(\us11\/_0383_ ), .D(\us11\/_0464_ ), .X(\us11\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1460_ ( .A1(\us11\/_0051_ ), .A2(\us11\/_0293_ ), .B1(\us11\/_0084_ ), .B2(\us11\/_0705_ ), .Y(\us11\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1461_ ( .A1(\us11\/_0017_ ), .A2(\us11\/_0072_ ), .B1(\us11\/_0134_ ), .B2(\us11\/_0078_ ), .Y(\us11\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1462_ ( .A(\us11\/_0687_ ), .B(\us11\/_0236_ ), .C(\us11\/_0688_ ), .D(\us11\/_0689_ ), .X(\us11\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1463_ ( .A(\us11\/_0680_ ), .B(\us11\/_0682_ ), .C(\us11\/_0685_ ), .D(\us11\/_0690_ ), .X(\us11\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us11/_1464_ ( .A1(\us11\/_0532_ ), .A2(\us11\/_0380_ ), .B1(\us11\/_0102_ ), .C1(\us11\/_0355_ ), .X(\us11\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us11/_1465_ ( .A(\us11\/_0692_ ), .B(\us11\/_0338_ ), .C(\us11\/_0644_ ), .Y(\us11\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1466_ ( .A(\us11\/_0016_ ), .B(\us11\/_0020_ ), .Y(\us11\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1467_ ( .A1(\us11\/_0032_ ), .A2(\us11\/_0137_ ), .B1(\us11\/_0279_ ), .B2(\us11\/_0094_ ), .Y(\us11\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1468_ ( .A1(\us11\/_0575_ ), .A2(\us11\/_0153_ ), .B1(\us11\/_0161_ ), .B2(\us11\/_0293_ ), .Y(\us11\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1469_ ( .A(\us11\/_0259_ ), .B(\us11\/_0695_ ), .C(\us11\/_0696_ ), .D(\us11\/_0697_ ), .X(\us11\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us11/_1470_ ( .A1(\us11\/_0255_ ), .A2(\us11\/_0640_ ), .B1(\us11\/_0016_ ), .B2(\us11\/_0193_ ), .X(\us11\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1471_ ( .A1(\us11\/_0060_ ), .A2(\us11\/_0176_ ), .B1(\us11\/_0699_ ), .C1(\us11\/_0177_ ), .Y(\us11\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1472_ ( .A1(\us11\/_0091_ ), .A2(\us11\/_0499_ ), .B1(\us11\/_0092_ ), .B2(\us11\/_0705_ ), .Y(\us11\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us11/_1473_ ( .A1(\us11\/_0705_ ), .A2(\us11\/_0683_ ), .B1(\us11\/_0093_ ), .B2(\us11\/_0114_ ), .Y(\us11\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us11/_1474_ ( .A1(\us11\/_0683_ ), .A2(\us11\/_0084_ ), .B1(\us11\/_0094_ ), .Y(\us11\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us11/_1475_ ( .A1(\us11\/_0543_ ), .A2(\us11\/_0216_ ), .B1(\us11\/_0038_ ), .C1(\us11\/_0292_ ), .Y(\us11\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1476_ ( .A(\us11\/_0701_ ), .B(\us11\/_0702_ ), .C(\us11\/_0703_ ), .D(\us11\/_0704_ ), .X(\us11\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1477_ ( .A(\us11\/_0693_ ), .B(\us11\/_0698_ ), .C(\us11\/_0700_ ), .D(\us11\/_0706_ ), .X(\us11\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us11/_1478_ ( .A1(\us11\/_0113_ ), .A2(\us11\/_0640_ ), .B1(\us11\/_0364_ ), .B2(\us11\/_0058_ ), .X(\us11\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us11/_1479_ ( .A(\us11\/_0407_ ), .B(\us11\/_0708_ ), .C(\us11\/_0529_ ), .Y(\us11\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1480_ ( .A(\us11\/_0568_ ), .B(\us11\/_0175_ ), .Y(\us11\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us11/_1481_ ( .A1(\us11\/_0247_ ), .A2(\us11\/_0114_ ), .A3(\us11\/_0051_ ), .B1(\us11\/_0130_ ), .Y(\us11\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1482_ ( .A(\us11\/_0709_ ), .B(\us11\/_0550_ ), .C(\us11\/_0710_ ), .D(\us11\/_0711_ ), .X(\us11\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us11/_1483_ ( .A1(\us11\/_0114_ ), .A2(\us11\/_0064_ ), .B1(\us11\/_0261_ ), .B2(\us11\/_0089_ ), .X(\us11\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1484_ ( .A1(\us11\/_0355_ ), .A2(\us11\/_0261_ ), .B1(\us11\/_0198_ ), .C1(\us11\/_0713_ ), .Y(\us11\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1485_ ( .A(\us11\/_0586_ ), .B(\us11\/_0478_ ), .Y(\us11\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us11/_1486_ ( .A_N(\us11\/_0541_ ), .B(\us11\/_0267_ ), .C(\us11\/_0715_ ), .D(\us11\/_0320_ ), .X(\us11\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1487_ ( .A(\us11\/_0586_ ), .B(\us11\/_0070_ ), .Y(\us11\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us11/_1488_ ( .A_N(\us11\/_0211_ ), .B(\us11\/_0155_ ), .C(\us11\/_0202_ ), .D(\us11\/_0718_ ), .X(\us11\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us11/_1489_ ( .A(\us11\/_0150_ ), .B(\us11\/_0216_ ), .C(\us11\/_0380_ ), .Y(\us11\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us11/_1490_ ( .A(\us11\/_0411_ ), .B(\us11\/_0720_ ), .X(\us11\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us11/_1491_ ( .A1(\us11\/_0017_ ), .A2(\us11\/_0022_ ), .B1(\us11\/_0078_ ), .X(\us11\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us11/_1492_ ( .A1(\us11\/_0134_ ), .A2(\us11\/_0738_ ), .B1(\us11\/_0101_ ), .C1(\us11\/_0722_ ), .Y(\us11\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1493_ ( .A(\us11\/_0717_ ), .B(\us11\/_0719_ ), .C(\us11\/_0721_ ), .D(\us11\/_0723_ ), .X(\us11\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us11/_1494_ ( .A(\us11\/_0739_ ), .B(\us11\/_0193_ ), .Y(\us11\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1495_ ( .A(\us11\/_0344_ ), .B(\us11\/_0184_ ), .C(\us11\/_0449_ ), .D(\us11\/_0725_ ), .X(\us11\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us11/_1496_ ( .A(\us11\/_0712_ ), .B(\us11\/_0714_ ), .C(\us11\/_0724_ ), .D(\us11\/_0726_ ), .X(\us11\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \us11/_1497_ ( .A(\us11\/_0691_ ), .B(\us11\/_0707_ ), .C(\us11\/_0728_ ), .Y(\us11\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \us12/_0753_ ( .A(\sa12\[2\] ), .B_N(\sa12\[3\] ), .Y(\us12\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0755_ ( .A(\sa12\[1\] ), .B(\sa12\[0\] ), .X(\us12\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0756_ ( .A(\us12\/_0096_ ), .B(\us12\/_0118_ ), .X(\us12\/_0129_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0757_ ( .A(\sa12\[7\] ), .B(\sa12\[6\] ), .X(\us12\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_0758_ ( .A(\sa12\[4\] ), .B(\sa12\[5\] ), .Y(\us12\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0759_ ( .A(\us12\/_0140_ ), .B(\us12\/_0151_ ), .X(\us12\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0761_ ( .A(\us12\/_0129_ ), .B(\us12\/_0162_ ), .X(\us12\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0762_ ( .A(\us12\/_0096_ ), .X(\us12\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \us12/_0763_ ( .A(\sa12\[1\] ), .B_N(\sa12\[0\] ), .Y(\us12\/_0205_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0764_ ( .A(\us12\/_0205_ ), .X(\us12\/_0216_ ) );
sky130_fd_sc_hd__and3_1 \us12/_0765_ ( .A(\us12\/_0162_ ), .B(\us12\/_0194_ ), .C(\us12\/_0216_ ), .X(\us12\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us12/_0766_ ( .A(\us12\/_0183_ ), .SLEEP(\us12\/_0227_ ), .X(\us12\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \us12/_0767_ ( .A(\sa12\[0\] ), .B_N(\sa12\[1\] ), .Y(\us12\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_0768_ ( .A(\sa12\[2\] ), .B(\sa12\[3\] ), .Y(\us12\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0769_ ( .A(\us12\/_0249_ ), .B(\us12\/_0260_ ), .X(\us12\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0771_ ( .A(\us12\/_0271_ ), .X(\us12\/_0293_ ) );
sky130_fd_sc_hd__buf_2 \us12/_0772_ ( .A(\us12\/_0162_ ), .X(\us12\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_0773_ ( .A(\us12\/_0293_ ), .B(\us12\/_0304_ ), .Y(\us12\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us12/_0774_ ( .A(\sa12\[1\] ), .Y(\us12\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us12/_0776_ ( .A(\sa12\[0\] ), .Y(\us12\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0777_ ( .A(\sa12\[2\] ), .B(\sa12\[3\] ), .X(\us12\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0779_ ( .A(\us12\/_0358_ ), .X(\us12\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_0780_ ( .A1(\us12\/_0325_ ), .A2(\us12\/_0347_ ), .B1(\us12\/_0380_ ), .C1(\us12\/_0304_ ), .Y(\us12\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us12/_0781_ ( .A_N(\us12\/_0238_ ), .B(\us12\/_0314_ ), .C(\us12\/_0391_ ), .X(\us12\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us12/_0782_ ( .A(\sa12\[3\] ), .B_N(\sa12\[2\] ), .Y(\us12\/_0412_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0783_ ( .A(\us12\/_0412_ ), .X(\us12\/_0423_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0784_ ( .A(\us12\/_0423_ ), .B(\us12\/_0205_ ), .X(\us12\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \us12/_0787_ ( .A(\sa12\[5\] ), .B_N(\sa12\[4\] ), .Y(\us12\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0788_ ( .A(\us12\/_0467_ ), .B(\us12\/_0140_ ), .X(\us12\/_0478_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0789_ ( .A(\us12\/_0478_ ), .X(\us12\/_0489_ ) );
sky130_fd_sc_hd__buf_2 \us12/_0790_ ( .A(\us12\/_0489_ ), .X(\us12\/_0499_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_0791_ ( .A(\us12\/_0134_ ), .B(\us12\/_0499_ ), .Y(\us12\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_0792_ ( .A(\us12\/_0489_ ), .B(\us12\/_0271_ ), .Y(\us12\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0793_ ( .A(\us12\/_0194_ ), .X(\us12\/_0532_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0794_ ( .A(\us12\/_0249_ ), .X(\us12\/_0543_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0795_ ( .A(\us12\/_0543_ ), .B(\us12\/_0358_ ), .X(\us12\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0797_ ( .A(\us12\/_0554_ ), .X(\us12\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0798_ ( .A(\us12\/_0216_ ), .B(\us12\/_0358_ ), .X(\us12\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0800_ ( .A(\us12\/_0586_ ), .X(\us12\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_0801_ ( .A1(\us12\/_0532_ ), .A2(\us12\/_0575_ ), .A3(\us12\/_0608_ ), .B1(\us12\/_0499_ ), .Y(\us12\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us12/_0802_ ( .A(\us12\/_0401_ ), .B(\us12\/_0510_ ), .C(\us12\/_0521_ ), .D(\us12\/_0619_ ), .X(\us12\/_0629_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0803_ ( .A(\us12\/_0358_ ), .B(\sa12\[1\] ), .X(\us12\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0805_ ( .A(\us12\/_0205_ ), .B(\us12\/_0260_ ), .X(\us12\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0807_ ( .A(\us12\/_0662_ ), .X(\us12\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us12/_0808_ ( .A(\sa12\[6\] ), .B_N(\sa12\[7\] ), .Y(\us12\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0809_ ( .A(\us12\/_0467_ ), .B(\us12\/_0694_ ), .X(\us12\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0811_ ( .A(\us12\/_0705_ ), .X(\us12\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_0812_ ( .A1(\us12\/_0640_ ), .A2(\us12\/_0293_ ), .A3(\us12\/_0683_ ), .B1(\us12\/_0727_ ), .Y(\us12\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_0813_ ( .A(\sa12\[1\] ), .B(\sa12\[0\] ), .Y(\us12\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0814_ ( .A(\us12\/_0730_ ), .B(\us12\/_0260_ ), .X(\us12\/_0731_ ) );
sky130_fd_sc_hd__buf_1 \us12/_0815_ ( .A(\us12\/_0731_ ), .X(\us12\/_0732_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0816_ ( .A(\us12\/_0732_ ), .X(\us12\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0817_ ( .A(\sa12\[0\] ), .X(\us12\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us12/_0818_ ( .A1(\us12\/_0325_ ), .A2(\us12\/_0734_ ), .B1(\us12\/_0423_ ), .X(\us12\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0819_ ( .A(\us12\/_0694_ ), .B(\us12\/_0151_ ), .X(\us12\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0821_ ( .A(\us12\/_0736_ ), .X(\us12\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0822_ ( .A(\us12\/_0738_ ), .X(\us12\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_0823_ ( .A1(\us12\/_0733_ ), .A2(\us12\/_0735_ ), .A3(\us12\/_0293_ ), .B1(\us12\/_0739_ ), .Y(\us12\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us12/_0824_ ( .A(\us12\/_0730_ ), .B_N(\us12\/_0358_ ), .Y(\us12\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_0825_ ( .A(\us12\/_0741_ ), .B(\us12\/_0739_ ), .Y(\us12\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_0827_ ( .A1(\us12\/_0118_ ), .A2(\us12\/_0216_ ), .B1(\us12\/_0532_ ), .C1(\us12\/_0739_ ), .Y(\us12\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us12/_0828_ ( .A(\us12\/_0729_ ), .B(\us12\/_0740_ ), .C(\us12\/_0742_ ), .D(\us12\/_0744_ ), .X(\us12\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0829_ ( .A(\us12\/_0423_ ), .B(\us12\/_0730_ ), .X(\us12\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0830_ ( .A(\us12\/_0746_ ), .X(\us12\/_0747_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0831_ ( .A(\us12\/_0747_ ), .X(\us12\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us12/_0832_ ( .A(\sa12\[4\] ), .B_N(\sa12\[5\] ), .Y(\us12\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0833_ ( .A(\us12\/_0749_ ), .B(\us12\/_0694_ ), .X(\us12\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0835_ ( .A(\us12\/_0750_ ), .X(\us12\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0836_ ( .A(\us12\/_0752_ ), .X(\us12\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0837_ ( .A(\us12\/_0118_ ), .B(\us12\/_0358_ ), .X(\us12\/_0017_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0838_ ( .A(\us12\/_0017_ ), .X(\us12\/_0018_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0839_ ( .A(\us12\/_0752_ ), .B(\us12\/_0018_ ), .X(\us12\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0840_ ( .A(\us12\/_0358_ ), .B(\us12\/_0325_ ), .X(\us12\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0842_ ( .A(\us12\/_0096_ ), .B(\us12\/_0205_ ), .X(\us12\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \us12/_0844_ ( .A1(\us12\/_0020_ ), .A2(\us12\/_0022_ ), .B1(\us12\/_0752_ ), .X(\us12\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_0845_ ( .A1(\us12\/_0748_ ), .A2(\us12\/_0016_ ), .B1(\us12\/_0019_ ), .C1(\us12\/_0024_ ), .Y(\us12\/_0025_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0846_ ( .A(\sa12\[4\] ), .B(\sa12\[5\] ), .X(\us12\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0847_ ( .A(\us12\/_0694_ ), .B(\us12\/_0026_ ), .X(\us12\/_0027_ ) );
sky130_fd_sc_hd__buf_2 \us12/_0849_ ( .A(\us12\/_0027_ ), .X(\us12\/_0029_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0850_ ( .A(\us12\/_0358_ ), .B(\us12\/_0730_ ), .X(\us12\/_0030_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0852_ ( .A(\us12\/_0030_ ), .X(\us12\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_0853_ ( .A(\us12\/_0029_ ), .B(\us12\/_0032_ ), .Y(\us12\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_0854_ ( .A(\us12\/_0029_ ), .B(\us12\/_0735_ ), .Y(\us12\/_0034_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0855_ ( .A(\us12\/_0118_ ), .B(\us12\/_0260_ ), .X(\us12\/_0035_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0857_ ( .A(\us12\/_0027_ ), .B(\us12\/_0035_ ), .X(\us12\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0858_ ( .A(\us12\/_0260_ ), .X(\us12\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_0859_ ( .A(\us12\/_0038_ ), .B(\us12\/_0347_ ), .Y(\us12\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us12/_0860_ ( .A_N(\us12\/_0039_ ), .B(\us12\/_0027_ ), .X(\us12\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_0861_ ( .A(\us12\/_0037_ ), .B(\us12\/_0040_ ), .Y(\us12\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us12/_0862_ ( .A(\us12\/_0025_ ), .B(\us12\/_0033_ ), .C(\us12\/_0034_ ), .D(\us12\/_0041_ ), .X(\us12\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0863_ ( .A(\us12\/_0749_ ), .B(\us12\/_0140_ ), .X(\us12\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us12/_0865_ ( .A(\sa12\[0\] ), .B(\sa12\[2\] ), .C(\sa12\[3\] ), .X(\us12\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0866_ ( .A(\us12\/_0043_ ), .B(\us12\/_0045_ ), .X(\us12\/_0046_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0867_ ( .A(\us12\/_0096_ ), .B(\us12\/_0543_ ), .X(\us12\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0869_ ( .A(\us12\/_0047_ ), .B(\us12\/_0043_ ), .X(\us12\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0870_ ( .A(\us12\/_0730_ ), .X(\us12\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0871_ ( .A(\us12\/_0043_ ), .X(\us12\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_0872_ ( .A1(\us12\/_0118_ ), .A2(\us12\/_0050_ ), .B1(\us12\/_0194_ ), .C1(\us12\/_0051_ ), .Y(\us12\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us12/_0873_ ( .A(\us12\/_0046_ ), .B(\us12\/_0049_ ), .C_N(\us12\/_0052_ ), .Y(\us12\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0874_ ( .A(\us12\/_0026_ ), .B(\us12\/_0140_ ), .X(\us12\/_0054_ ) );
sky130_fd_sc_hd__buf_2 \us12/_0876_ ( .A(\us12\/_0054_ ), .X(\us12\/_0056_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_0877_ ( .A1(\us12\/_0532_ ), .A2(\us12\/_0575_ ), .B1(\us12\/_0056_ ), .Y(\us12\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0878_ ( .A(\us12\/_0423_ ), .B(\us12\/_0325_ ), .X(\us12\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0880_ ( .A(\us12\/_0051_ ), .X(\us12\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_0881_ ( .A1(\us12\/_0732_ ), .A2(\us12\/_0035_ ), .A3(\us12\/_0058_ ), .B1(\us12\/_0060_ ), .Y(\us12\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0882_ ( .A(\us12\/_0260_ ), .B(\sa12\[1\] ), .X(\us12\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0884_ ( .A(\us12\/_0062_ ), .X(\us12\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_0885_ ( .A1(\us12\/_0064_ ), .A2(\us12\/_0748_ ), .A3(\us12\/_0683_ ), .B1(\us12\/_0056_ ), .Y(\us12\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us12/_0886_ ( .A(\us12\/_0053_ ), .B(\us12\/_0057_ ), .C(\us12\/_0061_ ), .D(\us12\/_0065_ ), .X(\us12\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us12/_0887_ ( .A(\us12\/_0629_ ), .B(\us12\/_0745_ ), .C(\us12\/_0042_ ), .D(\us12\/_0066_ ), .X(\us12\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us12/_0889_ ( .A(\sa12\[7\] ), .B_N(\sa12\[6\] ), .Y(\us12\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0890_ ( .A(\us12\/_0069_ ), .B(\us12\/_0151_ ), .X(\us12\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0892_ ( .A(\us12\/_0070_ ), .X(\us12\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_0893_ ( .A1(\us12\/_0129_ ), .A2(\us12\/_0586_ ), .B1(\us12\/_0072_ ), .Y(\us12\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_0894_ ( .A1(\us12\/_0380_ ), .A2(\us12\/_0347_ ), .B1(\us12\/_0194_ ), .B2(\us12\/_0216_ ), .Y(\us12\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us12/_0895_ ( .A(\us12\/_0074_ ), .B_N(\us12\/_0070_ ), .Y(\us12\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us12/_0896_ ( .A(\us12\/_0073_ ), .SLEEP(\us12\/_0075_ ), .X(\us12\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0897_ ( .A(\us12\/_0467_ ), .B(\us12\/_0069_ ), .X(\us12\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0898_ ( .A(\us12\/_0077_ ), .X(\us12\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0899_ ( .A(\us12\/_0412_ ), .B(\us12\/_0118_ ), .X(\us12\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0901_ ( .A(\us12\/_0078_ ), .B(\us12\/_0079_ ), .X(\us12\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0902_ ( .A(\us12\/_0412_ ), .B(\us12\/_0249_ ), .X(\us12\/_0082_ ) );
sky130_fd_sc_hd__buf_2 \us12/_0904_ ( .A(\us12\/_0082_ ), .X(\us12\/_0084_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0905_ ( .A(\us12\/_0084_ ), .B(\us12\/_0078_ ), .X(\us12\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us12/_0906_ ( .A1(\sa12\[0\] ), .A2(\us12\/_0325_ ), .B1(\us12\/_0260_ ), .Y(\us12\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us12/_0907_ ( .A_N(\us12\/_0086_ ), .B(\us12\/_0078_ ), .X(\us12\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us12/_0908_ ( .A(\us12\/_0081_ ), .B(\us12\/_0085_ ), .C(\us12\/_0087_ ), .Y(\us12\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0909_ ( .A(\us12\/_0072_ ), .X(\us12\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_0910_ ( .A1(\us12\/_0733_ ), .A2(\us12\/_0748_ ), .A3(\us12\/_0683_ ), .B1(\us12\/_0089_ ), .Y(\us12\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0911_ ( .A(\us12\/_0129_ ), .X(\us12\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0912_ ( .A(\us12\/_0018_ ), .X(\us12\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0913_ ( .A(\us12\/_0022_ ), .X(\us12\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0914_ ( .A(\us12\/_0078_ ), .X(\us12\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_0915_ ( .A1(\us12\/_0091_ ), .A2(\us12\/_0092_ ), .A3(\us12\/_0093_ ), .B1(\us12\/_0094_ ), .Y(\us12\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us12/_0916_ ( .A(\us12\/_0076_ ), .B(\us12\/_0088_ ), .C(\us12\/_0090_ ), .D(\us12\/_0095_ ), .X(\us12\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0917_ ( .A(\us12\/_0069_ ), .B(\us12\/_0026_ ), .X(\us12\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \us12/_0918_ ( .A(\us12\/_0098_ ), .X(\us12\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0919_ ( .A(\us12\/_0434_ ), .B(\us12\/_0099_ ), .X(\us12\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0920_ ( .A(\us12\/_0079_ ), .B(\us12\/_0098_ ), .X(\us12\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0921_ ( .A(\us12\/_0325_ ), .X(\us12\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_0922_ ( .A1(\us12\/_0102_ ), .A2(\us12\/_0734_ ), .B1(\us12\/_0038_ ), .C1(\us12\/_0099_ ), .Y(\us12\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us12/_0923_ ( .A(\us12\/_0100_ ), .B(\us12\/_0101_ ), .C_N(\us12\/_0103_ ), .Y(\us12\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_0924_ ( .A1(\us12\/_0554_ ), .A2(\us12\/_0586_ ), .B1(\us12\/_0099_ ), .Y(\us12\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_0925_ ( .A(\us12\/_0129_ ), .B(\us12\/_0099_ ), .Y(\us12\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0926_ ( .A(\us12\/_0105_ ), .B(\us12\/_0106_ ), .X(\us12\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0927_ ( .A(\us12\/_0423_ ), .X(\us12\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0928_ ( .A(\us12\/_0260_ ), .B(\sa12\[0\] ), .X(\us12\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0929_ ( .A(\us12\/_0069_ ), .B(\us12\/_0749_ ), .X(\us12\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0931_ ( .A(\us12\/_0111_ ), .X(\us12\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0932_ ( .A(\us12\/_0113_ ), .X(\us12\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_0933_ ( .A1(\us12\/_0109_ ), .A2(\us12\/_0110_ ), .B1(\us12\/_0114_ ), .Y(\us12\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us12/_0934_ ( .A(\us12\/_0022_ ), .Y(\us12\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us12/_0935_ ( .A(\us12\/_0554_ ), .Y(\us12\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us12/_0936_ ( .A1(\us12\/_0050_ ), .A2(\us12\/_0118_ ), .B1(\us12\/_0194_ ), .Y(\us12\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us12/_0937_ ( .A(\us12\/_0113_ ), .Y(\us12\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us12/_0938_ ( .A1(\us12\/_0116_ ), .A2(\us12\/_0117_ ), .A3(\us12\/_0119_ ), .B1(\us12\/_0120_ ), .X(\us12\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us12/_0939_ ( .A(\us12\/_0104_ ), .B(\us12\/_0108_ ), .C(\us12\/_0115_ ), .D(\us12\/_0121_ ), .X(\us12\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_0940_ ( .A(\sa12\[7\] ), .B(\sa12\[6\] ), .Y(\us12\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0941_ ( .A(\us12\/_0749_ ), .B(\us12\/_0123_ ), .X(\us12\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0943_ ( .A(\us12\/_0082_ ), .B(\us12\/_0124_ ), .X(\us12\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_0944_ ( .A(\us12\/_0271_ ), .B(\us12\/_0124_ ), .Y(\us12\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0945_ ( .A(\us12\/_0124_ ), .X(\us12\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0946_ ( .A(\us12\/_0260_ ), .B(\us12\/_0325_ ), .X(\us12\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_0948_ ( .A(\us12\/_0128_ ), .B(\us12\/_0130_ ), .Y(\us12\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_0949_ ( .A(\us12\/_0127_ ), .B(\us12\/_0132_ ), .Y(\us12\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us12/_0950_ ( .A(\us12\/_0434_ ), .X(\us12\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_0951_ ( .A(\us12\/_0134_ ), .B(\us12\/_0128_ ), .Y(\us12\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us12/_0952_ ( .A(\us12\/_0126_ ), .B(\us12\/_0133_ ), .C_N(\us12\/_0135_ ), .Y(\us12\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0953_ ( .A(\us12\/_0026_ ), .B(\us12\/_0123_ ), .X(\us12\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0955_ ( .A(\us12\/_0137_ ), .X(\us12\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_0956_ ( .A1(\us12\/_0110_ ), .A2(\us12\/_0293_ ), .A3(\us12\/_0084_ ), .B1(\us12\/_0139_ ), .Y(\us12\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0957_ ( .A(\us12\/_0096_ ), .B(\us12\/_0730_ ), .X(\us12\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0959_ ( .A(\us12\/_0142_ ), .X(\us12\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_0960_ ( .A1(\us12\/_0020_ ), .A2(\us12\/_0144_ ), .A3(\us12\/_0018_ ), .B1(\us12\/_0139_ ), .Y(\us12\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \us12/_0961_ ( .A(\sa12\[2\] ), .B(\us12\/_0050_ ), .C_N(\sa12\[3\] ), .Y(\us12\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0962_ ( .A(\us12\/_0128_ ), .X(\us12\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_0963_ ( .A1(\us12\/_0146_ ), .A2(\us12\/_0032_ ), .A3(\us12\/_0640_ ), .B1(\us12\/_0147_ ), .Y(\us12\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us12/_0964_ ( .A(\us12\/_0136_ ), .B(\us12\/_0141_ ), .C(\us12\/_0145_ ), .D(\us12\/_0148_ ), .X(\us12\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0965_ ( .A(\us12\/_0123_ ), .B(\us12\/_0151_ ), .X(\us12\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0967_ ( .A(\us12\/_0150_ ), .X(\us12\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0968_ ( .A(\us12\/_0150_ ), .B(\us12\/_0062_ ), .X(\us12\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_0969_ ( .A(\us12\/_0079_ ), .B(\us12\/_0150_ ), .Y(\us12\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us12/_0970_ ( .A(\us12\/_0150_ ), .B(\us12\/_0423_ ), .C(\us12\/_0543_ ), .Y(\us12\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_0971_ ( .A(\us12\/_0155_ ), .B(\us12\/_0156_ ), .Y(\us12\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_0972_ ( .A1(\us12\/_0153_ ), .A2(\us12\/_0134_ ), .B1(\us12\/_0154_ ), .C1(\us12\/_0157_ ), .Y(\us12\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0973_ ( .A(\us12\/_0467_ ), .B(\us12\/_0123_ ), .X(\us12\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_0975_ ( .A(\us12\/_0159_ ), .X(\us12\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us12/_0976_ ( .A_N(\us12\/_0119_ ), .B(\us12\/_0161_ ), .X(\us12\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us12/_0977_ ( .A(\us12\/_0163_ ), .Y(\us12\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_0978_ ( .A1(\us12\/_0146_ ), .A2(\us12\/_0575_ ), .A3(\us12\/_0608_ ), .B1(\us12\/_0153_ ), .Y(\us12\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_0979_ ( .A1(\us12\/_0062_ ), .A2(\us12\/_0084_ ), .A3(\us12\/_0134_ ), .B1(\us12\/_0161_ ), .Y(\us12\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us12/_0980_ ( .A(\us12\/_0158_ ), .B(\us12\/_0164_ ), .C(\us12\/_0165_ ), .D(\us12\/_0166_ ), .X(\us12\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us12/_0981_ ( .A(\us12\/_0097_ ), .B(\us12\/_0122_ ), .C(\us12\/_0149_ ), .D(\us12\/_0167_ ), .X(\us12\/_0168_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0982_ ( .A(\us12\/_0662_ ), .B(\us12\/_0150_ ), .X(\us12\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_0983_ ( .A(\us12\/_0154_ ), .B(\us12\/_0169_ ), .Y(\us12\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us12/_0984_ ( .A(\us12\/_0123_ ), .B(\us12\/_0151_ ), .C(\us12\/_0038_ ), .X(\us12\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0985_ ( .A(\us12\/_0170_ ), .B(\us12\/_0171_ ), .X(\us12\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \us12/_0986_ ( .A(\us12\/_0172_ ), .Y(\us12\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \us12/_0987_ ( .A(\us12\/_0067_ ), .B(\us12\/_0168_ ), .C(\us12\/_0174_ ), .Y(\us12\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us12/_0988_ ( .A(\sa12\[1\] ), .B(\sa12\[0\] ), .Y(\us12\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us12/_0989_ ( .A(\us12\/_0175_ ), .B(\us12\/_0358_ ), .X(\us12\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0990_ ( .A(\us12\/_0176_ ), .B(\us12\/_0489_ ), .X(\us12\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_0991_ ( .A(\us12\/_0084_ ), .B(\us12\/_0113_ ), .Y(\us12\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0992_ ( .A(\us12\/_0111_ ), .B(\us12\/_0062_ ), .X(\us12\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0993_ ( .A(\us12\/_0111_ ), .B(\us12\/_0662_ ), .X(\us12\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_0994_ ( .A(\us12\/_0179_ ), .B(\us12\/_0180_ ), .Y(\us12\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0995_ ( .A(\us12\/_0054_ ), .B(\us12\/_0058_ ), .X(\us12\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us12/_0996_ ( .A(\us12\/_0182_ ), .Y(\us12\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us12/_0997_ ( .A_N(\us12\/_0177_ ), .B(\us12\/_0178_ ), .C(\us12\/_0181_ ), .D(\us12\/_0184_ ), .X(\us12\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0998_ ( .A(\us12\/_0098_ ), .B(\us12\/_0741_ ), .X(\us12\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us12/_0999_ ( .A(\us12\/_0047_ ), .B(\us12\/_0098_ ), .X(\us12\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us12/_1000_ ( .A(\us12\/_0186_ ), .B(\us12\/_0187_ ), .X(\us12\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1001_ ( .A(\us12\/_0188_ ), .Y(\us12\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1002_ ( .A(\us12\/_0738_ ), .B(\us12\/_0735_ ), .X(\us12\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1003_ ( .A(\us12\/_0271_ ), .B(\us12\/_0736_ ), .X(\us12\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_1004_ ( .A(\us12\/_0190_ ), .B(\us12\/_0191_ ), .Y(\us12\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us12/_1005_ ( .A(\us12\/_0096_ ), .B(\us12\/_0325_ ), .X(\us12\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1006_ ( .A1(\us12\/_0193_ ), .A2(\us12\/_0176_ ), .B1(\us12\/_0043_ ), .Y(\us12\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1007_ ( .A(\us12\/_0185_ ), .B(\us12\/_0189_ ), .C(\us12\/_0192_ ), .D(\us12\/_0195_ ), .X(\us12\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us12/_1008_ ( .A_N(\sa12\[3\] ), .B(\us12\/_0734_ ), .C(\sa12\[2\] ), .X(\us12\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1009_ ( .A(\us12\/_0137_ ), .B(\us12\/_0197_ ), .X(\us12\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_1010_ ( .A(\us12\/_0198_ ), .B(\us12\/_0040_ ), .Y(\us12\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1011_ ( .A(\us12\/_0293_ ), .B(\us12\/_0137_ ), .X(\us12\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1012_ ( .A(\us12\/_0200_ ), .Y(\us12\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1013_ ( .A(\us12\/_0137_ ), .B(\us12\/_0110_ ), .Y(\us12\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1014_ ( .A(\us12\/_0139_ ), .B(\us12\/_0020_ ), .Y(\us12\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1015_ ( .A(\us12\/_0199_ ), .B(\us12\/_0201_ ), .C(\us12\/_0202_ ), .D(\us12\/_0203_ ), .X(\us12\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us12/_1016_ ( .A1(\us12\/_0532_ ), .A2(\us12\/_0109_ ), .B1(\us12\/_0102_ ), .C1(\us12\/_0727_ ), .X(\us12\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1017_ ( .A(\us12\/_0022_ ), .B(\us12\/_0078_ ), .Y(\us12\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1018_ ( .A(\us12\/_0078_ ), .B(\us12\/_0142_ ), .Y(\us12\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1019_ ( .A(\us12\/_0207_ ), .B(\us12\/_0208_ ), .Y(\us12\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1020_ ( .A1(\us12\/_0094_ ), .A2(\us12\/_0176_ ), .B1(\us12\/_0206_ ), .C1(\us12\/_0209_ ), .Y(\us12\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1021_ ( .A(\us12\/_0662_ ), .B(\us12\/_0070_ ), .X(\us12\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us12/_1022_ ( .A(\us12\/_0732_ ), .B(\us12\/_0123_ ), .C(\us12\/_0749_ ), .Y(\us12\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us12/_1023_ ( .A(\us12\/_0732_ ), .B(\us12\/_0467_ ), .C(\us12\/_0069_ ), .Y(\us12\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us12/_1024_ ( .A_N(\us12\/_0211_ ), .B(\us12\/_0127_ ), .C(\us12\/_0212_ ), .D(\us12\/_0213_ ), .X(\us12\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1025_ ( .A(\us12\/_0137_ ), .Y(\us12\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1026_ ( .A(\us12\/_0128_ ), .B(\us12\/_0035_ ), .Y(\us12\/_0217_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1028_ ( .A1(\us12\/_0159_ ), .A2(\us12\/_0747_ ), .B1(\us12\/_0434_ ), .B2(\us12\/_0499_ ), .Y(\us12\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us12/_1029_ ( .A1(\us12\/_0116_ ), .A2(\us12\/_0215_ ), .B1(\us12\/_0217_ ), .C1(\us12\/_0219_ ), .X(\us12\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1030_ ( .A(\us12\/_0113_ ), .B(\us12\/_0746_ ), .X(\us12\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us12/_1031_ ( .A1(\us12\/_0098_ ), .A2(\us12\/_0746_ ), .B1(\us12\/_0434_ ), .B2(\us12\/_0750_ ), .X(\us12\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1032_ ( .A1(\us12\/_0047_ ), .A2(\us12\/_0113_ ), .B1(\us12\/_0221_ ), .C1(\us12\/_0222_ ), .Y(\us12\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us12/_1033_ ( .A1(\us12\/_0129_ ), .A2(\us12\/_0162_ ), .B1(\us12\/_0271_ ), .B2(\us12\/_0705_ ), .X(\us12\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1034_ ( .A1(\us12\/_0093_ ), .A2(\us12\/_0738_ ), .B1(\us12\/_0081_ ), .C1(\us12\/_0224_ ), .Y(\us12\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1035_ ( .A(\us12\/_0214_ ), .B(\us12\/_0220_ ), .C(\us12\/_0223_ ), .D(\us12\/_0225_ ), .X(\us12\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1036_ ( .A(\us12\/_0196_ ), .B(\us12\/_0204_ ), .C(\us12\/_0210_ ), .D(\us12\/_0226_ ), .X(\us12\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1037_ ( .A(\us12\/_0111_ ), .B(\us12\/_0554_ ), .X(\us12\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1038_ ( .A(\us12\/_0229_ ), .Y(\us12\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1039_ ( .A(\us12\/_0111_ ), .B(\us12\/_0129_ ), .Y(\us12\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1040_ ( .A(\us12\/_0018_ ), .B(\us12\/_0738_ ), .Y(\us12\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1041_ ( .A(\us12\/_0030_ ), .B(\us12\/_0304_ ), .Y(\us12\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1042_ ( .A(\us12\/_0230_ ), .B(\us12\/_0231_ ), .C(\us12\/_0232_ ), .D(\us12\/_0233_ ), .X(\us12\/_0234_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1043_ ( .A(\us12\/_0047_ ), .B(\us12\/_0489_ ), .X(\us12\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1044_ ( .A1(\us12\/_0129_ ), .A2(\us12\/_0554_ ), .B1(\us12\/_0137_ ), .Y(\us12\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us12/_1045_ ( .A(\us12\/_0235_ ), .B(\us12\/_0049_ ), .C_N(\us12\/_0236_ ), .Y(\us12\/_0237_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1046_ ( .A(\us12\/_0047_ ), .B(\us12\/_0077_ ), .X(\us12\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1047_ ( .A(\us12\/_0070_ ), .B(\us12\/_0035_ ), .X(\us12\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us12/_1048_ ( .A1(\us12\/_0047_ ), .A2(\us12\/_0736_ ), .B1(\us12\/_0022_ ), .B2(\us12\/_0099_ ), .X(\us12\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us12/_1049_ ( .A(\us12\/_0239_ ), .B(\us12\/_0240_ ), .C(\us12\/_0241_ ), .Y(\us12\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1050_ ( .A(\us12\/_0554_ ), .B(\us12\/_0072_ ), .X(\us12\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us12/_1051_ ( .A1(\us12\/_0142_ ), .A2(\us12\/_0137_ ), .B1(\us12\/_0159_ ), .B2(\us12\/_0082_ ), .X(\us12\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1052_ ( .A1(\us12\/_0608_ ), .A2(\us12\/_0072_ ), .B1(\us12\/_0243_ ), .C1(\us12\/_0244_ ), .Y(\us12\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1053_ ( .A(\us12\/_0234_ ), .B(\us12\/_0237_ ), .C(\us12\/_0242_ ), .D(\us12\/_0245_ ), .X(\us12\/_0246_ ) );
sky130_fd_sc_hd__o21a_1 \us12/_1055_ ( .A1(\us12\/_0554_ ), .A2(\us12\/_0586_ ), .B1(\us12\/_0029_ ), .X(\us12\/_0248_ ) );
sky130_fd_sc_hd__and2_1 \us12/_1056_ ( .A(\us12\/_0082_ ), .B(\us12\/_0489_ ), .X(\us12\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_1057_ ( .A(\us12\/_0079_ ), .X(\us12\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1058_ ( .A(\us12\/_0251_ ), .B(\us12\/_0489_ ), .X(\us12\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_1059_ ( .A(\us12\/_0250_ ), .B(\us12\/_0252_ ), .Y(\us12\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1060_ ( .A(\us12\/_0016_ ), .B(\us12\/_0064_ ), .Y(\us12\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_1061_ ( .A(\us12\/_0304_ ), .X(\us12\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1062_ ( .A(\us12\/_0255_ ), .B(\us12\/_0640_ ), .Y(\us12\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us12/_1063_ ( .A_N(\us12\/_0248_ ), .B(\us12\/_0253_ ), .C(\us12\/_0254_ ), .D(\us12\/_0256_ ), .X(\us12\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1064_ ( .A(\us12\/_0099_ ), .B(\us12\/_0110_ ), .X(\us12\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us12/_1065_ ( .A1(\us12\/_0161_ ), .A2(\us12\/_0130_ ), .B1(\us12\/_0258_ ), .Y(\us12\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1066_ ( .A(\us12\/_0194_ ), .B(\sa12\[1\] ), .X(\us12\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1068_ ( .A(\us12\/_0261_ ), .B(\us12\/_0153_ ), .Y(\us12\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us12/_1069_ ( .A_N(\us12\/_0154_ ), .B(\us12\/_0259_ ), .C(\us12\/_0263_ ), .X(\us12\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1070_ ( .A(\us12\/_0246_ ), .B(\us12\/_0174_ ), .C(\us12\/_0257_ ), .D(\us12\/_0264_ ), .X(\us12\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us12/_1071_ ( .A1(\us12\/_0261_ ), .A2(\us12\/_0554_ ), .B1(\us12\/_0159_ ), .X(\us12\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1072_ ( .A(\us12\/_0747_ ), .B(\us12\/_0150_ ), .Y(\us12\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1073_ ( .A(\us12\/_0175_ ), .Y(\us12\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us12/_1074_ ( .A(\us12\/_0423_ ), .B(\us12\/_0123_ ), .C(\us12\/_0151_ ), .X(\us12\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1075_ ( .A(\us12\/_0268_ ), .B(\us12\/_0269_ ), .Y(\us12\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us12/_1076_ ( .A_N(\us12\/_0266_ ), .B(\us12\/_0267_ ), .C(\us12\/_0270_ ), .X(\us12\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1077_ ( .A(\us12\/_0554_ ), .B(\us12\/_0150_ ), .X(\us12\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1078_ ( .A(\us12\/_0273_ ), .Y(\us12\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1079_ ( .A1(\us12\/_0734_ ), .A2(\us12\/_0325_ ), .B1(\us12\/_0380_ ), .Y(\us12\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1080_ ( .A(\us12\/_0275_ ), .Y(\us12\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1081_ ( .A(\us12\/_0276_ ), .B(\us12\/_0153_ ), .Y(\us12\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us12/_1082_ ( .A(\us12\/_0272_ ), .B(\us12\/_0274_ ), .C(\us12\/_0277_ ), .X(\us12\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_1083_ ( .A(\us12\/_0035_ ), .X(\us12\/_0279_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1085_ ( .A1(\us12\/_0499_ ), .A2(\us12\/_0279_ ), .B1(\us12\/_0084_ ), .B2(\us12\/_0060_ ), .Y(\us12\/_0281_ ) );
sky130_fd_sc_hd__o21ai_1 \us12/_1086_ ( .A1(\us12\/_0251_ ), .A2(\us12\/_0434_ ), .B1(\us12\/_0304_ ), .Y(\us12\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1087_ ( .A(\us12\/_0091_ ), .B(\us12\/_0056_ ), .Y(\us12\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1088_ ( .A1(\us12\/_0118_ ), .A2(\us12\/_0050_ ), .B1(\us12\/_0038_ ), .C1(\us12\/_0255_ ), .Y(\us12\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1089_ ( .A(\us12\/_0281_ ), .B(\us12\/_0283_ ), .C(\us12\/_0284_ ), .D(\us12\/_0285_ ), .X(\us12\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1090_ ( .A(\us12\/_0082_ ), .B(\us12\/_0027_ ), .X(\us12\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1091_ ( .A(\us12\/_0129_ ), .B(\us12\/_0027_ ), .X(\us12\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_1092_ ( .A(\us12\/_0287_ ), .B(\us12\/_0288_ ), .Y(\us12\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1093_ ( .A1(\us12\/_0752_ ), .A2(\us12\/_0683_ ), .B1(\us12\/_0093_ ), .B2(\us12\/_0029_ ), .Y(\us12\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1094_ ( .A1(\us12\/_0092_ ), .A2(\us12\/_0575_ ), .B1(\us12\/_0056_ ), .Y(\us12\/_0291_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1096_ ( .A1(\us12\/_0499_ ), .A2(\us12\/_0662_ ), .B1(\us12\/_0084_ ), .B2(\us12\/_0056_ ), .Y(\us12\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1097_ ( .A(\us12\/_0289_ ), .B(\us12\/_0290_ ), .C(\us12\/_0291_ ), .D(\us12\/_0294_ ), .X(\us12\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1098_ ( .A(\us12\/_0750_ ), .B(\us12\/_0193_ ), .X(\us12\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1099_ ( .A(\us12\/_0705_ ), .B(\us12\/_0380_ ), .X(\us12\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1100_ ( .A(\us12\/_0752_ ), .B(\us12\/_0129_ ), .Y(\us12\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us12/_1101_ ( .A(\us12\/_0296_ ), .B(\us12\/_0297_ ), .C_N(\us12\/_0298_ ), .Y(\us12\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1102_ ( .A(\us12\/_0089_ ), .B(\us12\/_0532_ ), .Y(\us12\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1103_ ( .A(\sa12\[2\] ), .Y(\us12\/_0301_ ) );
sky130_fd_sc_hd__nor3_2 \us12/_1104_ ( .A(\us12\/_0301_ ), .B(\sa12\[3\] ), .C(\us12\/_0118_ ), .Y(\us12\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1105_ ( .A(\us12\/_0072_ ), .B(\us12\/_0302_ ), .X(\us12\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1106_ ( .A(\us12\/_0303_ ), .Y(\us12\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1107_ ( .A(\us12\/_0147_ ), .B(\us12\/_0302_ ), .Y(\us12\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1108_ ( .A(\us12\/_0299_ ), .B(\us12\/_0300_ ), .C(\us12\/_0305_ ), .D(\us12\/_0306_ ), .X(\us12\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1109_ ( .A(\us12\/_0278_ ), .B(\us12\/_0286_ ), .C(\us12\/_0295_ ), .D(\us12\/_0307_ ), .X(\us12\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us12/_1110_ ( .A(\us12\/_0228_ ), .B(\us12\/_0265_ ), .C(\us12\/_0308_ ), .Y(\us12\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1111_ ( .A(\us12\/_0235_ ), .Y(\us12\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1112_ ( .A(\us12\/_0489_ ), .B(\us12\/_0640_ ), .X(\us12\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1113_ ( .A(\us12\/_0310_ ), .Y(\us12\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1114_ ( .A(\us12\/_0022_ ), .B(\us12\/_0499_ ), .Y(\us12\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1115_ ( .A(\us12\/_0499_ ), .B(\us12\/_0032_ ), .Y(\us12\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1116_ ( .A(\us12\/_0309_ ), .B(\us12\/_0311_ ), .C(\us12\/_0312_ ), .D(\us12\/_0313_ ), .X(\us12\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1117_ ( .A(\us12\/_0499_ ), .B(\us12\/_0064_ ), .Y(\us12\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1118_ ( .A(\us12\/_0499_ ), .B(\us12\/_0683_ ), .Y(\us12\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1119_ ( .A(\us12\/_0315_ ), .B(\us12\/_0316_ ), .C(\us12\/_0317_ ), .D(\us12\/_0253_ ), .X(\us12\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1120_ ( .A(\us12\/_0047_ ), .B(\us12\/_0304_ ), .Y(\us12\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1121_ ( .A(\us12\/_0586_ ), .B(\us12\/_0162_ ), .Y(\us12\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1122_ ( .A(\us12\/_0319_ ), .B(\us12\/_0320_ ), .Y(\us12\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_1123_ ( .A(\us12\/_0321_ ), .B(\us12\/_0238_ ), .Y(\us12\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1124_ ( .A(\us12\/_0304_ ), .B(\us12\/_0062_ ), .Y(\us12\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_1125_ ( .A(\us12\/_0251_ ), .X(\us12\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1126_ ( .A1(\us12\/_0324_ ), .A2(\us12\/_0084_ ), .B1(\us12\/_0255_ ), .Y(\us12\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1127_ ( .A1(\us12\/_0050_ ), .A2(\us12\/_0216_ ), .B1(\us12\/_0109_ ), .C1(\us12\/_0255_ ), .Y(\us12\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1128_ ( .A(\us12\/_0322_ ), .B(\us12\/_0323_ ), .C(\us12\/_0326_ ), .D(\us12\/_0327_ ), .X(\us12\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1129_ ( .A1(\us12\/_0733_ ), .A2(\us12\/_0279_ ), .A3(\us12\/_0058_ ), .B1(\us12\/_0056_ ), .Y(\us12\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_1130_ ( .A(\us12\/_0047_ ), .X(\us12\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1131_ ( .A(\us12\/_0330_ ), .B(\us12\/_0056_ ), .Y(\us12\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1132_ ( .A(\us12\/_0054_ ), .B(\us12\/_0045_ ), .Y(\us12\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1133_ ( .A(\us12\/_0329_ ), .B(\us12\/_0331_ ), .C(\us12\/_0284_ ), .D(\us12\/_0332_ ), .X(\us12\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us12/_1134_ ( .A1(\us12\/_0543_ ), .A2(\us12\/_0216_ ), .B1(\us12\/_0532_ ), .C1(\us12\/_0060_ ), .X(\us12\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1135_ ( .A(\us12\/_0084_ ), .B(\us12\/_0060_ ), .Y(\us12\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1136_ ( .A(\us12\/_0324_ ), .B(\us12\/_0060_ ), .Y(\us12\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1137_ ( .A(\us12\/_0335_ ), .B(\us12\/_0337_ ), .Y(\us12\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1138_ ( .A1(\us12\/_0276_ ), .A2(\us12\/_0060_ ), .B1(\us12\/_0334_ ), .C1(\us12\/_0338_ ), .Y(\us12\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1139_ ( .A(\us12\/_0318_ ), .B(\us12\/_0328_ ), .C(\us12\/_0333_ ), .D(\us12\/_0339_ ), .X(\us12\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us12/_1140_ ( .A1(\us12\/_0747_ ), .A2(\us12\/_0134_ ), .B1(\us12\/_0128_ ), .X(\us12\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us12/_1141_ ( .A_N(\us12\/_0086_ ), .B(\us12\/_0128_ ), .X(\us12\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1142_ ( .A(\us12\/_0079_ ), .B(\us12\/_0124_ ), .X(\us12\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_1143_ ( .A(\us12\/_0126_ ), .B(\us12\/_0343_ ), .Y(\us12\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us12/_1144_ ( .A(\us12\/_0341_ ), .B(\us12\/_0342_ ), .C_N(\us12\/_0344_ ), .Y(\us12\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1146_ ( .A1(\us12\/_0193_ ), .A2(\us12\/_0092_ ), .A3(\us12\/_0330_ ), .B1(\us12\/_0147_ ), .Y(\us12\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1147_ ( .A1(\us12\/_0130_ ), .A2(\us12\/_0084_ ), .A3(\us12\/_0134_ ), .B1(\us12\/_0139_ ), .Y(\us12\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1148_ ( .A1(\us12\/_0144_ ), .A2(\us12\/_0608_ ), .A3(\us12\/_0092_ ), .B1(\us12\/_0139_ ), .Y(\us12\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1149_ ( .A(\us12\/_0345_ ), .B(\us12\/_0348_ ), .C(\us12\/_0349_ ), .D(\us12\/_0350_ ), .X(\us12\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us12/_1150_ ( .A(\us12\/_0150_ ), .B(\us12\/_0194_ ), .C(\us12\/_0543_ ), .X(\us12\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us12/_1151_ ( .A(\us12\/_0277_ ), .SLEEP(\us12\/_0352_ ), .X(\us12\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us12/_1152_ ( .A1(\us12\/_0268_ ), .A2(\us12\/_0171_ ), .B1(\us12\/_0157_ ), .Y(\us12\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us12/_1153_ ( .A(\us12\/_0161_ ), .X(\us12\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1154_ ( .A1(\us12\/_0279_ ), .A2(\us12\/_0084_ ), .B1(\us12\/_0355_ ), .Y(\us12\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1155_ ( .A1(\us12\/_0020_ ), .A2(\us12\/_0193_ ), .A3(\us12\/_0091_ ), .B1(\us12\/_0355_ ), .Y(\us12\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1156_ ( .A(\us12\/_0353_ ), .B(\us12\/_0354_ ), .C(\us12\/_0356_ ), .D(\us12\/_0357_ ), .X(\us12\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1157_ ( .A(\us12\/_0111_ ), .B(\us12\/_0586_ ), .X(\us12\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1158_ ( .A(\us12\/_0360_ ), .Y(\us12\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us12/_1159_ ( .A1(\us12\/_0119_ ), .A2(\us12\/_0120_ ), .B1(\us12\/_0230_ ), .C1(\us12\/_0361_ ), .X(\us12\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1160_ ( .A1(\us12\/_0662_ ), .A2(\us12\/_0251_ ), .A3(\us12\/_0134_ ), .B1(\us12\/_0114_ ), .Y(\us12\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1162_ ( .A1(\us12\/_0035_ ), .A2(\us12\/_0251_ ), .A3(\us12\/_0134_ ), .B1(\us12\/_0099_ ), .Y(\us12\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1163_ ( .A1(\us12\/_0193_ ), .A2(\us12\/_0608_ ), .B1(\us12\/_0099_ ), .Y(\us12\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1164_ ( .A(\us12\/_0362_ ), .B(\us12\/_0363_ ), .C(\us12\/_0365_ ), .D(\us12\/_0366_ ), .X(\us12\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1165_ ( .A1(\us12\/_0575_ ), .A2(\us12\/_0092_ ), .A3(\us12\/_0330_ ), .B1(\us12\/_0089_ ), .Y(\us12\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1166_ ( .A1(\us12\/_0586_ ), .A2(\us12\/_0018_ ), .A3(\us12\/_0330_ ), .B1(\us12\/_0094_ ), .Y(\us12\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \us12/_1167_ ( .A1(\us12\/_0293_ ), .A2(\us12\/_0134_ ), .B1(\us12\/_0089_ ), .Y(\us12\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1168_ ( .A1(\us12\/_0279_ ), .A2(\us12\/_0134_ ), .B1(\us12\/_0094_ ), .Y(\us12\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1169_ ( .A(\us12\/_0368_ ), .B(\us12\/_0370_ ), .C(\us12\/_0371_ ), .D(\us12\/_0372_ ), .X(\us12\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1170_ ( .A(\us12\/_0351_ ), .B(\us12\/_0359_ ), .C(\us12\/_0367_ ), .D(\us12\/_0373_ ), .X(\us12\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1171_ ( .A1(\us12\/_0102_ ), .A2(\us12\/_0347_ ), .B1(\us12\/_0109_ ), .C1(\us12\/_0029_ ), .Y(\us12\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1172_ ( .A1(\us12\/_0102_ ), .A2(\us12\/_0347_ ), .B1(\us12\/_0532_ ), .C1(\us12\/_0029_ ), .Y(\us12\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1173_ ( .A1(\us12\/_0050_ ), .A2(\us12\/_0543_ ), .B1(\us12\/_0380_ ), .C1(\us12\/_0029_ ), .Y(\us12\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1174_ ( .A(\us12\/_0041_ ), .B(\us12\/_0375_ ), .C(\us12\/_0376_ ), .D(\us12\/_0377_ ), .X(\us12\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1175_ ( .A(\us12\/_0047_ ), .B(\us12\/_0750_ ), .X(\us12\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1176_ ( .A(\us12\/_0379_ ), .Y(\us12\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1177_ ( .A(\us12\/_0016_ ), .B(\us12\/_0608_ ), .Y(\us12\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1178_ ( .A(\us12\/_0752_ ), .B(\us12\/_0554_ ), .Y(\us12\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1179_ ( .A1(\sa12\[1\] ), .A2(\us12\/_0734_ ), .B1(\us12\/_0109_ ), .C1(\us12\/_0016_ ), .Y(\us12\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1180_ ( .A(\us12\/_0381_ ), .B(\us12\/_0382_ ), .C(\us12\/_0383_ ), .D(\us12\/_0384_ ), .X(\us12\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us12/_1181_ ( .A(\us12\/_0086_ ), .B_N(\us12\/_0736_ ), .X(\us12\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1182_ ( .A1(\us12\/_0748_ ), .A2(\us12\/_0134_ ), .B1(\us12\/_0739_ ), .Y(\us12\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1183_ ( .A1(\us12\/_0118_ ), .A2(\us12\/_0543_ ), .B1(\us12\/_0109_ ), .C1(\us12\/_0739_ ), .Y(\us12\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1184_ ( .A1(\us12\/_0102_ ), .A2(\us12\/_0301_ ), .B1(\sa12\[3\] ), .C1(\us12\/_0739_ ), .Y(\us12\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1185_ ( .A(\us12\/_0386_ ), .B(\us12\/_0387_ ), .C(\us12\/_0388_ ), .D(\us12\/_0389_ ), .X(\us12\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1186_ ( .A(\us12\/_0020_ ), .Y(\us12\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1187_ ( .A(\us12\/_0727_ ), .Y(\us12\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1188_ ( .A(\us12\/_0727_ ), .B(\us12\/_0064_ ), .Y(\us12\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1189_ ( .A1(\us12\/_0102_ ), .A2(\us12\/_0734_ ), .B1(\us12\/_0532_ ), .C1(\us12\/_0727_ ), .Y(\us12\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us12/_1190_ ( .A1(\us12\/_0392_ ), .A2(\us12\/_0393_ ), .B1(\us12\/_0394_ ), .C1(\us12\/_0395_ ), .X(\us12\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1191_ ( .A(\us12\/_0378_ ), .B(\us12\/_0385_ ), .C(\us12\/_0390_ ), .D(\us12\/_0396_ ), .X(\us12\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us12/_1192_ ( .A(\us12\/_0340_ ), .B(\us12\/_0374_ ), .C(\us12\/_0397_ ), .Y(\us12\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1193_ ( .A(\us12\/_0077_ ), .B(\us12\/_0129_ ), .X(\us12\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_1194_ ( .A(\us12\/_0398_ ), .B(\us12\/_0239_ ), .Y(\us12\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1195_ ( .A(\us12\/_0022_ ), .B(\us12\/_0111_ ), .X(\us12\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us12/_1196_ ( .A_N(\us12\/_0400_ ), .B(\us12\/_0231_ ), .Y(\us12\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us12/_1197_ ( .A(\us12\/_0399_ ), .SLEEP(\us12\/_0402_ ), .X(\us12\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_1198_ ( .A(\us12\/_0747_ ), .B(\us12\/_0251_ ), .Y(\us12\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us12/_1199_ ( .A_N(\us12\/_0404_ ), .B(\us12\/_0752_ ), .Y(\us12\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us12/_1200_ ( .A(\us12\/_0467_ ), .B(\us12\/_0194_ ), .C(\us12\/_0694_ ), .X(\us12\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us12/_1201_ ( .A_N(\us12\/_0175_ ), .B(\us12\/_0406_ ), .X(\us12\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1202_ ( .A(\us12\/_0407_ ), .Y(\us12\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1203_ ( .A1(\us12\/_0094_ ), .A2(\us12\/_0197_ ), .B1(\us12\/_0114_ ), .B2(\us12\/_0640_ ), .Y(\us12\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1204_ ( .A(\us12\/_0403_ ), .B(\us12\/_0405_ ), .C(\us12\/_0408_ ), .D(\us12\/_0409_ ), .X(\us12\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1205_ ( .A(\us12\/_0030_ ), .B(\us12\/_0150_ ), .Y(\us12\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us12/_1206_ ( .A_N(\us12\/_0169_ ), .B(\us12\/_0289_ ), .C(\us12\/_0411_ ), .X(\us12\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us12/_1207_ ( .A1(\us12\/_0467_ ), .A2(\us12\/_0151_ ), .B1(\us12\/_0140_ ), .C1(\us12\/_0129_ ), .X(\us12\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1208_ ( .A1(\us12\/_0608_ ), .A2(\us12\/_0099_ ), .B1(\us12\/_0037_ ), .C1(\us12\/_0414_ ), .Y(\us12\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1209_ ( .A(\us12\/_0738_ ), .Y(\us12\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1210_ ( .A(\us12\/_0586_ ), .B(\us12\/_0736_ ), .Y(\us12\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1211_ ( .A1(\us12\/_0194_ ), .A2(\us12\/_0038_ ), .B1(\us12\/_0118_ ), .C1(\us12\/_0153_ ), .Y(\us12\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us12/_1212_ ( .A1(\us12\/_0416_ ), .A2(\us12\/_0117_ ), .B1(\us12\/_0417_ ), .C1(\us12\/_0418_ ), .X(\us12\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1213_ ( .A(\us12\/_0077_ ), .B(\us12\/_0035_ ), .X(\us12\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1214_ ( .A(\us12\/_0662_ ), .B(\us12\/_0124_ ), .Y(\us12\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1215_ ( .A(\us12\/_0030_ ), .B(\us12\/_0137_ ), .Y(\us12\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1216_ ( .A(\us12\/_0072_ ), .B(\us12\/_0732_ ), .Y(\us12\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us12/_1217_ ( .A_N(\us12\/_0420_ ), .B(\us12\/_0421_ ), .C(\us12\/_0422_ ), .D(\us12\/_0424_ ), .X(\us12\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1218_ ( .A(\us12\/_0413_ ), .B(\us12\/_0415_ ), .C(\us12\/_0419_ ), .D(\us12\/_0425_ ), .X(\us12\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us12/_1219_ ( .A(\us12\/_0355_ ), .B(\us12\/_0102_ ), .C(\us12\/_0109_ ), .Y(\us12\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1220_ ( .A(\us12\/_0077_ ), .B(\us12\/_0018_ ), .X(\us12\/_0428_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1221_ ( .A(\us12\/_0077_ ), .B(\us12\/_0554_ ), .X(\us12\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us12/_1222_ ( .A1(\us12\/_0050_ ), .A2(\us12\/_0216_ ), .B1(\us12\/_0380_ ), .C1(\us12\/_0078_ ), .X(\us12\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us12/_1223_ ( .A(\us12\/_0428_ ), .B(\us12\/_0429_ ), .C(\us12\/_0430_ ), .Y(\us12\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us12/_1224_ ( .A_N(\us12\/_0209_ ), .B(\us12\/_0431_ ), .X(\us12\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us12/_1225_ ( .A1(\us12\/_0215_ ), .A2(\us12\/_0404_ ), .B1(\us12\/_0427_ ), .C1(\us12\/_0432_ ), .X(\us12\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1226_ ( .A(\us12\/_0043_ ), .B(\us12\/_0058_ ), .Y(\us12\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1227_ ( .A(\us12\/_0195_ ), .B(\us12\/_0233_ ), .C(\us12\/_0320_ ), .D(\us12\/_0435_ ), .X(\us12\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1228_ ( .A(\us12\/_0261_ ), .B(\us12\/_0738_ ), .Y(\us12\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1229_ ( .A1(\us12\/_0499_ ), .A2(\us12\/_0640_ ), .B1(\us12\/_0261_ ), .B2(\us12\/_0056_ ), .Y(\us12\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1230_ ( .A(\us12\/_0436_ ), .B(\us12\/_0394_ ), .C(\us12\/_0437_ ), .D(\us12\/_0438_ ), .X(\us12\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1231_ ( .A(\us12\/_0410_ ), .B(\us12\/_0426_ ), .C(\us12\/_0433_ ), .D(\us12\/_0439_ ), .X(\us12\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us12/_1232_ ( .A(\us12\/_0135_ ), .SLEEP(\us12\/_0273_ ), .X(\us12\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1233_ ( .A1(\us12\/_0279_ ), .A2(\us12\/_0134_ ), .B1(\us12\/_0099_ ), .Y(\us12\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1234_ ( .A(\us12\/_0441_ ), .B(\us12\/_0164_ ), .C(\us12\/_0270_ ), .D(\us12\/_0442_ ), .X(\us12\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1235_ ( .A(\us12\/_0051_ ), .B(\us12\/_0662_ ), .Y(\us12\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1236_ ( .A(\us12\/_0051_ ), .B(\us12\/_0271_ ), .Y(\us12\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1237_ ( .A(\us12\/_0444_ ), .B(\us12\/_0446_ ), .X(\us12\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1238_ ( .A(\us12\/_0193_ ), .B(\us12\/_0304_ ), .X(\us12\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1239_ ( .A(\us12\/_0448_ ), .Y(\us12\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1240_ ( .A(\us12\/_0162_ ), .B(\us12\/_0130_ ), .X(\us12\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1241_ ( .A(\us12\/_0450_ ), .Y(\us12\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1242_ ( .A1(\us12\/_0129_ ), .A2(\us12\/_0554_ ), .B1(\us12\/_0043_ ), .Y(\us12\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1243_ ( .A(\us12\/_0447_ ), .B(\us12\/_0449_ ), .C(\us12\/_0451_ ), .D(\us12\/_0452_ ), .X(\us12\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1244_ ( .A(\us12\/_0056_ ), .B(\us12\/_0064_ ), .Y(\us12\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us12/_1245_ ( .A_N(\us12\/_0248_ ), .B(\us12\/_0454_ ), .C(\us12\/_0254_ ), .D(\us12\/_0256_ ), .X(\us12\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1246_ ( .A1(\us12\/_0330_ ), .A2(\us12\/_0099_ ), .B1(\us12\/_0134_ ), .B2(\us12\/_0705_ ), .Y(\us12\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1247_ ( .A1(\us12\/_0748_ ), .A2(\us12\/_0738_ ), .B1(\us12\/_0092_ ), .B2(\us12\/_0752_ ), .Y(\us12\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1248_ ( .A1(\us12\/_0072_ ), .A2(\us12\/_0035_ ), .B1(\us12\/_0748_ ), .B2(\us12\/_0056_ ), .Y(\us12\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1249_ ( .A1(\us12\/_0748_ ), .A2(\us12\/_0251_ ), .B1(\us12\/_0029_ ), .Y(\us12\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1250_ ( .A(\us12\/_0457_ ), .B(\us12\/_0458_ ), .C(\us12\/_0459_ ), .D(\us12\/_0460_ ), .X(\us12\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1251_ ( .A(\us12\/_0443_ ), .B(\us12\/_0453_ ), .C(\us12\/_0455_ ), .D(\us12\/_0461_ ), .X(\us12\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1252_ ( .A(\us12\/_0705_ ), .B(\us12\/_0079_ ), .X(\us12\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1253_ ( .A(\us12\/_0586_ ), .B(\us12\/_0124_ ), .Y(\us12\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1254_ ( .A(\us12\/_0499_ ), .B(\us12\/_0747_ ), .Y(\us12\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us12/_1255_ ( .A_N(\us12\/_0463_ ), .B(\us12\/_0464_ ), .C(\us12\/_0465_ ), .X(\us12\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us12/_1256_ ( .A1(\us12\/_0271_ ), .A2(\us12\/_0072_ ), .B1(\us12\/_0142_ ), .B2(\us12\/_0027_ ), .X(\us12\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1257_ ( .A1(\us12\/_0144_ ), .A2(\us12\/_0099_ ), .B1(\us12\/_0360_ ), .C1(\us12\/_0468_ ), .Y(\us12\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us12/_1258_ ( .A1(\us12\/_0662_ ), .A2(\us12\/_0251_ ), .B1(\us12\/_0499_ ), .X(\us12\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1259_ ( .A1(\us12\/_0575_ ), .A2(\us12\/_0056_ ), .B1(\us12\/_0379_ ), .C1(\us12\/_0470_ ), .Y(\us12\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1260_ ( .A(\us12\/_0466_ ), .B(\us12\/_0469_ ), .C(\us12\/_0471_ ), .D(\us12\/_0305_ ), .X(\us12\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us12/_1261_ ( .A1(\us12\/_0029_ ), .A2(\us12\/_0683_ ), .B1(\us12\/_0324_ ), .B2(\us12\/_0056_ ), .X(\us12\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1262_ ( .A(\us12\/_0084_ ), .B(\us12\/_0099_ ), .X(\us12\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us12/_1263_ ( .A1(\us12\/_0092_ ), .A2(\us12\/_0029_ ), .B1(\us12\/_0474_ ), .X(\us12\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us12/_1264_ ( .A(\us12\/_0075_ ), .B(\us12\/_0473_ ), .C(\us12\/_0475_ ), .Y(\us12\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1265_ ( .A1(\us12\/_0279_ ), .A2(\us12\/_0255_ ), .B1(\us12\/_0084_ ), .B2(\us12\/_0060_ ), .Y(\us12\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1266_ ( .A1(\us12\/_0093_ ), .A2(\us12\/_0056_ ), .B1(\us12\/_0134_ ), .B2(\us12\/_0114_ ), .Y(\us12\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1267_ ( .A1(\us12\/_0161_ ), .A2(\us12\/_0032_ ), .B1(\us12\/_0324_ ), .B2(\us12\/_0147_ ), .Y(\us12\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1268_ ( .A1(\us12\/_0054_ ), .A2(\us12\/_0732_ ), .B1(\us12\/_0748_ ), .B2(\us12\/_0304_ ), .Y(\us12\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1269_ ( .A(\us12\/_0477_ ), .B(\us12\/_0479_ ), .C(\us12\/_0480_ ), .D(\us12\/_0481_ ), .X(\us12\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1270_ ( .A(\us12\/_0161_ ), .B(\us12\/_0064_ ), .Y(\us12\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us12/_1271_ ( .A(\us12\/_0732_ ), .B(\us12\/_0123_ ), .C(\us12\/_0467_ ), .Y(\us12\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1272_ ( .A(\us12\/_0483_ ), .B(\us12\/_0484_ ), .Y(\us12\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1273_ ( .A(\us12\/_0297_ ), .Y(\us12\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us12/_1274_ ( .A_N(\us12\/_0485_ ), .B(\us12\/_0181_ ), .C(\us12\/_0486_ ), .D(\us12\/_0386_ ), .X(\us12\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1275_ ( .A(\us12\/_0472_ ), .B(\us12\/_0476_ ), .C(\us12\/_0482_ ), .D(\us12\/_0487_ ), .X(\us12\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \us12/_1276_ ( .A(\us12\/_0440_ ), .B(\us12\/_0462_ ), .C(\us12\/_0488_ ), .Y(\us12\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1277_ ( .A(\us12\/_0403_ ), .B(\us12\/_0230_ ), .C(\us12\/_0451_ ), .D(\us12\/_0361_ ), .X(\us12\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1278_ ( .A1(\us12\/_0118_ ), .A2(\us12\/_0050_ ), .B1(\us12\/_0109_ ), .C1(\us12\/_0139_ ), .Y(\us12\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1279_ ( .A(\us12\/_0447_ ), .B(\us12\/_0437_ ), .C(\us12\/_0491_ ), .D(\us12\/_0427_ ), .X(\us12\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1280_ ( .A1(\us12\/_0084_ ), .A2(\us12\/_0255_ ), .B1(\us12\/_0608_ ), .B2(\us12\/_0029_ ), .Y(\us12\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1281_ ( .A1(\us12\/_0144_ ), .A2(\us12\/_0147_ ), .B1(\us12\/_0355_ ), .B2(\us12\/_0093_ ), .Y(\us12\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1282_ ( .A1(\us12\/_0705_ ), .A2(\us12\/_0279_ ), .B1(\us12\/_0330_ ), .B2(\us12\/_0029_ ), .Y(\us12\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1283_ ( .A1(\us12\/_0279_ ), .A2(\us12\/_0084_ ), .B1(\us12\/_0114_ ), .Y(\us12\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1284_ ( .A(\us12\/_0493_ ), .B(\us12\/_0494_ ), .C(\us12\/_0495_ ), .D(\us12\/_0496_ ), .X(\us12\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1285_ ( .A1(\us12\/_0134_ ), .A2(\us12\/_0137_ ), .B1(\us12\/_0355_ ), .B2(\us12\/_0575_ ), .Y(\us12\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1286_ ( .A1(\us12\/_0099_ ), .A2(\us12\/_0733_ ), .B1(\us12\/_0093_ ), .B2(\us12\/_0499_ ), .Y(\us12\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1287_ ( .A(\us12\/_0147_ ), .B(\us12\/_0640_ ), .Y(\us12\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1288_ ( .A1(\us12\/_0153_ ), .A2(\us12\/_0056_ ), .B1(\us12\/_0748_ ), .Y(\us12\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1289_ ( .A(\us12\/_0498_ ), .B(\us12\/_0500_ ), .C(\us12\/_0501_ ), .D(\us12\/_0502_ ), .X(\us12\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1290_ ( .A(\us12\/_0490_ ), .B(\us12\/_0492_ ), .C(\us12\/_0497_ ), .D(\us12\/_0503_ ), .X(\us12\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us12/_1291_ ( .A_N(\us12\/_0275_ ), .B(\us12\/_0705_ ), .X(\us12\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1292_ ( .A(\us12\/_0505_ ), .Y(\us12\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1293_ ( .A(\us12\/_0380_ ), .B(\us12\/_0347_ ), .X(\us12\/_0507_ ) );
sky130_fd_sc_hd__o21ai_1 \us12/_1294_ ( .A1(\us12\/_0507_ ), .A2(\us12\/_0093_ ), .B1(\us12\/_0056_ ), .Y(\us12\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1295_ ( .A(\us12\/_0322_ ), .B(\us12\/_0277_ ), .C(\us12\/_0506_ ), .D(\us12\/_0508_ ), .X(\us12\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1296_ ( .A(\us12\/_0084_ ), .B(\us12\/_0705_ ), .X(\us12\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1297_ ( .A1(\us12\/_0733_ ), .A2(\us12\/_0114_ ), .B1(\us12\/_0429_ ), .C1(\us12\/_0511_ ), .Y(\us12\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_1298_ ( .A(\us12\/_0019_ ), .B(\us12\/_0024_ ), .Y(\us12\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1299_ ( .A(\us12\/_0512_ ), .B(\us12\/_0513_ ), .C(\us12\/_0742_ ), .D(\us12\/_0306_ ), .X(\us12\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1300_ ( .A1(\us12\/_0532_ ), .A2(\us12\/_0089_ ), .B1(\us12\/_0154_ ), .C1(\us12\/_0169_ ), .Y(\us12\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us12/_1301_ ( .A1(\us12\/_0749_ ), .A2(\us12\/_0026_ ), .B1(\us12\/_0069_ ), .C1(\us12\/_0032_ ), .X(\us12\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us12/_1302_ ( .A1(\us12\/_0324_ ), .A2(\us12\/_0355_ ), .B1(\us12\/_0330_ ), .B2(\us12\/_0727_ ), .X(\us12\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us12/_1303_ ( .A(\us12\/_0133_ ), .B(\us12\/_0516_ ), .C(\us12\/_0517_ ), .Y(\us12\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1304_ ( .A(\us12\/_0509_ ), .B(\us12\/_0514_ ), .C(\us12\/_0515_ ), .D(\us12\/_0518_ ), .X(\us12\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1305_ ( .A(\us12\/_0747_ ), .B(\us12\/_0072_ ), .Y(\us12\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1306_ ( .A1(\us12\/_0082_ ), .A2(\us12\/_0070_ ), .B1(\us12\/_0043_ ), .B2(\us12\/_0193_ ), .Y(\us12\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1307_ ( .A(\us12\/_0311_ ), .B(\us12\/_0520_ ), .C(\us12\/_0332_ ), .D(\us12\/_0522_ ), .X(\us12\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1308_ ( .A(\us12\/_0129_ ), .B(\us12\/_0499_ ), .X(\us12\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_1309_ ( .A(\us12\/_0235_ ), .B(\us12\/_0524_ ), .Y(\us12\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us12/_1310_ ( .A(\us12\/_0081_ ), .B(\us12\/_0085_ ), .Y(\us12\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1311_ ( .A1(\us12\/_0051_ ), .A2(\us12\/_0045_ ), .B1(\us12\/_0130_ ), .B2(\us12\/_0094_ ), .Y(\us12\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1312_ ( .A(\us12\/_0523_ ), .B(\us12\/_0525_ ), .C(\us12\/_0526_ ), .D(\us12\/_0527_ ), .X(\us12\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us12/_1313_ ( .A_N(\us12\/_0250_ ), .B(\us12\/_0521_ ), .Y(\us12\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1314_ ( .A(\us12\/_0128_ ), .B(\us12\/_0020_ ), .X(\us12\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1315_ ( .A(\us12\/_0530_ ), .Y(\us12\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1316_ ( .A(\us12\/_0099_ ), .B(\us12\/_0058_ ), .X(\us12\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1317_ ( .A(\us12\/_0533_ ), .Y(\us12\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us12/_1318_ ( .A_N(\us12\/_0529_ ), .B(\us12\/_0531_ ), .C(\us12\/_0534_ ), .D(\us12\/_0192_ ), .X(\us12\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1319_ ( .A(\us12\/_0434_ ), .B(\us12\/_0078_ ), .X(\us12\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us12/_1320_ ( .A1(\us12\/_0750_ ), .A2(\us12\/_0079_ ), .B1(\us12\/_0129_ ), .B2(\us12\/_0705_ ), .X(\us12\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1321_ ( .A1(\us12\/_0161_ ), .A2(\us12\/_0032_ ), .B1(\us12\/_0536_ ), .C1(\us12\/_0537_ ), .Y(\us12\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us12/_1322_ ( .A1(\us12\/_0747_ ), .A2(\us12\/_0162_ ), .B1(\us12\/_0079_ ), .B2(\us12\/_0043_ ), .X(\us12\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1323_ ( .A1(\us12\/_0093_ ), .A2(\us12\/_0029_ ), .B1(\us12\/_0240_ ), .C1(\us12\/_0539_ ), .Y(\us12\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1324_ ( .A(\us12\/_0434_ ), .B(\us12\/_0043_ ), .X(\us12\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us12/_1325_ ( .A1(\us12\/_0142_ ), .A2(\us12\/_0150_ ), .B1(\us12\/_0022_ ), .B2(\us12\/_0137_ ), .X(\us12\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1326_ ( .A1(\us12\/_0279_ ), .A2(\us12\/_0051_ ), .B1(\us12\/_0541_ ), .C1(\us12\/_0542_ ), .Y(\us12\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1327_ ( .A(\us12\/_0159_ ), .B(\us12\/_0035_ ), .X(\us12\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us12/_1328_ ( .A1(\us12\/_0271_ ), .A2(\us12\/_0434_ ), .B1(\us12\/_0027_ ), .X(\us12\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1329_ ( .A1(\us12\/_0091_ ), .A2(\us12\/_0128_ ), .B1(\us12\/_0545_ ), .C1(\us12\/_0546_ ), .Y(\us12\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1330_ ( .A(\us12\/_0538_ ), .B(\us12\/_0540_ ), .C(\us12\/_0544_ ), .D(\us12\/_0547_ ), .X(\us12\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1331_ ( .A(\us12\/_0099_ ), .B(\us12\/_0193_ ), .X(\us12\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us12/_1332_ ( .A(\us12\/_0549_ ), .B(\us12\/_0186_ ), .C(\us12\/_0187_ ), .Y(\us12\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1333_ ( .A(\us12\/_0062_ ), .B(\us12\/_0347_ ), .C(\us12\/_0749_ ), .D(\us12\/_0694_ ), .X(\us12\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1334_ ( .A1(\us12\/_0130_ ), .A2(\us12\/_0499_ ), .B1(\us12\/_0551_ ), .C1(\us12\/_0101_ ), .Y(\us12\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1335_ ( .A(\us12\/_0139_ ), .B(\us12\/_0640_ ), .Y(\us12\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1336_ ( .A1(\us12\/_0752_ ), .A2(\us12\/_0662_ ), .B1(\us12\/_0084_ ), .B2(\us12\/_0099_ ), .Y(\us12\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1337_ ( .A(\us12\/_0550_ ), .B(\us12\/_0552_ ), .C(\us12\/_0553_ ), .D(\us12\/_0555_ ), .X(\us12\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1338_ ( .A(\us12\/_0528_ ), .B(\us12\/_0535_ ), .C(\us12\/_0548_ ), .D(\us12\/_0556_ ), .X(\us12\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us12/_1339_ ( .A(\us12\/_0504_ ), .B(\us12\/_0519_ ), .C(\us12\/_0557_ ), .Y(\us12\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1340_ ( .A(\us12\/_0054_ ), .B(\us12\/_0507_ ), .X(\us12\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us12/_1341_ ( .A_N(\us12\/_0558_ ), .B(\us12\/_0408_ ), .C(\us12\/_0451_ ), .D(\us12\/_0452_ ), .X(\us12\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1342_ ( .A(\us12\/_0549_ ), .Y(\us12\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1343_ ( .A(\us12\/_0559_ ), .B(\us12\/_0403_ ), .C(\us12\/_0560_ ), .D(\us12\/_0371_ ), .X(\us12\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1344_ ( .A(\us12\/_0181_ ), .B(\us12\/_0178_ ), .X(\us12\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1345_ ( .A(\us12\/_0562_ ), .B(\us12\/_0552_ ), .C(\us12\/_0553_ ), .D(\us12\/_0555_ ), .X(\us12\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1346_ ( .A(\us12\/_0029_ ), .B(\us12\/_0020_ ), .Y(\us12\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1347_ ( .A(\us12\/_0051_ ), .B(\us12\/_0130_ ), .X(\us12\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1348_ ( .A(\us12\/_0566_ ), .Y(\us12\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1349_ ( .A(\us12\/_0159_ ), .B(\us12\/_0423_ ), .X(\us12\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1350_ ( .A1(\us12\/_0752_ ), .A2(\us12\/_0640_ ), .B1(\us12\/_0568_ ), .B2(\us12\/_0175_ ), .Y(\us12\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1351_ ( .A(\us12\/_0076_ ), .B(\us12\/_0565_ ), .C(\us12\/_0567_ ), .D(\us12\/_0569_ ), .X(\us12\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us12/_1352_ ( .A1(\us12\/_0035_ ), .A2(\us12\/_0142_ ), .B1(\us12\/_0161_ ), .X(\us12\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1353_ ( .A(\us12\/_0099_ ), .B(\us12\/_0662_ ), .Y(\us12\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us12/_1354_ ( .A(\us12\/_0420_ ), .B(\us12\/_0571_ ), .C_N(\us12\/_0572_ ), .Y(\us12\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1355_ ( .A(\us12\/_0051_ ), .B(\us12\/_0747_ ), .Y(\us12\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1356_ ( .A(\us12\/_0574_ ), .B(\us12\/_0319_ ), .C(\us12\/_0320_ ), .D(\us12\/_0411_ ), .X(\us12\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1357_ ( .A(\us12\/_0736_ ), .B(\us12\/_0035_ ), .Y(\us12\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1358_ ( .A(\us12\/_0736_ ), .B(\us12\/_0030_ ), .Y(\us12\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1359_ ( .A(\us12\/_0298_ ), .B(\us12\/_0208_ ), .C(\us12\/_0577_ ), .D(\us12\/_0578_ ), .X(\us12\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1360_ ( .A1(\us12\/_0020_ ), .A2(\us12\/_0137_ ), .B1(\us12\/_0261_ ), .B2(\us12\/_0128_ ), .Y(\us12\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1361_ ( .A(\us12\/_0573_ ), .B(\us12\/_0576_ ), .C(\us12\/_0579_ ), .D(\us12\/_0580_ ), .X(\us12\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1362_ ( .A(\us12\/_0561_ ), .B(\us12\/_0563_ ), .C(\us12\/_0570_ ), .D(\us12\/_0581_ ), .X(\us12\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1363_ ( .A(\us12\/_0128_ ), .B(\us12\/_0193_ ), .X(\us12\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1364_ ( .A(\us12\/_0082_ ), .B(\us12\/_0162_ ), .X(\us12\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us12/_1365_ ( .A(\us12\/_0583_ ), .B(\us12\/_0584_ ), .C_N(\us12\/_0437_ ), .Y(\us12\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us12/_1366_ ( .A(\us12\/_0150_ ), .B(\us12\/_0118_ ), .C(\us12\/_0380_ ), .Y(\us12\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us12/_1367_ ( .A_N(\us12\/_0182_ ), .B(\us12\/_0587_ ), .C(\us12\/_0323_ ), .X(\us12\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1368_ ( .A1(\us12\/_0575_ ), .A2(\us12\/_0153_ ), .B1(\us12\/_0727_ ), .B2(\us12\/_0058_ ), .Y(\us12\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1369_ ( .A1(\us12\/_0499_ ), .A2(\us12\/_0064_ ), .B1(\us12\/_0134_ ), .B2(\us12\/_0255_ ), .Y(\us12\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1370_ ( .A(\us12\/_0585_ ), .B(\us12\/_0588_ ), .C(\us12\/_0589_ ), .D(\us12\/_0590_ ), .X(\us12\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us12/_1371_ ( .A1(\us12\/_0091_ ), .A2(\us12\/_0139_ ), .B1(\us12\/_0250_ ), .Y(\us12\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1372_ ( .A1(\us12\/_0092_ ), .A2(\us12\/_0739_ ), .B1(\us12\/_0324_ ), .B2(\us12\/_0029_ ), .Y(\us12\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1373_ ( .A1(\us12\/_0144_ ), .A2(\us12\/_0153_ ), .B1(\us12\/_0683_ ), .B2(\us12\/_0056_ ), .Y(\us12\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1374_ ( .A1(\us12\/_0091_ ), .A2(\us12\/_0499_ ), .B1(\us12\/_0330_ ), .B2(\us12\/_0056_ ), .Y(\us12\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1375_ ( .A(\us12\/_0592_ ), .B(\us12\/_0593_ ), .C(\us12\/_0594_ ), .D(\us12\/_0595_ ), .X(\us12\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1376_ ( .A(\us12\/_0499_ ), .B(\us12\/_0144_ ), .Y(\us12\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1377_ ( .A(\us12\/_0312_ ), .B(\us12\/_0598_ ), .Y(\us12\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1378_ ( .A(\us12\/_0575_ ), .B(\us12\/_0147_ ), .Y(\us12\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1379_ ( .A1(\us12\/_0293_ ), .A2(\us12\/_0137_ ), .B1(\us12\/_0093_ ), .B2(\us12\/_0739_ ), .Y(\us12\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1380_ ( .A1(\us12\/_0734_ ), .A2(\us12\/_0531_ ), .B1(\us12\/_0600_ ), .C1(\us12\/_0601_ ), .Y(\us12\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1381_ ( .A1(\us12\/_0153_ ), .A2(\us12\/_0261_ ), .B1(\us12\/_0599_ ), .C1(\us12\/_0602_ ), .Y(\us12\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1382_ ( .A(\us12\/_0591_ ), .B(\us12\/_0596_ ), .C(\us12\/_0174_ ), .D(\us12\/_0603_ ), .X(\us12\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1383_ ( .A(\us12\/_0029_ ), .B(\us12\/_0144_ ), .Y(\us12\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1384_ ( .A(\us12\/_0113_ ), .B(\us12\/_0018_ ), .Y(\us12\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1385_ ( .A(\us12\/_0381_ ), .B(\us12\/_0605_ ), .C(\us12\/_0361_ ), .D(\us12\/_0606_ ), .X(\us12\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1386_ ( .A1(\us12\/_0016_ ), .A2(\us12\/_0727_ ), .B1(\us12\/_0733_ ), .Y(\us12\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1387_ ( .A1(\us12\/_0586_ ), .A2(\us12\/_0159_ ), .B1(\us12\/_0082_ ), .B2(\us12\/_0750_ ), .Y(\us12\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1388_ ( .A1(\us12\/_0142_ ), .A2(\us12\/_0162_ ), .B1(\us12\/_0079_ ), .B2(\us12\/_0054_ ), .Y(\us12\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1389_ ( .A(\us12\/_0610_ ), .B(\us12\/_0611_ ), .C(\us12\/_0105_ ), .D(\us12\/_0106_ ), .X(\us12\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1390_ ( .A1(\us12\/_0094_ ), .A2(\us12\/_0302_ ), .B1(\us12\/_0324_ ), .B2(\us12\/_0089_ ), .Y(\us12\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1391_ ( .A(\us12\/_0607_ ), .B(\us12\/_0609_ ), .C(\us12\/_0612_ ), .D(\us12\/_0613_ ), .X(\us12\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1392_ ( .A(\us12\/_0041_ ), .B(\us12\/_0170_ ), .X(\us12\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1393_ ( .A(\us12\/_0554_ ), .B(\us12\/_0027_ ), .X(\us12\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1394_ ( .A(\us12\/_0027_ ), .B(\us12\/_0261_ ), .Y(\us12\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us12/_1395_ ( .A_N(\us12\/_0616_ ), .B(\us12\/_0617_ ), .Y(\us12\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1396_ ( .A1(\us12\/_0147_ ), .A2(\us12\/_0302_ ), .B1(\us12\/_0342_ ), .C1(\us12\/_0618_ ), .Y(\us12\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1397_ ( .A(\us12\/_0614_ ), .B(\us12\/_0272_ ), .C(\us12\/_0615_ ), .D(\us12\/_0620_ ), .X(\us12\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us12/_1398_ ( .A(\us12\/_0582_ ), .B(\us12\/_0604_ ), .C(\us12\/_0621_ ), .Y(\us12\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1399_ ( .A1(\us12\/_0084_ ), .A2(\us12\/_0134_ ), .B1(\us12\/_0089_ ), .Y(\us12\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1400_ ( .A1(\us12\/_0144_ ), .A2(\us12\/_0608_ ), .A3(\us12\/_0330_ ), .B1(\us12\/_0089_ ), .Y(\us12\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1401_ ( .A1(\us12\/_0197_ ), .A2(\us12\/_0130_ ), .A3(\us12\/_0110_ ), .B1(\us12\/_0094_ ), .Y(\us12\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1402_ ( .A(\us12\/_0432_ ), .B(\us12\/_0622_ ), .C(\us12\/_0623_ ), .D(\us12\/_0624_ ), .X(\us12\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us12/_1403_ ( .A1(\us12\/_0554_ ), .A2(\us12\/_0018_ ), .A3(\us12\/_0022_ ), .B1(\us12\/_0161_ ), .X(\us12\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us12/_1404_ ( .A_N(\us12\/_0269_ ), .B(\us12\/_0170_ ), .X(\us12\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1405_ ( .A1(\us12\/_0109_ ), .A2(\us12\/_0064_ ), .A3(\us12\/_0733_ ), .B1(\us12\/_0355_ ), .Y(\us12\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us12/_1406_ ( .A_N(\us12\/_0626_ ), .B(\us12\/_0627_ ), .C(\us12\/_0353_ ), .D(\us12\/_0628_ ), .X(\us12\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1407_ ( .A1(\us12\/_0091_ ), .A2(\us12\/_0110_ ), .A3(\us12\/_0176_ ), .B1(\us12\/_0139_ ), .Y(\us12\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1408_ ( .A1(\us12\/_0020_ ), .A2(\us12\/_0261_ ), .B1(\us12\/_0147_ ), .Y(\us12\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1409_ ( .A(\us12\/_0631_ ), .B(\us12\/_0344_ ), .C(\us12\/_0421_ ), .D(\us12\/_0632_ ), .X(\us12\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us12/_1410_ ( .A1(\us12\/_0325_ ), .A2(\us12\/_0734_ ), .B1(\us12\/_0038_ ), .C1(\us12\/_0113_ ), .X(\us12\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1411_ ( .A1(\us12\/_0134_ ), .A2(\us12\/_0114_ ), .B1(\us12\/_0221_ ), .C1(\us12\/_0634_ ), .Y(\us12\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us12/_1412_ ( .A(\us12\/_0119_ ), .B_N(\us12\/_0111_ ), .Y(\us12\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1413_ ( .A1(\us12\/_0032_ ), .A2(\us12\/_0113_ ), .B1(\us12\/_0636_ ), .C1(\us12\/_0400_ ), .Y(\us12\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1414_ ( .A1(\us12\/_0732_ ), .A2(\us12\/_0293_ ), .A3(\us12\/_0251_ ), .B1(\us12\/_0099_ ), .Y(\us12\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1415_ ( .A(\us12\/_0189_ ), .B(\us12\/_0635_ ), .C(\us12\/_0637_ ), .D(\us12\/_0638_ ), .X(\us12\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1416_ ( .A(\us12\/_0625_ ), .B(\us12\/_0630_ ), .C(\us12\/_0633_ ), .D(\us12\/_0639_ ), .X(\us12\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1417_ ( .A(\us12\/_0747_ ), .B(\us12\/_0738_ ), .X(\us12\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1418_ ( .A(\us12\/_0736_ ), .B(\us12\/_0731_ ), .X(\us12\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us12/_1419_ ( .A_N(\us12\/_0643_ ), .B(\us12\/_0577_ ), .Y(\us12\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1420_ ( .A1(\us12\/_0084_ ), .A2(\us12\/_0739_ ), .B1(\us12\/_0642_ ), .C1(\us12\/_0644_ ), .Y(\us12\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1421_ ( .A1(\us12\/_0050_ ), .A2(\us12\/_0543_ ), .B1(\us12\/_0194_ ), .C1(\us12\/_0738_ ), .Y(\us12\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1422_ ( .A(\us12\/_0646_ ), .B(\us12\/_0232_ ), .C(\us12\/_0417_ ), .D(\us12\/_0578_ ), .X(\us12\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1423_ ( .A1(\us12\/_0064_ ), .A2(\us12\/_0733_ ), .B1(\us12\/_0727_ ), .Y(\us12\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1424_ ( .A1(\us12\/_0193_ ), .A2(\us12\/_0276_ ), .B1(\us12\/_0727_ ), .Y(\us12\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1425_ ( .A(\us12\/_0645_ ), .B(\us12\/_0647_ ), .C(\us12\/_0648_ ), .D(\us12\/_0649_ ), .X(\us12\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1426_ ( .A1(\us12\/_0325_ ), .A2(\us12\/_0734_ ), .B1(\us12\/_0038_ ), .C1(\us12\/_0029_ ), .Y(\us12\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1427_ ( .A1(\us12\/_0543_ ), .A2(\us12\/_0216_ ), .B1(\us12\/_0423_ ), .C1(\us12\/_0029_ ), .Y(\us12\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1428_ ( .A(\us12\/_0652_ ), .B(\us12\/_0653_ ), .X(\us12\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1429_ ( .A1(\us12\/_0733_ ), .A2(\us12\/_0748_ ), .A3(\us12\/_0324_ ), .B1(\us12\/_0016_ ), .Y(\us12\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1430_ ( .A1(\us12\/_0640_ ), .A2(\us12\/_0193_ ), .A3(\us12\/_0091_ ), .B1(\us12\/_0016_ ), .Y(\us12\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1431_ ( .A1(\us12\/_0102_ ), .A2(\us12\/_0301_ ), .B1(\sa12\[3\] ), .C1(\us12\/_0029_ ), .Y(\us12\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1432_ ( .A(\us12\/_0654_ ), .B(\us12\/_0655_ ), .C(\us12\/_0656_ ), .D(\us12\/_0657_ ), .X(\us12\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1433_ ( .A1(\us12\/_0118_ ), .A2(\us12\/_0050_ ), .B1(\us12\/_0038_ ), .C1(\us12\/_0489_ ), .Y(\us12\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us12/_1434_ ( .A_N(\us12\/_0250_ ), .B(\us12\/_0465_ ), .C(\us12\/_0659_ ), .X(\us12\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1435_ ( .A1(\us12\/_0683_ ), .A2(\us12\/_0324_ ), .B1(\us12\/_0255_ ), .Y(\us12\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1436_ ( .A1(\us12\/_0032_ ), .A2(\us12\/_0193_ ), .A3(\us12\/_0047_ ), .B1(\us12\/_0255_ ), .Y(\us12\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1437_ ( .A1(\us12\/_0144_ ), .A2(\us12\/_0586_ ), .A3(\us12\/_0047_ ), .B1(\us12\/_0499_ ), .Y(\us12\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1438_ ( .A(\us12\/_0660_ ), .B(\us12\/_0661_ ), .C(\us12\/_0663_ ), .D(\us12\/_0664_ ), .X(\us12\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1439_ ( .A1(\us12\/_0091_ ), .A2(\us12\/_0276_ ), .B1(\us12\/_0060_ ), .Y(\us12\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1440_ ( .A1(\us12\/_0144_ ), .A2(\us12\/_0608_ ), .B1(\us12\/_0056_ ), .Y(\us12\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1441_ ( .A1(\us12\/_0423_ ), .A2(\us12\/_0038_ ), .B1(\us12\/_0102_ ), .C1(\us12\/_0060_ ), .Y(\us12\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1442_ ( .A1(\sa12\[1\] ), .A2(\us12\/_0734_ ), .B1(\us12\/_0109_ ), .C1(\us12\/_0056_ ), .Y(\us12\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1443_ ( .A(\us12\/_0666_ ), .B(\us12\/_0667_ ), .C(\us12\/_0668_ ), .D(\us12\/_0669_ ), .X(\us12\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1444_ ( .A(\us12\/_0650_ ), .B(\us12\/_0658_ ), .C(\us12\/_0665_ ), .D(\us12\/_0670_ ), .X(\us12\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us12/_1445_ ( .A(\us12\/_0641_ ), .B(\us12\/_0174_ ), .C(\us12\/_0671_ ), .Y(\us12\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us12/_1446_ ( .A(\us12\/_0049_ ), .B(\us12\/_0618_ ), .C_N(\us12\/_0052_ ), .Y(\us12\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us12/_1447_ ( .A(\us12\/_0239_ ), .Y(\us12\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1448_ ( .A(\us12\/_0705_ ), .B(\us12\/_0032_ ), .Y(\us12\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1449_ ( .A1(\us12\/_0054_ ), .A2(\us12\/_0732_ ), .B1(\us12\/_0035_ ), .B2(\us12\/_0705_ ), .Y(\us12\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1450_ ( .A1(\us12\/_0304_ ), .A2(\us12\/_0732_ ), .B1(\us12\/_0047_ ), .B2(\us12\/_0750_ ), .Y(\us12\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1451_ ( .A(\us12\/_0674_ ), .B(\us12\/_0675_ ), .C(\us12\/_0676_ ), .D(\us12\/_0677_ ), .X(\us12\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us12/_1452_ ( .A_N(\us12\/_0584_ ), .B(\us12\/_0283_ ), .X(\us12\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1453_ ( .A(\us12\/_0673_ ), .B(\us12\/_0678_ ), .C(\us12\/_0679_ ), .D(\us12\/_0508_ ), .X(\us12\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1454_ ( .A1(\us12\/_0016_ ), .A2(\us12\/_0733_ ), .B1(\us12\/_0355_ ), .B2(\us12\/_0092_ ), .Y(\us12\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1455_ ( .A(\us12\/_0681_ ), .B(\us12\/_0034_ ), .X(\us12\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us12/_1456_ ( .A1(\us12\/_0330_ ), .A2(\us12\/_0139_ ), .B1(\us12\/_0324_ ), .B2(\us12\/_0089_ ), .X(\us12\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1457_ ( .A1(\us12\/_0146_ ), .A2(\us12\/_0147_ ), .B1(\us12\/_0133_ ), .C1(\us12\/_0684_ ), .Y(\us12\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1458_ ( .A(\us12\/_0113_ ), .B(\us12\/_0251_ ), .Y(\us12\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us12/_1459_ ( .A_N(\us12\/_0463_ ), .B(\us12\/_0686_ ), .C(\us12\/_0383_ ), .D(\us12\/_0464_ ), .X(\us12\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1460_ ( .A1(\us12\/_0051_ ), .A2(\us12\/_0293_ ), .B1(\us12\/_0084_ ), .B2(\us12\/_0705_ ), .Y(\us12\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1461_ ( .A1(\us12\/_0018_ ), .A2(\us12\/_0072_ ), .B1(\us12\/_0134_ ), .B2(\us12\/_0078_ ), .Y(\us12\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1462_ ( .A(\us12\/_0687_ ), .B(\us12\/_0236_ ), .C(\us12\/_0688_ ), .D(\us12\/_0689_ ), .X(\us12\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1463_ ( .A(\us12\/_0680_ ), .B(\us12\/_0682_ ), .C(\us12\/_0685_ ), .D(\us12\/_0690_ ), .X(\us12\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us12/_1464_ ( .A1(\us12\/_0532_ ), .A2(\us12\/_0380_ ), .B1(\us12\/_0102_ ), .C1(\us12\/_0355_ ), .X(\us12\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us12/_1465_ ( .A(\us12\/_0692_ ), .B(\us12\/_0338_ ), .C(\us12\/_0644_ ), .Y(\us12\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1466_ ( .A(\us12\/_0016_ ), .B(\us12\/_0020_ ), .Y(\us12\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1467_ ( .A1(\us12\/_0032_ ), .A2(\us12\/_0137_ ), .B1(\us12\/_0279_ ), .B2(\us12\/_0094_ ), .Y(\us12\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1468_ ( .A1(\us12\/_0575_ ), .A2(\us12\/_0153_ ), .B1(\us12\/_0161_ ), .B2(\us12\/_0293_ ), .Y(\us12\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1469_ ( .A(\us12\/_0259_ ), .B(\us12\/_0695_ ), .C(\us12\/_0696_ ), .D(\us12\/_0697_ ), .X(\us12\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us12/_1470_ ( .A1(\us12\/_0255_ ), .A2(\us12\/_0640_ ), .B1(\us12\/_0016_ ), .B2(\us12\/_0193_ ), .X(\us12\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1471_ ( .A1(\us12\/_0060_ ), .A2(\us12\/_0176_ ), .B1(\us12\/_0699_ ), .C1(\us12\/_0177_ ), .Y(\us12\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1472_ ( .A1(\us12\/_0091_ ), .A2(\us12\/_0499_ ), .B1(\us12\/_0092_ ), .B2(\us12\/_0705_ ), .Y(\us12\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us12/_1473_ ( .A1(\us12\/_0705_ ), .A2(\us12\/_0683_ ), .B1(\us12\/_0093_ ), .B2(\us12\/_0114_ ), .Y(\us12\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us12/_1474_ ( .A1(\us12\/_0683_ ), .A2(\us12\/_0084_ ), .B1(\us12\/_0094_ ), .Y(\us12\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us12/_1475_ ( .A1(\us12\/_0543_ ), .A2(\us12\/_0216_ ), .B1(\us12\/_0038_ ), .C1(\us12\/_0056_ ), .Y(\us12\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1476_ ( .A(\us12\/_0701_ ), .B(\us12\/_0702_ ), .C(\us12\/_0703_ ), .D(\us12\/_0704_ ), .X(\us12\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1477_ ( .A(\us12\/_0693_ ), .B(\us12\/_0698_ ), .C(\us12\/_0700_ ), .D(\us12\/_0706_ ), .X(\us12\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us12/_1478_ ( .A1(\us12\/_0113_ ), .A2(\us12\/_0640_ ), .B1(\us12\/_0099_ ), .B2(\us12\/_0058_ ), .X(\us12\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us12/_1479_ ( .A(\us12\/_0407_ ), .B(\us12\/_0708_ ), .C(\us12\/_0529_ ), .Y(\us12\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1480_ ( .A(\us12\/_0568_ ), .B(\us12\/_0175_ ), .Y(\us12\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us12/_1481_ ( .A1(\us12\/_0029_ ), .A2(\us12\/_0114_ ), .A3(\us12\/_0051_ ), .B1(\us12\/_0130_ ), .Y(\us12\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1482_ ( .A(\us12\/_0709_ ), .B(\us12\/_0550_ ), .C(\us12\/_0710_ ), .D(\us12\/_0711_ ), .X(\us12\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us12/_1483_ ( .A1(\us12\/_0114_ ), .A2(\us12\/_0064_ ), .B1(\us12\/_0261_ ), .B2(\us12\/_0089_ ), .X(\us12\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1484_ ( .A1(\us12\/_0355_ ), .A2(\us12\/_0261_ ), .B1(\us12\/_0198_ ), .C1(\us12\/_0713_ ), .Y(\us12\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1485_ ( .A(\us12\/_0586_ ), .B(\us12\/_0489_ ), .Y(\us12\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us12/_1486_ ( .A_N(\us12\/_0541_ ), .B(\us12\/_0267_ ), .C(\us12\/_0715_ ), .D(\us12\/_0320_ ), .X(\us12\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1487_ ( .A(\us12\/_0586_ ), .B(\us12\/_0070_ ), .Y(\us12\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us12/_1488_ ( .A_N(\us12\/_0211_ ), .B(\us12\/_0155_ ), .C(\us12\/_0202_ ), .D(\us12\/_0718_ ), .X(\us12\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us12/_1489_ ( .A(\us12\/_0150_ ), .B(\us12\/_0216_ ), .C(\us12\/_0380_ ), .Y(\us12\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us12/_1490_ ( .A(\us12\/_0411_ ), .B(\us12\/_0720_ ), .X(\us12\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us12/_1491_ ( .A1(\us12\/_0018_ ), .A2(\us12\/_0022_ ), .B1(\us12\/_0078_ ), .X(\us12\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us12/_1492_ ( .A1(\us12\/_0134_ ), .A2(\us12\/_0738_ ), .B1(\us12\/_0101_ ), .C1(\us12\/_0722_ ), .Y(\us12\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1493_ ( .A(\us12\/_0717_ ), .B(\us12\/_0719_ ), .C(\us12\/_0721_ ), .D(\us12\/_0723_ ), .X(\us12\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us12/_1494_ ( .A(\us12\/_0739_ ), .B(\us12\/_0193_ ), .Y(\us12\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1495_ ( .A(\us12\/_0344_ ), .B(\us12\/_0184_ ), .C(\us12\/_0449_ ), .D(\us12\/_0725_ ), .X(\us12\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us12/_1496_ ( .A(\us12\/_0712_ ), .B(\us12\/_0714_ ), .C(\us12\/_0724_ ), .D(\us12\/_0726_ ), .X(\us12\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \us12/_1497_ ( .A(\us12\/_0691_ ), .B(\us12\/_0707_ ), .C(\us12\/_0728_ ), .Y(\us12\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \us13/_0753_ ( .A(\sa13\[2\] ), .B_N(\sa13\[3\] ), .Y(\us13\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \us13/_0755_ ( .A(\sa13\[1\] ), .B(\sa13\[0\] ), .X(\us13\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us13/_0756_ ( .A(\us13\/_0096_ ), .B(\us13\/_0118_ ), .X(\us13\/_0129_ ) );
sky130_fd_sc_hd__and2_1 \us13/_0757_ ( .A(\sa13\[7\] ), .B(\sa13\[6\] ), .X(\us13\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_0758_ ( .A(\sa13\[4\] ), .B(\sa13\[5\] ), .Y(\us13\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0759_ ( .A(\us13\/_0140_ ), .B(\us13\/_0151_ ), .X(\us13\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0761_ ( .A(\us13\/_0129_ ), .B(\us13\/_0162_ ), .X(\us13\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0762_ ( .A(\us13\/_0096_ ), .X(\us13\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \us13/_0763_ ( .A(\sa13\[1\] ), .B_N(\sa13\[0\] ), .Y(\us13\/_0205_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0764_ ( .A(\us13\/_0205_ ), .X(\us13\/_0216_ ) );
sky130_fd_sc_hd__and3_1 \us13/_0765_ ( .A(\us13\/_0162_ ), .B(\us13\/_0194_ ), .C(\us13\/_0216_ ), .X(\us13\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us13/_0766_ ( .A(\us13\/_0183_ ), .SLEEP(\us13\/_0227_ ), .X(\us13\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \us13/_0767_ ( .A(\sa13\[0\] ), .B_N(\sa13\[1\] ), .Y(\us13\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_0768_ ( .A(\sa13\[2\] ), .B(\sa13\[3\] ), .Y(\us13\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0769_ ( .A(\us13\/_0249_ ), .B(\us13\/_0260_ ), .X(\us13\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0771_ ( .A(\us13\/_0271_ ), .X(\us13\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0772_ ( .A(\us13\/_0162_ ), .X(\us13\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_0773_ ( .A(\us13\/_0293_ ), .B(\us13\/_0304_ ), .Y(\us13\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us13/_0774_ ( .A(\sa13\[1\] ), .Y(\us13\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us13/_0776_ ( .A(\sa13\[0\] ), .Y(\us13\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0777_ ( .A(\sa13\[2\] ), .B(\sa13\[3\] ), .X(\us13\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0779_ ( .A(\us13\/_0358_ ), .X(\us13\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_0780_ ( .A1(\us13\/_0325_ ), .A2(\us13\/_0347_ ), .B1(\us13\/_0380_ ), .C1(\us13\/_0304_ ), .Y(\us13\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us13/_0781_ ( .A_N(\us13\/_0238_ ), .B(\us13\/_0314_ ), .C(\us13\/_0391_ ), .X(\us13\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us13/_0782_ ( .A(\sa13\[3\] ), .B_N(\sa13\[2\] ), .Y(\us13\/_0412_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0783_ ( .A(\us13\/_0412_ ), .X(\us13\/_0423_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0784_ ( .A(\us13\/_0423_ ), .B(\us13\/_0205_ ), .X(\us13\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \us13/_0787_ ( .A(\sa13\[5\] ), .B_N(\sa13\[4\] ), .Y(\us13\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0788_ ( .A(\us13\/_0467_ ), .B(\us13\/_0140_ ), .X(\us13\/_0478_ ) );
sky130_fd_sc_hd__buf_2 \us13/_0790_ ( .A(\us13\/_0478_ ), .X(\us13\/_0499_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_0791_ ( .A(\us13\/_0134_ ), .B(\us13\/_0499_ ), .Y(\us13\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_0792_ ( .A(\us13\/_0478_ ), .B(\us13\/_0271_ ), .Y(\us13\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0793_ ( .A(\us13\/_0194_ ), .X(\us13\/_0532_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0794_ ( .A(\us13\/_0249_ ), .X(\us13\/_0543_ ) );
sky130_fd_sc_hd__and2_1 \us13/_0795_ ( .A(\us13\/_0543_ ), .B(\us13\/_0358_ ), .X(\us13\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0797_ ( .A(\us13\/_0554_ ), .X(\us13\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us13/_0798_ ( .A(\us13\/_0216_ ), .B(\us13\/_0358_ ), .X(\us13\/_0586_ ) );
sky130_fd_sc_hd__buf_2 \us13/_0800_ ( .A(\us13\/_0586_ ), .X(\us13\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_0801_ ( .A1(\us13\/_0532_ ), .A2(\us13\/_0575_ ), .A3(\us13\/_0608_ ), .B1(\us13\/_0499_ ), .Y(\us13\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us13/_0802_ ( .A(\us13\/_0401_ ), .B(\us13\/_0510_ ), .C(\us13\/_0521_ ), .D(\us13\/_0619_ ), .X(\us13\/_0629_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0803_ ( .A(\us13\/_0358_ ), .B(\sa13\[1\] ), .X(\us13\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0805_ ( .A(\us13\/_0205_ ), .B(\us13\/_0260_ ), .X(\us13\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0807_ ( .A(\us13\/_0662_ ), .X(\us13\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us13/_0808_ ( .A(\sa13\[6\] ), .B_N(\sa13\[7\] ), .Y(\us13\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \us13/_0809_ ( .A(\us13\/_0467_ ), .B(\us13\/_0694_ ), .X(\us13\/_0705_ ) );
sky130_fd_sc_hd__buf_2 \us13/_0810_ ( .A(\us13\/_0705_ ), .X(\us13\/_0716_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0811_ ( .A(\us13\/_0716_ ), .X(\us13\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_0812_ ( .A1(\us13\/_0640_ ), .A2(\us13\/_0293_ ), .A3(\us13\/_0683_ ), .B1(\us13\/_0727_ ), .Y(\us13\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_0813_ ( .A(\sa13\[1\] ), .B(\sa13\[0\] ), .Y(\us13\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0814_ ( .A(\us13\/_0730_ ), .B(\us13\/_0260_ ), .X(\us13\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0815_ ( .A(\us13\/_0731_ ), .X(\us13\/_0732_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0816_ ( .A(\us13\/_0732_ ), .X(\us13\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0817_ ( .A(\sa13\[0\] ), .X(\us13\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us13/_0818_ ( .A1(\us13\/_0325_ ), .A2(\us13\/_0734_ ), .B1(\us13\/_0423_ ), .X(\us13\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0819_ ( .A(\us13\/_0694_ ), .B(\us13\/_0151_ ), .X(\us13\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0821_ ( .A(\us13\/_0736_ ), .X(\us13\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0822_ ( .A(\us13\/_0738_ ), .X(\us13\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_0823_ ( .A1(\us13\/_0733_ ), .A2(\us13\/_0735_ ), .A3(\us13\/_0293_ ), .B1(\us13\/_0739_ ), .Y(\us13\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us13/_0824_ ( .A(\us13\/_0730_ ), .B_N(\us13\/_0358_ ), .Y(\us13\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_0825_ ( .A(\us13\/_0741_ ), .B(\us13\/_0739_ ), .Y(\us13\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_0827_ ( .A1(\us13\/_0118_ ), .A2(\us13\/_0216_ ), .B1(\us13\/_0532_ ), .C1(\us13\/_0739_ ), .Y(\us13\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us13/_0828_ ( .A(\us13\/_0729_ ), .B(\us13\/_0740_ ), .C(\us13\/_0742_ ), .D(\us13\/_0744_ ), .X(\us13\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0829_ ( .A(\us13\/_0423_ ), .B(\us13\/_0730_ ), .X(\us13\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0830_ ( .A(\us13\/_0746_ ), .X(\us13\/_0747_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0831_ ( .A(\us13\/_0747_ ), .X(\us13\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us13/_0832_ ( .A(\sa13\[4\] ), .B_N(\sa13\[5\] ), .Y(\us13\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0833_ ( .A(\us13\/_0749_ ), .B(\us13\/_0694_ ), .X(\us13\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0835_ ( .A(\us13\/_0750_ ), .X(\us13\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0836_ ( .A(\us13\/_0752_ ), .X(\us13\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0837_ ( .A(\us13\/_0118_ ), .B(\us13\/_0358_ ), .X(\us13\/_0017_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0838_ ( .A(\us13\/_0017_ ), .X(\us13\/_0018_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0839_ ( .A(\us13\/_0752_ ), .B(\us13\/_0018_ ), .X(\us13\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0840_ ( .A(\us13\/_0358_ ), .B(\us13\/_0325_ ), .X(\us13\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0842_ ( .A(\us13\/_0096_ ), .B(\us13\/_0205_ ), .X(\us13\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \us13/_0844_ ( .A1(\us13\/_0020_ ), .A2(\us13\/_0022_ ), .B1(\us13\/_0752_ ), .X(\us13\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_0845_ ( .A1(\us13\/_0748_ ), .A2(\us13\/_0016_ ), .B1(\us13\/_0019_ ), .C1(\us13\/_0024_ ), .Y(\us13\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \us13/_0846_ ( .A(\sa13\[4\] ), .B(\sa13\[5\] ), .X(\us13\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0847_ ( .A(\us13\/_0694_ ), .B(\us13\/_0026_ ), .X(\us13\/_0027_ ) );
sky130_fd_sc_hd__buf_2 \us13/_0849_ ( .A(\us13\/_0027_ ), .X(\us13\/_0029_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0850_ ( .A(\us13\/_0358_ ), .B(\us13\/_0730_ ), .X(\us13\/_0030_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0852_ ( .A(\us13\/_0030_ ), .X(\us13\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_0853_ ( .A(\us13\/_0029_ ), .B(\us13\/_0032_ ), .Y(\us13\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_0854_ ( .A(\us13\/_0029_ ), .B(\us13\/_0735_ ), .Y(\us13\/_0034_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0855_ ( .A(\us13\/_0118_ ), .B(\us13\/_0260_ ), .X(\us13\/_0035_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0856_ ( .A(\us13\/_0035_ ), .X(\us13\/_0036_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0857_ ( .A(\us13\/_0027_ ), .B(\us13\/_0036_ ), .X(\us13\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0858_ ( .A(\us13\/_0260_ ), .X(\us13\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_0859_ ( .A(\us13\/_0038_ ), .B(\us13\/_0347_ ), .Y(\us13\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us13/_0860_ ( .A_N(\us13\/_0039_ ), .B(\us13\/_0027_ ), .X(\us13\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_0861_ ( .A(\us13\/_0037_ ), .B(\us13\/_0040_ ), .Y(\us13\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us13/_0862_ ( .A(\us13\/_0025_ ), .B(\us13\/_0033_ ), .C(\us13\/_0034_ ), .D(\us13\/_0041_ ), .X(\us13\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0863_ ( .A(\us13\/_0749_ ), .B(\us13\/_0140_ ), .X(\us13\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us13/_0865_ ( .A(\sa13\[0\] ), .B(\sa13\[2\] ), .C(\sa13\[3\] ), .X(\us13\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0866_ ( .A(\us13\/_0043_ ), .B(\us13\/_0045_ ), .X(\us13\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0867_ ( .A(\us13\/_0096_ ), .B(\us13\/_0543_ ), .X(\us13\/_0047_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0868_ ( .A(\us13\/_0047_ ), .X(\us13\/_0048_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0869_ ( .A(\us13\/_0048_ ), .B(\us13\/_0043_ ), .X(\us13\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0870_ ( .A(\us13\/_0730_ ), .X(\us13\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0871_ ( .A(\us13\/_0043_ ), .X(\us13\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_0872_ ( .A1(\us13\/_0118_ ), .A2(\us13\/_0050_ ), .B1(\us13\/_0194_ ), .C1(\us13\/_0051_ ), .Y(\us13\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us13/_0873_ ( .A(\us13\/_0046_ ), .B(\us13\/_0049_ ), .C_N(\us13\/_0052_ ), .Y(\us13\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0874_ ( .A(\us13\/_0026_ ), .B(\us13\/_0140_ ), .X(\us13\/_0054_ ) );
sky130_fd_sc_hd__buf_2 \us13/_0876_ ( .A(\us13\/_0054_ ), .X(\us13\/_0056_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_0877_ ( .A1(\us13\/_0532_ ), .A2(\us13\/_0575_ ), .B1(\us13\/_0056_ ), .Y(\us13\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0878_ ( .A(\us13\/_0423_ ), .B(\us13\/_0325_ ), .X(\us13\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0880_ ( .A(\us13\/_0051_ ), .X(\us13\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_0881_ ( .A1(\us13\/_0732_ ), .A2(\us13\/_0036_ ), .A3(\us13\/_0058_ ), .B1(\us13\/_0060_ ), .Y(\us13\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0882_ ( .A(\us13\/_0260_ ), .B(\sa13\[1\] ), .X(\us13\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0884_ ( .A(\us13\/_0062_ ), .X(\us13\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_0885_ ( .A1(\us13\/_0064_ ), .A2(\us13\/_0748_ ), .A3(\us13\/_0683_ ), .B1(\us13\/_0056_ ), .Y(\us13\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us13/_0886_ ( .A(\us13\/_0053_ ), .B(\us13\/_0057_ ), .C(\us13\/_0061_ ), .D(\us13\/_0065_ ), .X(\us13\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us13/_0887_ ( .A(\us13\/_0629_ ), .B(\us13\/_0745_ ), .C(\us13\/_0042_ ), .D(\us13\/_0066_ ), .X(\us13\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us13/_0889_ ( .A(\sa13\[7\] ), .B_N(\sa13\[6\] ), .Y(\us13\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0890_ ( .A(\us13\/_0069_ ), .B(\us13\/_0151_ ), .X(\us13\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0892_ ( .A(\us13\/_0070_ ), .X(\us13\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_0893_ ( .A1(\us13\/_0129_ ), .A2(\us13\/_0586_ ), .B1(\us13\/_0072_ ), .Y(\us13\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_0894_ ( .A1(\us13\/_0380_ ), .A2(\us13\/_0347_ ), .B1(\us13\/_0194_ ), .B2(\us13\/_0216_ ), .Y(\us13\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us13/_0895_ ( .A(\us13\/_0074_ ), .B_N(\us13\/_0070_ ), .Y(\us13\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us13/_0896_ ( .A(\us13\/_0073_ ), .SLEEP(\us13\/_0075_ ), .X(\us13\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us13/_0897_ ( .A(\us13\/_0467_ ), .B(\us13\/_0069_ ), .X(\us13\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0898_ ( .A(\us13\/_0077_ ), .X(\us13\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0899_ ( .A(\us13\/_0412_ ), .B(\us13\/_0118_ ), .X(\us13\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0901_ ( .A(\us13\/_0078_ ), .B(\us13\/_0079_ ), .X(\us13\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0902_ ( .A(\us13\/_0412_ ), .B(\us13\/_0249_ ), .X(\us13\/_0082_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0903_ ( .A(\us13\/_0082_ ), .X(\us13\/_0083_ ) );
sky130_fd_sc_hd__buf_2 \us13/_0904_ ( .A(\us13\/_0083_ ), .X(\us13\/_0084_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0905_ ( .A(\us13\/_0084_ ), .B(\us13\/_0078_ ), .X(\us13\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us13/_0906_ ( .A1(\sa13\[0\] ), .A2(\us13\/_0325_ ), .B1(\us13\/_0260_ ), .Y(\us13\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us13/_0907_ ( .A_N(\us13\/_0086_ ), .B(\us13\/_0078_ ), .X(\us13\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us13/_0908_ ( .A(\us13\/_0081_ ), .B(\us13\/_0085_ ), .C(\us13\/_0087_ ), .Y(\us13\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0909_ ( .A(\us13\/_0072_ ), .X(\us13\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_0910_ ( .A1(\us13\/_0733_ ), .A2(\us13\/_0748_ ), .A3(\us13\/_0683_ ), .B1(\us13\/_0089_ ), .Y(\us13\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0911_ ( .A(\us13\/_0129_ ), .X(\us13\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0912_ ( .A(\us13\/_0018_ ), .X(\us13\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0913_ ( .A(\us13\/_0022_ ), .X(\us13\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0914_ ( .A(\us13\/_0078_ ), .X(\us13\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_0915_ ( .A1(\us13\/_0091_ ), .A2(\us13\/_0092_ ), .A3(\us13\/_0093_ ), .B1(\us13\/_0094_ ), .Y(\us13\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us13/_0916_ ( .A(\us13\/_0076_ ), .B(\us13\/_0088_ ), .C(\us13\/_0090_ ), .D(\us13\/_0095_ ), .X(\us13\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us13/_0917_ ( .A(\us13\/_0069_ ), .B(\us13\/_0026_ ), .X(\us13\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \us13/_0918_ ( .A(\us13\/_0098_ ), .X(\us13\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0919_ ( .A(\us13\/_0434_ ), .B(\us13\/_0099_ ), .X(\us13\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0920_ ( .A(\us13\/_0079_ ), .B(\us13\/_0098_ ), .X(\us13\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0921_ ( .A(\us13\/_0325_ ), .X(\us13\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_0922_ ( .A1(\us13\/_0102_ ), .A2(\us13\/_0734_ ), .B1(\us13\/_0038_ ), .C1(\us13\/_0099_ ), .Y(\us13\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us13/_0923_ ( .A(\us13\/_0100_ ), .B(\us13\/_0101_ ), .C_N(\us13\/_0103_ ), .Y(\us13\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_0924_ ( .A1(\us13\/_0554_ ), .A2(\us13\/_0586_ ), .B1(\us13\/_0099_ ), .Y(\us13\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_0925_ ( .A(\us13\/_0129_ ), .B(\us13\/_0099_ ), .Y(\us13\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0926_ ( .A(\us13\/_0105_ ), .B(\us13\/_0106_ ), .X(\us13\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0927_ ( .A(\us13\/_0423_ ), .X(\us13\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us13/_0928_ ( .A(\us13\/_0260_ ), .B(\sa13\[0\] ), .X(\us13\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0929_ ( .A(\us13\/_0069_ ), .B(\us13\/_0749_ ), .X(\us13\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0931_ ( .A(\us13\/_0111_ ), .X(\us13\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0932_ ( .A(\us13\/_0113_ ), .X(\us13\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_0933_ ( .A1(\us13\/_0109_ ), .A2(\us13\/_0110_ ), .B1(\us13\/_0114_ ), .Y(\us13\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us13/_0934_ ( .A(\us13\/_0022_ ), .Y(\us13\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us13/_0935_ ( .A(\us13\/_0554_ ), .Y(\us13\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us13/_0936_ ( .A1(\us13\/_0050_ ), .A2(\us13\/_0118_ ), .B1(\us13\/_0194_ ), .Y(\us13\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us13/_0937_ ( .A(\us13\/_0113_ ), .Y(\us13\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us13/_0938_ ( .A1(\us13\/_0116_ ), .A2(\us13\/_0117_ ), .A3(\us13\/_0119_ ), .B1(\us13\/_0120_ ), .X(\us13\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us13/_0939_ ( .A(\us13\/_0104_ ), .B(\us13\/_0108_ ), .C(\us13\/_0115_ ), .D(\us13\/_0121_ ), .X(\us13\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_0940_ ( .A(\sa13\[7\] ), .B(\sa13\[6\] ), .Y(\us13\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0941_ ( .A(\us13\/_0749_ ), .B(\us13\/_0123_ ), .X(\us13\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0943_ ( .A(\us13\/_0083_ ), .B(\us13\/_0124_ ), .X(\us13\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_0944_ ( .A(\us13\/_0271_ ), .B(\us13\/_0124_ ), .Y(\us13\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0945_ ( .A(\us13\/_0124_ ), .X(\us13\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0946_ ( .A(\us13\/_0260_ ), .B(\us13\/_0325_ ), .X(\us13\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_0948_ ( .A(\us13\/_0128_ ), .B(\us13\/_0130_ ), .Y(\us13\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_0949_ ( .A(\us13\/_0127_ ), .B(\us13\/_0132_ ), .Y(\us13\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us13/_0950_ ( .A(\us13\/_0434_ ), .X(\us13\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_0951_ ( .A(\us13\/_0134_ ), .B(\us13\/_0128_ ), .Y(\us13\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us13/_0952_ ( .A(\us13\/_0126_ ), .B(\us13\/_0133_ ), .C_N(\us13\/_0135_ ), .Y(\us13\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us13/_0953_ ( .A(\us13\/_0026_ ), .B(\us13\/_0123_ ), .X(\us13\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0955_ ( .A(\us13\/_0137_ ), .X(\us13\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_0956_ ( .A1(\us13\/_0110_ ), .A2(\us13\/_0293_ ), .A3(\us13\/_0084_ ), .B1(\us13\/_0139_ ), .Y(\us13\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0957_ ( .A(\us13\/_0096_ ), .B(\us13\/_0730_ ), .X(\us13\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0959_ ( .A(\us13\/_0142_ ), .X(\us13\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_0960_ ( .A1(\us13\/_0020_ ), .A2(\us13\/_0144_ ), .A3(\us13\/_0018_ ), .B1(\us13\/_0139_ ), .Y(\us13\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \us13/_0961_ ( .A(\sa13\[2\] ), .B(\us13\/_0050_ ), .C_N(\sa13\[3\] ), .Y(\us13\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0962_ ( .A(\us13\/_0128_ ), .X(\us13\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_0963_ ( .A1(\us13\/_0146_ ), .A2(\us13\/_0032_ ), .A3(\us13\/_0640_ ), .B1(\us13\/_0147_ ), .Y(\us13\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us13/_0964_ ( .A(\us13\/_0136_ ), .B(\us13\/_0141_ ), .C(\us13\/_0145_ ), .D(\us13\/_0148_ ), .X(\us13\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0965_ ( .A(\us13\/_0123_ ), .B(\us13\/_0151_ ), .X(\us13\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0967_ ( .A(\us13\/_0150_ ), .X(\us13\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \us13/_0968_ ( .A(\us13\/_0150_ ), .B(\us13\/_0062_ ), .X(\us13\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_0969_ ( .A(\us13\/_0079_ ), .B(\us13\/_0150_ ), .Y(\us13\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us13/_0970_ ( .A(\us13\/_0150_ ), .B(\us13\/_0423_ ), .C(\us13\/_0543_ ), .Y(\us13\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_0971_ ( .A(\us13\/_0155_ ), .B(\us13\/_0156_ ), .Y(\us13\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_0972_ ( .A1(\us13\/_0153_ ), .A2(\us13\/_0134_ ), .B1(\us13\/_0154_ ), .C1(\us13\/_0157_ ), .Y(\us13\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0973_ ( .A(\us13\/_0467_ ), .B(\us13\/_0123_ ), .X(\us13\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_0975_ ( .A(\us13\/_0159_ ), .X(\us13\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us13/_0976_ ( .A_N(\us13\/_0119_ ), .B(\us13\/_0161_ ), .X(\us13\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us13/_0977_ ( .A(\us13\/_0163_ ), .Y(\us13\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_0978_ ( .A1(\us13\/_0146_ ), .A2(\us13\/_0575_ ), .A3(\us13\/_0608_ ), .B1(\us13\/_0153_ ), .Y(\us13\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_0979_ ( .A1(\us13\/_0062_ ), .A2(\us13\/_0084_ ), .A3(\us13\/_0134_ ), .B1(\us13\/_0161_ ), .Y(\us13\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us13/_0980_ ( .A(\us13\/_0158_ ), .B(\us13\/_0164_ ), .C(\us13\/_0165_ ), .D(\us13\/_0166_ ), .X(\us13\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us13/_0981_ ( .A(\us13\/_0097_ ), .B(\us13\/_0122_ ), .C(\us13\/_0149_ ), .D(\us13\/_0167_ ), .X(\us13\/_0168_ ) );
sky130_fd_sc_hd__and2_1 \us13/_0982_ ( .A(\us13\/_0662_ ), .B(\us13\/_0150_ ), .X(\us13\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_0983_ ( .A(\us13\/_0154_ ), .B(\us13\/_0169_ ), .Y(\us13\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us13/_0984_ ( .A(\us13\/_0123_ ), .B(\us13\/_0151_ ), .C(\us13\/_0038_ ), .X(\us13\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0985_ ( .A(\us13\/_0170_ ), .B(\us13\/_0171_ ), .X(\us13\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \us13/_0986_ ( .A(\us13\/_0172_ ), .Y(\us13\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \us13/_0987_ ( .A(\us13\/_0067_ ), .B(\us13\/_0168_ ), .C(\us13\/_0174_ ), .Y(\us13\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us13/_0988_ ( .A(\sa13\[1\] ), .B(\sa13\[0\] ), .Y(\us13\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us13/_0989_ ( .A(\us13\/_0175_ ), .B(\us13\/_0358_ ), .X(\us13\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0990_ ( .A(\us13\/_0176_ ), .B(\us13\/_0478_ ), .X(\us13\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_0991_ ( .A(\us13\/_0084_ ), .B(\us13\/_0113_ ), .Y(\us13\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0992_ ( .A(\us13\/_0111_ ), .B(\us13\/_0062_ ), .X(\us13\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0993_ ( .A(\us13\/_0111_ ), .B(\us13\/_0662_ ), .X(\us13\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_0994_ ( .A(\us13\/_0179_ ), .B(\us13\/_0180_ ), .Y(\us13\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0995_ ( .A(\us13\/_0054_ ), .B(\us13\/_0058_ ), .X(\us13\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us13/_0996_ ( .A(\us13\/_0182_ ), .Y(\us13\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us13/_0997_ ( .A_N(\us13\/_0177_ ), .B(\us13\/_0178_ ), .C(\us13\/_0181_ ), .D(\us13\/_0184_ ), .X(\us13\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0998_ ( .A(\us13\/_0098_ ), .B(\us13\/_0741_ ), .X(\us13\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us13/_0999_ ( .A(\us13\/_0047_ ), .B(\us13\/_0098_ ), .X(\us13\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us13/_1000_ ( .A(\us13\/_0186_ ), .B(\us13\/_0187_ ), .X(\us13\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1001_ ( .A(\us13\/_0188_ ), .Y(\us13\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1002_ ( .A(\us13\/_0738_ ), .B(\us13\/_0735_ ), .X(\us13\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1003_ ( .A(\us13\/_0271_ ), .B(\us13\/_0736_ ), .X(\us13\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_1004_ ( .A(\us13\/_0190_ ), .B(\us13\/_0191_ ), .Y(\us13\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us13/_1005_ ( .A(\us13\/_0096_ ), .B(\us13\/_0325_ ), .X(\us13\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1006_ ( .A1(\us13\/_0193_ ), .A2(\us13\/_0176_ ), .B1(\us13\/_0043_ ), .Y(\us13\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1007_ ( .A(\us13\/_0185_ ), .B(\us13\/_0189_ ), .C(\us13\/_0192_ ), .D(\us13\/_0195_ ), .X(\us13\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us13/_1008_ ( .A_N(\sa13\[3\] ), .B(\us13\/_0734_ ), .C(\sa13\[2\] ), .X(\us13\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1009_ ( .A(\us13\/_0137_ ), .B(\us13\/_0197_ ), .X(\us13\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_1010_ ( .A(\us13\/_0198_ ), .B(\us13\/_0040_ ), .Y(\us13\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1011_ ( .A(\us13\/_0293_ ), .B(\us13\/_0137_ ), .X(\us13\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1012_ ( .A(\us13\/_0200_ ), .Y(\us13\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1013_ ( .A(\us13\/_0137_ ), .B(\us13\/_0110_ ), .Y(\us13\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1014_ ( .A(\us13\/_0139_ ), .B(\us13\/_0020_ ), .Y(\us13\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1015_ ( .A(\us13\/_0199_ ), .B(\us13\/_0201_ ), .C(\us13\/_0202_ ), .D(\us13\/_0203_ ), .X(\us13\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us13/_1016_ ( .A1(\us13\/_0532_ ), .A2(\us13\/_0109_ ), .B1(\us13\/_0102_ ), .C1(\us13\/_0727_ ), .X(\us13\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1017_ ( .A(\us13\/_0022_ ), .B(\us13\/_0078_ ), .Y(\us13\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1018_ ( .A(\us13\/_0078_ ), .B(\us13\/_0142_ ), .Y(\us13\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1019_ ( .A(\us13\/_0207_ ), .B(\us13\/_0208_ ), .Y(\us13\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1020_ ( .A1(\us13\/_0094_ ), .A2(\us13\/_0176_ ), .B1(\us13\/_0206_ ), .C1(\us13\/_0209_ ), .Y(\us13\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1021_ ( .A(\us13\/_0662_ ), .B(\us13\/_0070_ ), .X(\us13\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us13/_1022_ ( .A(\us13\/_0732_ ), .B(\us13\/_0123_ ), .C(\us13\/_0749_ ), .Y(\us13\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us13/_1023_ ( .A(\us13\/_0732_ ), .B(\us13\/_0467_ ), .C(\us13\/_0069_ ), .Y(\us13\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us13/_1024_ ( .A_N(\us13\/_0211_ ), .B(\us13\/_0127_ ), .C(\us13\/_0212_ ), .D(\us13\/_0213_ ), .X(\us13\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1025_ ( .A(\us13\/_0137_ ), .Y(\us13\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1026_ ( .A(\us13\/_0128_ ), .B(\us13\/_0036_ ), .Y(\us13\/_0217_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1028_ ( .A1(\us13\/_0159_ ), .A2(\us13\/_0747_ ), .B1(\us13\/_0434_ ), .B2(\us13\/_0499_ ), .Y(\us13\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us13/_1029_ ( .A1(\us13\/_0116_ ), .A2(\us13\/_0215_ ), .B1(\us13\/_0217_ ), .C1(\us13\/_0219_ ), .X(\us13\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1030_ ( .A(\us13\/_0113_ ), .B(\us13\/_0746_ ), .X(\us13\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us13/_1031_ ( .A1(\us13\/_0098_ ), .A2(\us13\/_0746_ ), .B1(\us13\/_0434_ ), .B2(\us13\/_0750_ ), .X(\us13\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1032_ ( .A1(\us13\/_0048_ ), .A2(\us13\/_0113_ ), .B1(\us13\/_0221_ ), .C1(\us13\/_0222_ ), .Y(\us13\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us13/_1033_ ( .A1(\us13\/_0129_ ), .A2(\us13\/_0162_ ), .B1(\us13\/_0271_ ), .B2(\us13\/_0705_ ), .X(\us13\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1034_ ( .A1(\us13\/_0093_ ), .A2(\us13\/_0738_ ), .B1(\us13\/_0081_ ), .C1(\us13\/_0224_ ), .Y(\us13\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1035_ ( .A(\us13\/_0214_ ), .B(\us13\/_0220_ ), .C(\us13\/_0223_ ), .D(\us13\/_0225_ ), .X(\us13\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1036_ ( .A(\us13\/_0196_ ), .B(\us13\/_0204_ ), .C(\us13\/_0210_ ), .D(\us13\/_0226_ ), .X(\us13\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1037_ ( .A(\us13\/_0111_ ), .B(\us13\/_0554_ ), .X(\us13\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1038_ ( .A(\us13\/_0229_ ), .Y(\us13\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1039_ ( .A(\us13\/_0111_ ), .B(\us13\/_0129_ ), .Y(\us13\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1040_ ( .A(\us13\/_0018_ ), .B(\us13\/_0738_ ), .Y(\us13\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1041_ ( .A(\us13\/_0030_ ), .B(\us13\/_0304_ ), .Y(\us13\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1042_ ( .A(\us13\/_0230_ ), .B(\us13\/_0231_ ), .C(\us13\/_0232_ ), .D(\us13\/_0233_ ), .X(\us13\/_0234_ ) );
sky130_fd_sc_hd__and2_1 \us13/_1043_ ( .A(\us13\/_0048_ ), .B(\us13\/_0478_ ), .X(\us13\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1044_ ( .A1(\us13\/_0129_ ), .A2(\us13\/_0554_ ), .B1(\us13\/_0137_ ), .Y(\us13\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us13/_1045_ ( .A(\us13\/_0235_ ), .B(\us13\/_0049_ ), .C_N(\us13\/_0236_ ), .Y(\us13\/_0237_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1046_ ( .A(\us13\/_0047_ ), .B(\us13\/_0077_ ), .X(\us13\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1047_ ( .A(\us13\/_0070_ ), .B(\us13\/_0036_ ), .X(\us13\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us13/_1048_ ( .A1(\us13\/_0048_ ), .A2(\us13\/_0736_ ), .B1(\us13\/_0022_ ), .B2(\us13\/_0099_ ), .X(\us13\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us13/_1049_ ( .A(\us13\/_0239_ ), .B(\us13\/_0240_ ), .C(\us13\/_0241_ ), .Y(\us13\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1050_ ( .A(\us13\/_0554_ ), .B(\us13\/_0072_ ), .X(\us13\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us13/_1051_ ( .A1(\us13\/_0142_ ), .A2(\us13\/_0137_ ), .B1(\us13\/_0159_ ), .B2(\us13\/_0083_ ), .X(\us13\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1052_ ( .A1(\us13\/_0608_ ), .A2(\us13\/_0072_ ), .B1(\us13\/_0243_ ), .C1(\us13\/_0244_ ), .Y(\us13\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1053_ ( .A(\us13\/_0234_ ), .B(\us13\/_0237_ ), .C(\us13\/_0242_ ), .D(\us13\/_0245_ ), .X(\us13\/_0246_ ) );
sky130_fd_sc_hd__o21a_1 \us13/_1055_ ( .A1(\us13\/_0554_ ), .A2(\us13\/_0586_ ), .B1(\us13\/_0029_ ), .X(\us13\/_0248_ ) );
sky130_fd_sc_hd__and2_1 \us13/_1056_ ( .A(\us13\/_0083_ ), .B(\us13\/_0478_ ), .X(\us13\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_1057_ ( .A(\us13\/_0079_ ), .X(\us13\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1058_ ( .A(\us13\/_0251_ ), .B(\us13\/_0478_ ), .X(\us13\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_1059_ ( .A(\us13\/_0250_ ), .B(\us13\/_0252_ ), .Y(\us13\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1060_ ( .A(\us13\/_0016_ ), .B(\us13\/_0064_ ), .Y(\us13\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_1061_ ( .A(\us13\/_0304_ ), .X(\us13\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1062_ ( .A(\us13\/_0255_ ), .B(\us13\/_0640_ ), .Y(\us13\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us13/_1063_ ( .A_N(\us13\/_0248_ ), .B(\us13\/_0253_ ), .C(\us13\/_0254_ ), .D(\us13\/_0256_ ), .X(\us13\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1064_ ( .A(\us13\/_0099_ ), .B(\us13\/_0110_ ), .X(\us13\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us13/_1065_ ( .A1(\us13\/_0161_ ), .A2(\us13\/_0130_ ), .B1(\us13\/_0258_ ), .Y(\us13\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1066_ ( .A(\us13\/_0194_ ), .B(\sa13\[1\] ), .X(\us13\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1068_ ( .A(\us13\/_0261_ ), .B(\us13\/_0153_ ), .Y(\us13\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us13/_1069_ ( .A_N(\us13\/_0154_ ), .B(\us13\/_0259_ ), .C(\us13\/_0263_ ), .X(\us13\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1070_ ( .A(\us13\/_0246_ ), .B(\us13\/_0174_ ), .C(\us13\/_0257_ ), .D(\us13\/_0264_ ), .X(\us13\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us13/_1071_ ( .A1(\us13\/_0261_ ), .A2(\us13\/_0554_ ), .B1(\us13\/_0159_ ), .X(\us13\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1072_ ( .A(\us13\/_0747_ ), .B(\us13\/_0150_ ), .Y(\us13\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1073_ ( .A(\us13\/_0175_ ), .Y(\us13\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us13/_1074_ ( .A(\us13\/_0423_ ), .B(\us13\/_0123_ ), .C(\us13\/_0151_ ), .X(\us13\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1075_ ( .A(\us13\/_0268_ ), .B(\us13\/_0269_ ), .Y(\us13\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us13/_1076_ ( .A_N(\us13\/_0266_ ), .B(\us13\/_0267_ ), .C(\us13\/_0270_ ), .X(\us13\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1077_ ( .A(\us13\/_0554_ ), .B(\us13\/_0150_ ), .X(\us13\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1078_ ( .A(\us13\/_0273_ ), .Y(\us13\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1079_ ( .A1(\us13\/_0734_ ), .A2(\us13\/_0325_ ), .B1(\us13\/_0380_ ), .Y(\us13\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1080_ ( .A(\us13\/_0275_ ), .Y(\us13\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1081_ ( .A(\us13\/_0276_ ), .B(\us13\/_0153_ ), .Y(\us13\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us13/_1082_ ( .A(\us13\/_0272_ ), .B(\us13\/_0274_ ), .C(\us13\/_0277_ ), .X(\us13\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_1083_ ( .A(\us13\/_0036_ ), .X(\us13\/_0279_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1085_ ( .A1(\us13\/_0499_ ), .A2(\us13\/_0279_ ), .B1(\us13\/_0084_ ), .B2(\us13\/_0060_ ), .Y(\us13\/_0281_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1086_ ( .A1(\us13\/_0251_ ), .A2(\us13\/_0434_ ), .B1(\us13\/_0304_ ), .Y(\us13\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1087_ ( .A(\us13\/_0091_ ), .B(\us13\/_0056_ ), .Y(\us13\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1088_ ( .A1(\us13\/_0118_ ), .A2(\us13\/_0050_ ), .B1(\us13\/_0038_ ), .C1(\us13\/_0255_ ), .Y(\us13\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1089_ ( .A(\us13\/_0281_ ), .B(\us13\/_0283_ ), .C(\us13\/_0284_ ), .D(\us13\/_0285_ ), .X(\us13\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1090_ ( .A(\us13\/_0083_ ), .B(\us13\/_0027_ ), .X(\us13\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1091_ ( .A(\us13\/_0129_ ), .B(\us13\/_0027_ ), .X(\us13\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_1092_ ( .A(\us13\/_0287_ ), .B(\us13\/_0288_ ), .Y(\us13\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1093_ ( .A1(\us13\/_0752_ ), .A2(\us13\/_0683_ ), .B1(\us13\/_0093_ ), .B2(\us13\/_0029_ ), .Y(\us13\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1094_ ( .A1(\us13\/_0092_ ), .A2(\us13\/_0575_ ), .B1(\us13\/_0056_ ), .Y(\us13\/_0291_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1096_ ( .A1(\us13\/_0499_ ), .A2(\us13\/_0662_ ), .B1(\us13\/_0084_ ), .B2(\us13\/_0056_ ), .Y(\us13\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1097_ ( .A(\us13\/_0289_ ), .B(\us13\/_0290_ ), .C(\us13\/_0291_ ), .D(\us13\/_0294_ ), .X(\us13\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1098_ ( .A(\us13\/_0750_ ), .B(\us13\/_0193_ ), .X(\us13\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1099_ ( .A(\us13\/_0716_ ), .B(\us13\/_0380_ ), .X(\us13\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1100_ ( .A(\us13\/_0752_ ), .B(\us13\/_0129_ ), .Y(\us13\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us13/_1101_ ( .A(\us13\/_0296_ ), .B(\us13\/_0297_ ), .C_N(\us13\/_0298_ ), .Y(\us13\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1102_ ( .A(\us13\/_0089_ ), .B(\us13\/_0532_ ), .Y(\us13\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1103_ ( .A(\sa13\[2\] ), .Y(\us13\/_0301_ ) );
sky130_fd_sc_hd__nor3_2 \us13/_1104_ ( .A(\us13\/_0301_ ), .B(\sa13\[3\] ), .C(\us13\/_0118_ ), .Y(\us13\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1105_ ( .A(\us13\/_0072_ ), .B(\us13\/_0302_ ), .X(\us13\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1106_ ( .A(\us13\/_0303_ ), .Y(\us13\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1107_ ( .A(\us13\/_0147_ ), .B(\us13\/_0302_ ), .Y(\us13\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1108_ ( .A(\us13\/_0299_ ), .B(\us13\/_0300_ ), .C(\us13\/_0305_ ), .D(\us13\/_0306_ ), .X(\us13\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1109_ ( .A(\us13\/_0278_ ), .B(\us13\/_0286_ ), .C(\us13\/_0295_ ), .D(\us13\/_0307_ ), .X(\us13\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us13/_1110_ ( .A(\us13\/_0228_ ), .B(\us13\/_0265_ ), .C(\us13\/_0308_ ), .Y(\us13\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1111_ ( .A(\us13\/_0235_ ), .Y(\us13\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1112_ ( .A(\us13\/_0478_ ), .B(\us13\/_0640_ ), .X(\us13\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1113_ ( .A(\us13\/_0310_ ), .Y(\us13\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1114_ ( .A(\us13\/_0022_ ), .B(\us13\/_0499_ ), .Y(\us13\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1115_ ( .A(\us13\/_0499_ ), .B(\us13\/_0032_ ), .Y(\us13\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1116_ ( .A(\us13\/_0309_ ), .B(\us13\/_0311_ ), .C(\us13\/_0312_ ), .D(\us13\/_0313_ ), .X(\us13\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1117_ ( .A(\us13\/_0499_ ), .B(\us13\/_0064_ ), .Y(\us13\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1118_ ( .A(\us13\/_0499_ ), .B(\us13\/_0683_ ), .Y(\us13\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1119_ ( .A(\us13\/_0315_ ), .B(\us13\/_0316_ ), .C(\us13\/_0317_ ), .D(\us13\/_0253_ ), .X(\us13\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1120_ ( .A(\us13\/_0048_ ), .B(\us13\/_0304_ ), .Y(\us13\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1121_ ( .A(\us13\/_0586_ ), .B(\us13\/_0162_ ), .Y(\us13\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1122_ ( .A(\us13\/_0319_ ), .B(\us13\/_0320_ ), .Y(\us13\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_1123_ ( .A(\us13\/_0321_ ), .B(\us13\/_0238_ ), .Y(\us13\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1124_ ( .A(\us13\/_0304_ ), .B(\us13\/_0062_ ), .Y(\us13\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_1125_ ( .A(\us13\/_0251_ ), .X(\us13\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1126_ ( .A1(\us13\/_0324_ ), .A2(\us13\/_0084_ ), .B1(\us13\/_0255_ ), .Y(\us13\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1127_ ( .A1(\us13\/_0050_ ), .A2(\us13\/_0216_ ), .B1(\us13\/_0109_ ), .C1(\us13\/_0255_ ), .Y(\us13\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1128_ ( .A(\us13\/_0322_ ), .B(\us13\/_0323_ ), .C(\us13\/_0326_ ), .D(\us13\/_0327_ ), .X(\us13\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1129_ ( .A1(\us13\/_0733_ ), .A2(\us13\/_0279_ ), .A3(\us13\/_0058_ ), .B1(\us13\/_0056_ ), .Y(\us13\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_1130_ ( .A(\us13\/_0048_ ), .X(\us13\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1131_ ( .A(\us13\/_0330_ ), .B(\us13\/_0056_ ), .Y(\us13\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1132_ ( .A(\us13\/_0054_ ), .B(\us13\/_0045_ ), .Y(\us13\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1133_ ( .A(\us13\/_0329_ ), .B(\us13\/_0331_ ), .C(\us13\/_0284_ ), .D(\us13\/_0332_ ), .X(\us13\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us13/_1134_ ( .A1(\us13\/_0543_ ), .A2(\us13\/_0216_ ), .B1(\us13\/_0532_ ), .C1(\us13\/_0060_ ), .X(\us13\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1135_ ( .A(\us13\/_0084_ ), .B(\us13\/_0060_ ), .Y(\us13\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1136_ ( .A(\us13\/_0324_ ), .B(\us13\/_0060_ ), .Y(\us13\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1137_ ( .A(\us13\/_0335_ ), .B(\us13\/_0337_ ), .Y(\us13\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1138_ ( .A1(\us13\/_0276_ ), .A2(\us13\/_0060_ ), .B1(\us13\/_0334_ ), .C1(\us13\/_0338_ ), .Y(\us13\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1139_ ( .A(\us13\/_0318_ ), .B(\us13\/_0328_ ), .C(\us13\/_0333_ ), .D(\us13\/_0339_ ), .X(\us13\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us13/_1140_ ( .A1(\us13\/_0747_ ), .A2(\us13\/_0134_ ), .B1(\us13\/_0128_ ), .X(\us13\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us13/_1141_ ( .A_N(\us13\/_0086_ ), .B(\us13\/_0128_ ), .X(\us13\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1142_ ( .A(\us13\/_0079_ ), .B(\us13\/_0124_ ), .X(\us13\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_1143_ ( .A(\us13\/_0126_ ), .B(\us13\/_0343_ ), .Y(\us13\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us13/_1144_ ( .A(\us13\/_0341_ ), .B(\us13\/_0342_ ), .C_N(\us13\/_0344_ ), .Y(\us13\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1146_ ( .A1(\us13\/_0193_ ), .A2(\us13\/_0092_ ), .A3(\us13\/_0330_ ), .B1(\us13\/_0147_ ), .Y(\us13\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1147_ ( .A1(\us13\/_0130_ ), .A2(\us13\/_0084_ ), .A3(\us13\/_0134_ ), .B1(\us13\/_0139_ ), .Y(\us13\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1148_ ( .A1(\us13\/_0144_ ), .A2(\us13\/_0608_ ), .A3(\us13\/_0092_ ), .B1(\us13\/_0139_ ), .Y(\us13\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1149_ ( .A(\us13\/_0345_ ), .B(\us13\/_0348_ ), .C(\us13\/_0349_ ), .D(\us13\/_0350_ ), .X(\us13\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us13/_1150_ ( .A(\us13\/_0150_ ), .B(\us13\/_0194_ ), .C(\us13\/_0543_ ), .X(\us13\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us13/_1151_ ( .A(\us13\/_0277_ ), .SLEEP(\us13\/_0352_ ), .X(\us13\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us13/_1152_ ( .A1(\us13\/_0268_ ), .A2(\us13\/_0171_ ), .B1(\us13\/_0157_ ), .Y(\us13\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us13/_1153_ ( .A(\us13\/_0161_ ), .X(\us13\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1154_ ( .A1(\us13\/_0279_ ), .A2(\us13\/_0084_ ), .B1(\us13\/_0355_ ), .Y(\us13\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1155_ ( .A1(\us13\/_0020_ ), .A2(\us13\/_0193_ ), .A3(\us13\/_0091_ ), .B1(\us13\/_0355_ ), .Y(\us13\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1156_ ( .A(\us13\/_0353_ ), .B(\us13\/_0354_ ), .C(\us13\/_0356_ ), .D(\us13\/_0357_ ), .X(\us13\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1157_ ( .A(\us13\/_0111_ ), .B(\us13\/_0586_ ), .X(\us13\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1158_ ( .A(\us13\/_0360_ ), .Y(\us13\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us13/_1159_ ( .A1(\us13\/_0119_ ), .A2(\us13\/_0120_ ), .B1(\us13\/_0230_ ), .C1(\us13\/_0361_ ), .X(\us13\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1160_ ( .A1(\us13\/_0662_ ), .A2(\us13\/_0251_ ), .A3(\us13\/_0134_ ), .B1(\us13\/_0114_ ), .Y(\us13\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1162_ ( .A1(\us13\/_0036_ ), .A2(\us13\/_0251_ ), .A3(\us13\/_0134_ ), .B1(\us13\/_0099_ ), .Y(\us13\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1163_ ( .A1(\us13\/_0193_ ), .A2(\us13\/_0608_ ), .B1(\us13\/_0099_ ), .Y(\us13\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1164_ ( .A(\us13\/_0362_ ), .B(\us13\/_0363_ ), .C(\us13\/_0365_ ), .D(\us13\/_0366_ ), .X(\us13\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1165_ ( .A1(\us13\/_0575_ ), .A2(\us13\/_0092_ ), .A3(\us13\/_0330_ ), .B1(\us13\/_0089_ ), .Y(\us13\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1166_ ( .A1(\us13\/_0586_ ), .A2(\us13\/_0018_ ), .A3(\us13\/_0330_ ), .B1(\us13\/_0094_ ), .Y(\us13\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \us13/_1167_ ( .A1(\us13\/_0293_ ), .A2(\us13\/_0134_ ), .B1(\us13\/_0089_ ), .Y(\us13\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1168_ ( .A1(\us13\/_0279_ ), .A2(\us13\/_0134_ ), .B1(\us13\/_0094_ ), .Y(\us13\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1169_ ( .A(\us13\/_0368_ ), .B(\us13\/_0370_ ), .C(\us13\/_0371_ ), .D(\us13\/_0372_ ), .X(\us13\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1170_ ( .A(\us13\/_0351_ ), .B(\us13\/_0359_ ), .C(\us13\/_0367_ ), .D(\us13\/_0373_ ), .X(\us13\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1171_ ( .A1(\us13\/_0102_ ), .A2(\us13\/_0347_ ), .B1(\us13\/_0109_ ), .C1(\us13\/_0029_ ), .Y(\us13\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1172_ ( .A1(\us13\/_0102_ ), .A2(\us13\/_0347_ ), .B1(\us13\/_0532_ ), .C1(\us13\/_0029_ ), .Y(\us13\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1173_ ( .A1(\us13\/_0050_ ), .A2(\us13\/_0543_ ), .B1(\us13\/_0380_ ), .C1(\us13\/_0029_ ), .Y(\us13\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1174_ ( .A(\us13\/_0041_ ), .B(\us13\/_0375_ ), .C(\us13\/_0376_ ), .D(\us13\/_0377_ ), .X(\us13\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1175_ ( .A(\us13\/_0048_ ), .B(\us13\/_0750_ ), .X(\us13\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1176_ ( .A(\us13\/_0379_ ), .Y(\us13\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1177_ ( .A(\us13\/_0016_ ), .B(\us13\/_0608_ ), .Y(\us13\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1178_ ( .A(\us13\/_0752_ ), .B(\us13\/_0554_ ), .Y(\us13\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1179_ ( .A1(\sa13\[1\] ), .A2(\us13\/_0734_ ), .B1(\us13\/_0109_ ), .C1(\us13\/_0016_ ), .Y(\us13\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1180_ ( .A(\us13\/_0381_ ), .B(\us13\/_0382_ ), .C(\us13\/_0383_ ), .D(\us13\/_0384_ ), .X(\us13\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us13/_1181_ ( .A(\us13\/_0086_ ), .B_N(\us13\/_0736_ ), .X(\us13\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1182_ ( .A1(\us13\/_0748_ ), .A2(\us13\/_0134_ ), .B1(\us13\/_0739_ ), .Y(\us13\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1183_ ( .A1(\us13\/_0118_ ), .A2(\us13\/_0543_ ), .B1(\us13\/_0109_ ), .C1(\us13\/_0739_ ), .Y(\us13\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1184_ ( .A1(\us13\/_0102_ ), .A2(\us13\/_0301_ ), .B1(\sa13\[3\] ), .C1(\us13\/_0739_ ), .Y(\us13\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1185_ ( .A(\us13\/_0386_ ), .B(\us13\/_0387_ ), .C(\us13\/_0388_ ), .D(\us13\/_0389_ ), .X(\us13\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1186_ ( .A(\us13\/_0020_ ), .Y(\us13\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1187_ ( .A(\us13\/_0727_ ), .Y(\us13\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1188_ ( .A(\us13\/_0727_ ), .B(\us13\/_0064_ ), .Y(\us13\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1189_ ( .A1(\us13\/_0102_ ), .A2(\us13\/_0734_ ), .B1(\us13\/_0532_ ), .C1(\us13\/_0727_ ), .Y(\us13\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us13/_1190_ ( .A1(\us13\/_0392_ ), .A2(\us13\/_0393_ ), .B1(\us13\/_0394_ ), .C1(\us13\/_0395_ ), .X(\us13\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1191_ ( .A(\us13\/_0378_ ), .B(\us13\/_0385_ ), .C(\us13\/_0390_ ), .D(\us13\/_0396_ ), .X(\us13\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us13/_1192_ ( .A(\us13\/_0340_ ), .B(\us13\/_0374_ ), .C(\us13\/_0397_ ), .Y(\us13\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1193_ ( .A(\us13\/_0077_ ), .B(\us13\/_0129_ ), .X(\us13\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_1194_ ( .A(\us13\/_0398_ ), .B(\us13\/_0239_ ), .Y(\us13\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1195_ ( .A(\us13\/_0022_ ), .B(\us13\/_0111_ ), .X(\us13\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us13/_1196_ ( .A_N(\us13\/_0400_ ), .B(\us13\/_0231_ ), .Y(\us13\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us13/_1197_ ( .A(\us13\/_0399_ ), .SLEEP(\us13\/_0402_ ), .X(\us13\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_1198_ ( .A(\us13\/_0747_ ), .B(\us13\/_0251_ ), .Y(\us13\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us13/_1199_ ( .A_N(\us13\/_0404_ ), .B(\us13\/_0752_ ), .Y(\us13\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us13/_1200_ ( .A(\us13\/_0467_ ), .B(\us13\/_0194_ ), .C(\us13\/_0694_ ), .X(\us13\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us13/_1201_ ( .A_N(\us13\/_0175_ ), .B(\us13\/_0406_ ), .X(\us13\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1202_ ( .A(\us13\/_0407_ ), .Y(\us13\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1203_ ( .A1(\us13\/_0094_ ), .A2(\us13\/_0197_ ), .B1(\us13\/_0114_ ), .B2(\us13\/_0640_ ), .Y(\us13\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1204_ ( .A(\us13\/_0403_ ), .B(\us13\/_0405_ ), .C(\us13\/_0408_ ), .D(\us13\/_0409_ ), .X(\us13\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1205_ ( .A(\us13\/_0030_ ), .B(\us13\/_0150_ ), .Y(\us13\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us13/_1206_ ( .A_N(\us13\/_0169_ ), .B(\us13\/_0289_ ), .C(\us13\/_0411_ ), .X(\us13\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us13/_1207_ ( .A1(\us13\/_0467_ ), .A2(\us13\/_0151_ ), .B1(\us13\/_0140_ ), .C1(\us13\/_0129_ ), .X(\us13\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1208_ ( .A1(\us13\/_0608_ ), .A2(\us13\/_0099_ ), .B1(\us13\/_0037_ ), .C1(\us13\/_0414_ ), .Y(\us13\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1209_ ( .A(\us13\/_0738_ ), .Y(\us13\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1210_ ( .A(\us13\/_0586_ ), .B(\us13\/_0736_ ), .Y(\us13\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1211_ ( .A1(\us13\/_0194_ ), .A2(\us13\/_0038_ ), .B1(\us13\/_0118_ ), .C1(\us13\/_0153_ ), .Y(\us13\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us13/_1212_ ( .A1(\us13\/_0416_ ), .A2(\us13\/_0117_ ), .B1(\us13\/_0417_ ), .C1(\us13\/_0418_ ), .X(\us13\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1213_ ( .A(\us13\/_0077_ ), .B(\us13\/_0035_ ), .X(\us13\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1214_ ( .A(\us13\/_0662_ ), .B(\us13\/_0124_ ), .Y(\us13\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1215_ ( .A(\us13\/_0030_ ), .B(\us13\/_0137_ ), .Y(\us13\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1216_ ( .A(\us13\/_0072_ ), .B(\us13\/_0732_ ), .Y(\us13\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us13/_1217_ ( .A_N(\us13\/_0420_ ), .B(\us13\/_0421_ ), .C(\us13\/_0422_ ), .D(\us13\/_0424_ ), .X(\us13\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1218_ ( .A(\us13\/_0413_ ), .B(\us13\/_0415_ ), .C(\us13\/_0419_ ), .D(\us13\/_0425_ ), .X(\us13\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us13/_1219_ ( .A(\us13\/_0355_ ), .B(\us13\/_0102_ ), .C(\us13\/_0109_ ), .Y(\us13\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1220_ ( .A(\us13\/_0077_ ), .B(\us13\/_0018_ ), .X(\us13\/_0428_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1221_ ( .A(\us13\/_0077_ ), .B(\us13\/_0554_ ), .X(\us13\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us13/_1222_ ( .A1(\us13\/_0050_ ), .A2(\us13\/_0216_ ), .B1(\us13\/_0380_ ), .C1(\us13\/_0078_ ), .X(\us13\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us13/_1223_ ( .A(\us13\/_0428_ ), .B(\us13\/_0429_ ), .C(\us13\/_0430_ ), .Y(\us13\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us13/_1224_ ( .A_N(\us13\/_0209_ ), .B(\us13\/_0431_ ), .X(\us13\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us13/_1225_ ( .A1(\us13\/_0215_ ), .A2(\us13\/_0404_ ), .B1(\us13\/_0427_ ), .C1(\us13\/_0432_ ), .X(\us13\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1226_ ( .A(\us13\/_0043_ ), .B(\us13\/_0058_ ), .Y(\us13\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1227_ ( .A(\us13\/_0195_ ), .B(\us13\/_0233_ ), .C(\us13\/_0320_ ), .D(\us13\/_0435_ ), .X(\us13\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1228_ ( .A(\us13\/_0261_ ), .B(\us13\/_0738_ ), .Y(\us13\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1229_ ( .A1(\us13\/_0499_ ), .A2(\us13\/_0640_ ), .B1(\us13\/_0261_ ), .B2(\us13\/_0056_ ), .Y(\us13\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1230_ ( .A(\us13\/_0436_ ), .B(\us13\/_0394_ ), .C(\us13\/_0437_ ), .D(\us13\/_0438_ ), .X(\us13\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1231_ ( .A(\us13\/_0410_ ), .B(\us13\/_0426_ ), .C(\us13\/_0433_ ), .D(\us13\/_0439_ ), .X(\us13\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us13/_1232_ ( .A(\us13\/_0135_ ), .SLEEP(\us13\/_0273_ ), .X(\us13\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1233_ ( .A1(\us13\/_0279_ ), .A2(\us13\/_0134_ ), .B1(\us13\/_0099_ ), .Y(\us13\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1234_ ( .A(\us13\/_0441_ ), .B(\us13\/_0164_ ), .C(\us13\/_0270_ ), .D(\us13\/_0442_ ), .X(\us13\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1235_ ( .A(\us13\/_0051_ ), .B(\us13\/_0662_ ), .Y(\us13\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1236_ ( .A(\us13\/_0051_ ), .B(\us13\/_0271_ ), .Y(\us13\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1237_ ( .A(\us13\/_0444_ ), .B(\us13\/_0446_ ), .X(\us13\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1238_ ( .A(\us13\/_0193_ ), .B(\us13\/_0304_ ), .X(\us13\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1239_ ( .A(\us13\/_0448_ ), .Y(\us13\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1240_ ( .A(\us13\/_0162_ ), .B(\us13\/_0130_ ), .X(\us13\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1241_ ( .A(\us13\/_0450_ ), .Y(\us13\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1242_ ( .A1(\us13\/_0129_ ), .A2(\us13\/_0554_ ), .B1(\us13\/_0043_ ), .Y(\us13\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1243_ ( .A(\us13\/_0447_ ), .B(\us13\/_0449_ ), .C(\us13\/_0451_ ), .D(\us13\/_0452_ ), .X(\us13\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1244_ ( .A(\us13\/_0056_ ), .B(\us13\/_0064_ ), .Y(\us13\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us13/_1245_ ( .A_N(\us13\/_0248_ ), .B(\us13\/_0454_ ), .C(\us13\/_0254_ ), .D(\us13\/_0256_ ), .X(\us13\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1246_ ( .A1(\us13\/_0330_ ), .A2(\us13\/_0099_ ), .B1(\us13\/_0134_ ), .B2(\us13\/_0716_ ), .Y(\us13\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1247_ ( .A1(\us13\/_0748_ ), .A2(\us13\/_0738_ ), .B1(\us13\/_0092_ ), .B2(\us13\/_0752_ ), .Y(\us13\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1248_ ( .A1(\us13\/_0072_ ), .A2(\us13\/_0036_ ), .B1(\us13\/_0748_ ), .B2(\us13\/_0056_ ), .Y(\us13\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1249_ ( .A1(\us13\/_0748_ ), .A2(\us13\/_0251_ ), .B1(\us13\/_0029_ ), .Y(\us13\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1250_ ( .A(\us13\/_0457_ ), .B(\us13\/_0458_ ), .C(\us13\/_0459_ ), .D(\us13\/_0460_ ), .X(\us13\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1251_ ( .A(\us13\/_0443_ ), .B(\us13\/_0453_ ), .C(\us13\/_0455_ ), .D(\us13\/_0461_ ), .X(\us13\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1252_ ( .A(\us13\/_0705_ ), .B(\us13\/_0079_ ), .X(\us13\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1253_ ( .A(\us13\/_0586_ ), .B(\us13\/_0124_ ), .Y(\us13\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1254_ ( .A(\us13\/_0499_ ), .B(\us13\/_0747_ ), .Y(\us13\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us13/_1255_ ( .A_N(\us13\/_0463_ ), .B(\us13\/_0464_ ), .C(\us13\/_0465_ ), .X(\us13\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us13/_1256_ ( .A1(\us13\/_0271_ ), .A2(\us13\/_0072_ ), .B1(\us13\/_0142_ ), .B2(\us13\/_0027_ ), .X(\us13\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1257_ ( .A1(\us13\/_0144_ ), .A2(\us13\/_0099_ ), .B1(\us13\/_0360_ ), .C1(\us13\/_0468_ ), .Y(\us13\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us13/_1258_ ( .A1(\us13\/_0662_ ), .A2(\us13\/_0251_ ), .B1(\us13\/_0499_ ), .X(\us13\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1259_ ( .A1(\us13\/_0575_ ), .A2(\us13\/_0056_ ), .B1(\us13\/_0379_ ), .C1(\us13\/_0470_ ), .Y(\us13\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1260_ ( .A(\us13\/_0466_ ), .B(\us13\/_0469_ ), .C(\us13\/_0471_ ), .D(\us13\/_0305_ ), .X(\us13\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us13/_1261_ ( .A1(\us13\/_0029_ ), .A2(\us13\/_0683_ ), .B1(\us13\/_0324_ ), .B2(\us13\/_0056_ ), .X(\us13\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1262_ ( .A(\us13\/_0084_ ), .B(\us13\/_0099_ ), .X(\us13\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us13/_1263_ ( .A1(\us13\/_0092_ ), .A2(\us13\/_0029_ ), .B1(\us13\/_0474_ ), .X(\us13\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us13/_1264_ ( .A(\us13\/_0075_ ), .B(\us13\/_0473_ ), .C(\us13\/_0475_ ), .Y(\us13\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1265_ ( .A1(\us13\/_0279_ ), .A2(\us13\/_0255_ ), .B1(\us13\/_0084_ ), .B2(\us13\/_0060_ ), .Y(\us13\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1266_ ( .A1(\us13\/_0093_ ), .A2(\us13\/_0056_ ), .B1(\us13\/_0134_ ), .B2(\us13\/_0114_ ), .Y(\us13\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1267_ ( .A1(\us13\/_0161_ ), .A2(\us13\/_0032_ ), .B1(\us13\/_0324_ ), .B2(\us13\/_0147_ ), .Y(\us13\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1268_ ( .A1(\us13\/_0054_ ), .A2(\us13\/_0732_ ), .B1(\us13\/_0748_ ), .B2(\us13\/_0304_ ), .Y(\us13\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1269_ ( .A(\us13\/_0477_ ), .B(\us13\/_0479_ ), .C(\us13\/_0480_ ), .D(\us13\/_0481_ ), .X(\us13\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1270_ ( .A(\us13\/_0161_ ), .B(\us13\/_0064_ ), .Y(\us13\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us13/_1271_ ( .A(\us13\/_0732_ ), .B(\us13\/_0123_ ), .C(\us13\/_0467_ ), .Y(\us13\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1272_ ( .A(\us13\/_0483_ ), .B(\us13\/_0484_ ), .Y(\us13\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1273_ ( .A(\us13\/_0297_ ), .Y(\us13\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us13/_1274_ ( .A_N(\us13\/_0485_ ), .B(\us13\/_0181_ ), .C(\us13\/_0486_ ), .D(\us13\/_0386_ ), .X(\us13\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1275_ ( .A(\us13\/_0472_ ), .B(\us13\/_0476_ ), .C(\us13\/_0482_ ), .D(\us13\/_0487_ ), .X(\us13\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \us13/_1276_ ( .A(\us13\/_0440_ ), .B(\us13\/_0462_ ), .C(\us13\/_0488_ ), .Y(\us13\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1277_ ( .A(\us13\/_0403_ ), .B(\us13\/_0230_ ), .C(\us13\/_0451_ ), .D(\us13\/_0361_ ), .X(\us13\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1278_ ( .A1(\us13\/_0118_ ), .A2(\us13\/_0050_ ), .B1(\us13\/_0109_ ), .C1(\us13\/_0139_ ), .Y(\us13\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1279_ ( .A(\us13\/_0447_ ), .B(\us13\/_0437_ ), .C(\us13\/_0491_ ), .D(\us13\/_0427_ ), .X(\us13\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1280_ ( .A1(\us13\/_0084_ ), .A2(\us13\/_0255_ ), .B1(\us13\/_0608_ ), .B2(\us13\/_0029_ ), .Y(\us13\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1281_ ( .A1(\us13\/_0144_ ), .A2(\us13\/_0147_ ), .B1(\us13\/_0355_ ), .B2(\us13\/_0093_ ), .Y(\us13\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1282_ ( .A1(\us13\/_0716_ ), .A2(\us13\/_0279_ ), .B1(\us13\/_0330_ ), .B2(\us13\/_0029_ ), .Y(\us13\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1283_ ( .A1(\us13\/_0279_ ), .A2(\us13\/_0084_ ), .B1(\us13\/_0114_ ), .Y(\us13\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1284_ ( .A(\us13\/_0493_ ), .B(\us13\/_0494_ ), .C(\us13\/_0495_ ), .D(\us13\/_0496_ ), .X(\us13\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1285_ ( .A1(\us13\/_0134_ ), .A2(\us13\/_0137_ ), .B1(\us13\/_0355_ ), .B2(\us13\/_0575_ ), .Y(\us13\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1286_ ( .A1(\us13\/_0099_ ), .A2(\us13\/_0733_ ), .B1(\us13\/_0093_ ), .B2(\us13\/_0499_ ), .Y(\us13\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1287_ ( .A(\us13\/_0147_ ), .B(\us13\/_0640_ ), .Y(\us13\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1288_ ( .A1(\us13\/_0153_ ), .A2(\us13\/_0056_ ), .B1(\us13\/_0748_ ), .Y(\us13\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1289_ ( .A(\us13\/_0498_ ), .B(\us13\/_0500_ ), .C(\us13\/_0501_ ), .D(\us13\/_0502_ ), .X(\us13\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1290_ ( .A(\us13\/_0490_ ), .B(\us13\/_0492_ ), .C(\us13\/_0497_ ), .D(\us13\/_0503_ ), .X(\us13\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us13/_1291_ ( .A_N(\us13\/_0275_ ), .B(\us13\/_0716_ ), .X(\us13\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1292_ ( .A(\us13\/_0505_ ), .Y(\us13\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1293_ ( .A(\us13\/_0380_ ), .B(\us13\/_0347_ ), .X(\us13\/_0507_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1294_ ( .A1(\us13\/_0507_ ), .A2(\us13\/_0093_ ), .B1(\us13\/_0056_ ), .Y(\us13\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1295_ ( .A(\us13\/_0322_ ), .B(\us13\/_0277_ ), .C(\us13\/_0506_ ), .D(\us13\/_0508_ ), .X(\us13\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1296_ ( .A(\us13\/_0084_ ), .B(\us13\/_0716_ ), .X(\us13\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1297_ ( .A1(\us13\/_0733_ ), .A2(\us13\/_0114_ ), .B1(\us13\/_0429_ ), .C1(\us13\/_0511_ ), .Y(\us13\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_1298_ ( .A(\us13\/_0019_ ), .B(\us13\/_0024_ ), .Y(\us13\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1299_ ( .A(\us13\/_0512_ ), .B(\us13\/_0513_ ), .C(\us13\/_0742_ ), .D(\us13\/_0306_ ), .X(\us13\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1300_ ( .A1(\us13\/_0532_ ), .A2(\us13\/_0089_ ), .B1(\us13\/_0154_ ), .C1(\us13\/_0169_ ), .Y(\us13\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us13/_1301_ ( .A1(\us13\/_0749_ ), .A2(\us13\/_0026_ ), .B1(\us13\/_0069_ ), .C1(\us13\/_0032_ ), .X(\us13\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us13/_1302_ ( .A1(\us13\/_0324_ ), .A2(\us13\/_0355_ ), .B1(\us13\/_0330_ ), .B2(\us13\/_0727_ ), .X(\us13\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us13/_1303_ ( .A(\us13\/_0133_ ), .B(\us13\/_0516_ ), .C(\us13\/_0517_ ), .Y(\us13\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1304_ ( .A(\us13\/_0509_ ), .B(\us13\/_0514_ ), .C(\us13\/_0515_ ), .D(\us13\/_0518_ ), .X(\us13\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1305_ ( .A(\us13\/_0747_ ), .B(\us13\/_0072_ ), .Y(\us13\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1306_ ( .A1(\us13\/_0083_ ), .A2(\us13\/_0070_ ), .B1(\us13\/_0043_ ), .B2(\us13\/_0193_ ), .Y(\us13\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1307_ ( .A(\us13\/_0311_ ), .B(\us13\/_0520_ ), .C(\us13\/_0332_ ), .D(\us13\/_0522_ ), .X(\us13\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1308_ ( .A(\us13\/_0129_ ), .B(\us13\/_0499_ ), .X(\us13\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_1309_ ( .A(\us13\/_0235_ ), .B(\us13\/_0524_ ), .Y(\us13\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us13/_1310_ ( .A(\us13\/_0081_ ), .B(\us13\/_0085_ ), .Y(\us13\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1311_ ( .A1(\us13\/_0051_ ), .A2(\us13\/_0045_ ), .B1(\us13\/_0130_ ), .B2(\us13\/_0094_ ), .Y(\us13\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1312_ ( .A(\us13\/_0523_ ), .B(\us13\/_0525_ ), .C(\us13\/_0526_ ), .D(\us13\/_0527_ ), .X(\us13\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us13/_1313_ ( .A_N(\us13\/_0250_ ), .B(\us13\/_0521_ ), .Y(\us13\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1314_ ( .A(\us13\/_0128_ ), .B(\us13\/_0020_ ), .X(\us13\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1315_ ( .A(\us13\/_0530_ ), .Y(\us13\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1316_ ( .A(\us13\/_0099_ ), .B(\us13\/_0058_ ), .X(\us13\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1317_ ( .A(\us13\/_0533_ ), .Y(\us13\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us13/_1318_ ( .A_N(\us13\/_0529_ ), .B(\us13\/_0531_ ), .C(\us13\/_0534_ ), .D(\us13\/_0192_ ), .X(\us13\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1319_ ( .A(\us13\/_0434_ ), .B(\us13\/_0078_ ), .X(\us13\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us13/_1320_ ( .A1(\us13\/_0750_ ), .A2(\us13\/_0079_ ), .B1(\us13\/_0129_ ), .B2(\us13\/_0705_ ), .X(\us13\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1321_ ( .A1(\us13\/_0161_ ), .A2(\us13\/_0032_ ), .B1(\us13\/_0536_ ), .C1(\us13\/_0537_ ), .Y(\us13\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us13/_1322_ ( .A1(\us13\/_0747_ ), .A2(\us13\/_0162_ ), .B1(\us13\/_0079_ ), .B2(\us13\/_0043_ ), .X(\us13\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1323_ ( .A1(\us13\/_0093_ ), .A2(\us13\/_0029_ ), .B1(\us13\/_0240_ ), .C1(\us13\/_0539_ ), .Y(\us13\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1324_ ( .A(\us13\/_0434_ ), .B(\us13\/_0043_ ), .X(\us13\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us13/_1325_ ( .A1(\us13\/_0142_ ), .A2(\us13\/_0150_ ), .B1(\us13\/_0022_ ), .B2(\us13\/_0137_ ), .X(\us13\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1326_ ( .A1(\us13\/_0279_ ), .A2(\us13\/_0051_ ), .B1(\us13\/_0541_ ), .C1(\us13\/_0542_ ), .Y(\us13\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1327_ ( .A(\us13\/_0159_ ), .B(\us13\/_0036_ ), .X(\us13\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us13/_1328_ ( .A1(\us13\/_0271_ ), .A2(\us13\/_0434_ ), .B1(\us13\/_0027_ ), .X(\us13\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1329_ ( .A1(\us13\/_0091_ ), .A2(\us13\/_0128_ ), .B1(\us13\/_0545_ ), .C1(\us13\/_0546_ ), .Y(\us13\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1330_ ( .A(\us13\/_0538_ ), .B(\us13\/_0540_ ), .C(\us13\/_0544_ ), .D(\us13\/_0547_ ), .X(\us13\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1331_ ( .A(\us13\/_0099_ ), .B(\us13\/_0193_ ), .X(\us13\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us13/_1332_ ( .A(\us13\/_0549_ ), .B(\us13\/_0186_ ), .C(\us13\/_0187_ ), .Y(\us13\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1333_ ( .A(\us13\/_0062_ ), .B(\us13\/_0347_ ), .C(\us13\/_0749_ ), .D(\us13\/_0694_ ), .X(\us13\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1334_ ( .A1(\us13\/_0130_ ), .A2(\us13\/_0499_ ), .B1(\us13\/_0551_ ), .C1(\us13\/_0101_ ), .Y(\us13\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1335_ ( .A(\us13\/_0139_ ), .B(\us13\/_0640_ ), .Y(\us13\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1336_ ( .A1(\us13\/_0752_ ), .A2(\us13\/_0662_ ), .B1(\us13\/_0084_ ), .B2(\us13\/_0099_ ), .Y(\us13\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1337_ ( .A(\us13\/_0550_ ), .B(\us13\/_0552_ ), .C(\us13\/_0553_ ), .D(\us13\/_0555_ ), .X(\us13\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1338_ ( .A(\us13\/_0528_ ), .B(\us13\/_0535_ ), .C(\us13\/_0548_ ), .D(\us13\/_0556_ ), .X(\us13\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us13/_1339_ ( .A(\us13\/_0504_ ), .B(\us13\/_0519_ ), .C(\us13\/_0557_ ), .Y(\us13\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1340_ ( .A(\us13\/_0054_ ), .B(\us13\/_0507_ ), .X(\us13\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us13/_1341_ ( .A_N(\us13\/_0558_ ), .B(\us13\/_0408_ ), .C(\us13\/_0451_ ), .D(\us13\/_0452_ ), .X(\us13\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1342_ ( .A(\us13\/_0549_ ), .Y(\us13\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1343_ ( .A(\us13\/_0559_ ), .B(\us13\/_0403_ ), .C(\us13\/_0560_ ), .D(\us13\/_0371_ ), .X(\us13\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1344_ ( .A(\us13\/_0181_ ), .B(\us13\/_0178_ ), .X(\us13\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1345_ ( .A(\us13\/_0562_ ), .B(\us13\/_0552_ ), .C(\us13\/_0553_ ), .D(\us13\/_0555_ ), .X(\us13\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1346_ ( .A(\us13\/_0029_ ), .B(\us13\/_0020_ ), .Y(\us13\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1347_ ( .A(\us13\/_0051_ ), .B(\us13\/_0130_ ), .X(\us13\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1348_ ( .A(\us13\/_0566_ ), .Y(\us13\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1349_ ( .A(\us13\/_0159_ ), .B(\us13\/_0423_ ), .X(\us13\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1350_ ( .A1(\us13\/_0752_ ), .A2(\us13\/_0640_ ), .B1(\us13\/_0568_ ), .B2(\us13\/_0175_ ), .Y(\us13\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1351_ ( .A(\us13\/_0076_ ), .B(\us13\/_0565_ ), .C(\us13\/_0567_ ), .D(\us13\/_0569_ ), .X(\us13\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us13/_1352_ ( .A1(\us13\/_0036_ ), .A2(\us13\/_0142_ ), .B1(\us13\/_0161_ ), .X(\us13\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1353_ ( .A(\us13\/_0099_ ), .B(\us13\/_0662_ ), .Y(\us13\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us13/_1354_ ( .A(\us13\/_0420_ ), .B(\us13\/_0571_ ), .C_N(\us13\/_0572_ ), .Y(\us13\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1355_ ( .A(\us13\/_0051_ ), .B(\us13\/_0747_ ), .Y(\us13\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1356_ ( .A(\us13\/_0574_ ), .B(\us13\/_0319_ ), .C(\us13\/_0320_ ), .D(\us13\/_0411_ ), .X(\us13\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1357_ ( .A(\us13\/_0736_ ), .B(\us13\/_0035_ ), .Y(\us13\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1358_ ( .A(\us13\/_0736_ ), .B(\us13\/_0030_ ), .Y(\us13\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1359_ ( .A(\us13\/_0298_ ), .B(\us13\/_0208_ ), .C(\us13\/_0577_ ), .D(\us13\/_0578_ ), .X(\us13\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1360_ ( .A1(\us13\/_0020_ ), .A2(\us13\/_0137_ ), .B1(\us13\/_0261_ ), .B2(\us13\/_0128_ ), .Y(\us13\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1361_ ( .A(\us13\/_0573_ ), .B(\us13\/_0576_ ), .C(\us13\/_0579_ ), .D(\us13\/_0580_ ), .X(\us13\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1362_ ( .A(\us13\/_0561_ ), .B(\us13\/_0563_ ), .C(\us13\/_0570_ ), .D(\us13\/_0581_ ), .X(\us13\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1363_ ( .A(\us13\/_0128_ ), .B(\us13\/_0193_ ), .X(\us13\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1364_ ( .A(\us13\/_0083_ ), .B(\us13\/_0162_ ), .X(\us13\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us13/_1365_ ( .A(\us13\/_0583_ ), .B(\us13\/_0584_ ), .C_N(\us13\/_0437_ ), .Y(\us13\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us13/_1366_ ( .A(\us13\/_0150_ ), .B(\us13\/_0118_ ), .C(\us13\/_0380_ ), .Y(\us13\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us13/_1367_ ( .A_N(\us13\/_0182_ ), .B(\us13\/_0587_ ), .C(\us13\/_0323_ ), .X(\us13\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1368_ ( .A1(\us13\/_0575_ ), .A2(\us13\/_0153_ ), .B1(\us13\/_0727_ ), .B2(\us13\/_0058_ ), .Y(\us13\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1369_ ( .A1(\us13\/_0499_ ), .A2(\us13\/_0064_ ), .B1(\us13\/_0134_ ), .B2(\us13\/_0255_ ), .Y(\us13\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1370_ ( .A(\us13\/_0585_ ), .B(\us13\/_0588_ ), .C(\us13\/_0589_ ), .D(\us13\/_0590_ ), .X(\us13\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us13/_1371_ ( .A1(\us13\/_0091_ ), .A2(\us13\/_0139_ ), .B1(\us13\/_0250_ ), .Y(\us13\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1372_ ( .A1(\us13\/_0092_ ), .A2(\us13\/_0739_ ), .B1(\us13\/_0324_ ), .B2(\us13\/_0029_ ), .Y(\us13\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1373_ ( .A1(\us13\/_0144_ ), .A2(\us13\/_0153_ ), .B1(\us13\/_0683_ ), .B2(\us13\/_0056_ ), .Y(\us13\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1374_ ( .A1(\us13\/_0091_ ), .A2(\us13\/_0499_ ), .B1(\us13\/_0330_ ), .B2(\us13\/_0056_ ), .Y(\us13\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1375_ ( .A(\us13\/_0592_ ), .B(\us13\/_0593_ ), .C(\us13\/_0594_ ), .D(\us13\/_0595_ ), .X(\us13\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1376_ ( .A(\us13\/_0499_ ), .B(\us13\/_0144_ ), .Y(\us13\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1377_ ( .A(\us13\/_0312_ ), .B(\us13\/_0598_ ), .Y(\us13\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1378_ ( .A(\us13\/_0575_ ), .B(\us13\/_0147_ ), .Y(\us13\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1379_ ( .A1(\us13\/_0293_ ), .A2(\us13\/_0137_ ), .B1(\us13\/_0093_ ), .B2(\us13\/_0739_ ), .Y(\us13\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1380_ ( .A1(\us13\/_0734_ ), .A2(\us13\/_0531_ ), .B1(\us13\/_0600_ ), .C1(\us13\/_0601_ ), .Y(\us13\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1381_ ( .A1(\us13\/_0153_ ), .A2(\us13\/_0261_ ), .B1(\us13\/_0599_ ), .C1(\us13\/_0602_ ), .Y(\us13\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1382_ ( .A(\us13\/_0591_ ), .B(\us13\/_0596_ ), .C(\us13\/_0174_ ), .D(\us13\/_0603_ ), .X(\us13\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1383_ ( .A(\us13\/_0029_ ), .B(\us13\/_0144_ ), .Y(\us13\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1384_ ( .A(\us13\/_0113_ ), .B(\us13\/_0018_ ), .Y(\us13\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1385_ ( .A(\us13\/_0381_ ), .B(\us13\/_0605_ ), .C(\us13\/_0361_ ), .D(\us13\/_0606_ ), .X(\us13\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1386_ ( .A1(\us13\/_0016_ ), .A2(\us13\/_0727_ ), .B1(\us13\/_0733_ ), .Y(\us13\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1387_ ( .A1(\us13\/_0586_ ), .A2(\us13\/_0159_ ), .B1(\us13\/_0083_ ), .B2(\us13\/_0750_ ), .Y(\us13\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1388_ ( .A1(\us13\/_0142_ ), .A2(\us13\/_0162_ ), .B1(\us13\/_0079_ ), .B2(\us13\/_0054_ ), .Y(\us13\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1389_ ( .A(\us13\/_0610_ ), .B(\us13\/_0611_ ), .C(\us13\/_0105_ ), .D(\us13\/_0106_ ), .X(\us13\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1390_ ( .A1(\us13\/_0094_ ), .A2(\us13\/_0302_ ), .B1(\us13\/_0324_ ), .B2(\us13\/_0089_ ), .Y(\us13\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1391_ ( .A(\us13\/_0607_ ), .B(\us13\/_0609_ ), .C(\us13\/_0612_ ), .D(\us13\/_0613_ ), .X(\us13\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1392_ ( .A(\us13\/_0041_ ), .B(\us13\/_0170_ ), .X(\us13\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1393_ ( .A(\us13\/_0554_ ), .B(\us13\/_0027_ ), .X(\us13\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1394_ ( .A(\us13\/_0027_ ), .B(\us13\/_0261_ ), .Y(\us13\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us13/_1395_ ( .A_N(\us13\/_0616_ ), .B(\us13\/_0617_ ), .Y(\us13\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1396_ ( .A1(\us13\/_0147_ ), .A2(\us13\/_0302_ ), .B1(\us13\/_0342_ ), .C1(\us13\/_0618_ ), .Y(\us13\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1397_ ( .A(\us13\/_0614_ ), .B(\us13\/_0272_ ), .C(\us13\/_0615_ ), .D(\us13\/_0620_ ), .X(\us13\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us13/_1398_ ( .A(\us13\/_0582_ ), .B(\us13\/_0604_ ), .C(\us13\/_0621_ ), .Y(\us13\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1399_ ( .A1(\us13\/_0084_ ), .A2(\us13\/_0134_ ), .B1(\us13\/_0089_ ), .Y(\us13\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1400_ ( .A1(\us13\/_0144_ ), .A2(\us13\/_0608_ ), .A3(\us13\/_0330_ ), .B1(\us13\/_0089_ ), .Y(\us13\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1401_ ( .A1(\us13\/_0197_ ), .A2(\us13\/_0130_ ), .A3(\us13\/_0110_ ), .B1(\us13\/_0094_ ), .Y(\us13\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1402_ ( .A(\us13\/_0432_ ), .B(\us13\/_0622_ ), .C(\us13\/_0623_ ), .D(\us13\/_0624_ ), .X(\us13\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us13/_1403_ ( .A1(\us13\/_0554_ ), .A2(\us13\/_0018_ ), .A3(\us13\/_0022_ ), .B1(\us13\/_0161_ ), .X(\us13\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us13/_1404_ ( .A_N(\us13\/_0269_ ), .B(\us13\/_0170_ ), .X(\us13\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1405_ ( .A1(\us13\/_0109_ ), .A2(\us13\/_0064_ ), .A3(\us13\/_0733_ ), .B1(\us13\/_0355_ ), .Y(\us13\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us13/_1406_ ( .A_N(\us13\/_0626_ ), .B(\us13\/_0627_ ), .C(\us13\/_0353_ ), .D(\us13\/_0628_ ), .X(\us13\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1407_ ( .A1(\us13\/_0091_ ), .A2(\us13\/_0110_ ), .A3(\us13\/_0176_ ), .B1(\us13\/_0139_ ), .Y(\us13\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1408_ ( .A1(\us13\/_0020_ ), .A2(\us13\/_0261_ ), .B1(\us13\/_0147_ ), .Y(\us13\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1409_ ( .A(\us13\/_0631_ ), .B(\us13\/_0344_ ), .C(\us13\/_0421_ ), .D(\us13\/_0632_ ), .X(\us13\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us13/_1410_ ( .A1(\us13\/_0325_ ), .A2(\us13\/_0734_ ), .B1(\us13\/_0038_ ), .C1(\us13\/_0113_ ), .X(\us13\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1411_ ( .A1(\us13\/_0134_ ), .A2(\us13\/_0114_ ), .B1(\us13\/_0221_ ), .C1(\us13\/_0634_ ), .Y(\us13\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us13/_1412_ ( .A(\us13\/_0119_ ), .B_N(\us13\/_0111_ ), .Y(\us13\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1413_ ( .A1(\us13\/_0032_ ), .A2(\us13\/_0113_ ), .B1(\us13\/_0636_ ), .C1(\us13\/_0400_ ), .Y(\us13\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1414_ ( .A1(\us13\/_0732_ ), .A2(\us13\/_0293_ ), .A3(\us13\/_0251_ ), .B1(\us13\/_0099_ ), .Y(\us13\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1415_ ( .A(\us13\/_0189_ ), .B(\us13\/_0635_ ), .C(\us13\/_0637_ ), .D(\us13\/_0638_ ), .X(\us13\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1416_ ( .A(\us13\/_0625_ ), .B(\us13\/_0630_ ), .C(\us13\/_0633_ ), .D(\us13\/_0639_ ), .X(\us13\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1417_ ( .A(\us13\/_0747_ ), .B(\us13\/_0738_ ), .X(\us13\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1418_ ( .A(\us13\/_0736_ ), .B(\us13\/_0731_ ), .X(\us13\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us13/_1419_ ( .A_N(\us13\/_0643_ ), .B(\us13\/_0577_ ), .Y(\us13\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1420_ ( .A1(\us13\/_0084_ ), .A2(\us13\/_0739_ ), .B1(\us13\/_0642_ ), .C1(\us13\/_0644_ ), .Y(\us13\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1421_ ( .A1(\us13\/_0050_ ), .A2(\us13\/_0543_ ), .B1(\us13\/_0194_ ), .C1(\us13\/_0738_ ), .Y(\us13\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1422_ ( .A(\us13\/_0646_ ), .B(\us13\/_0232_ ), .C(\us13\/_0417_ ), .D(\us13\/_0578_ ), .X(\us13\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1423_ ( .A1(\us13\/_0064_ ), .A2(\us13\/_0733_ ), .B1(\us13\/_0727_ ), .Y(\us13\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1424_ ( .A1(\us13\/_0193_ ), .A2(\us13\/_0276_ ), .B1(\us13\/_0727_ ), .Y(\us13\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1425_ ( .A(\us13\/_0645_ ), .B(\us13\/_0647_ ), .C(\us13\/_0648_ ), .D(\us13\/_0649_ ), .X(\us13\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1426_ ( .A1(\us13\/_0325_ ), .A2(\us13\/_0734_ ), .B1(\us13\/_0038_ ), .C1(\us13\/_0029_ ), .Y(\us13\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1427_ ( .A1(\us13\/_0543_ ), .A2(\us13\/_0216_ ), .B1(\us13\/_0423_ ), .C1(\us13\/_0029_ ), .Y(\us13\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1428_ ( .A(\us13\/_0652_ ), .B(\us13\/_0653_ ), .X(\us13\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1429_ ( .A1(\us13\/_0733_ ), .A2(\us13\/_0748_ ), .A3(\us13\/_0324_ ), .B1(\us13\/_0016_ ), .Y(\us13\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1430_ ( .A1(\us13\/_0640_ ), .A2(\us13\/_0193_ ), .A3(\us13\/_0091_ ), .B1(\us13\/_0016_ ), .Y(\us13\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1431_ ( .A1(\us13\/_0102_ ), .A2(\us13\/_0301_ ), .B1(\sa13\[3\] ), .C1(\us13\/_0029_ ), .Y(\us13\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1432_ ( .A(\us13\/_0654_ ), .B(\us13\/_0655_ ), .C(\us13\/_0656_ ), .D(\us13\/_0657_ ), .X(\us13\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1433_ ( .A1(\us13\/_0118_ ), .A2(\us13\/_0050_ ), .B1(\us13\/_0038_ ), .C1(\us13\/_0478_ ), .Y(\us13\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us13/_1434_ ( .A_N(\us13\/_0250_ ), .B(\us13\/_0465_ ), .C(\us13\/_0659_ ), .X(\us13\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1435_ ( .A1(\us13\/_0683_ ), .A2(\us13\/_0324_ ), .B1(\us13\/_0255_ ), .Y(\us13\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1436_ ( .A1(\us13\/_0032_ ), .A2(\us13\/_0193_ ), .A3(\us13\/_0048_ ), .B1(\us13\/_0255_ ), .Y(\us13\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1437_ ( .A1(\us13\/_0144_ ), .A2(\us13\/_0586_ ), .A3(\us13\/_0048_ ), .B1(\us13\/_0499_ ), .Y(\us13\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1438_ ( .A(\us13\/_0660_ ), .B(\us13\/_0661_ ), .C(\us13\/_0663_ ), .D(\us13\/_0664_ ), .X(\us13\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1439_ ( .A1(\us13\/_0091_ ), .A2(\us13\/_0276_ ), .B1(\us13\/_0060_ ), .Y(\us13\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1440_ ( .A1(\us13\/_0144_ ), .A2(\us13\/_0608_ ), .B1(\us13\/_0056_ ), .Y(\us13\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1441_ ( .A1(\us13\/_0423_ ), .A2(\us13\/_0038_ ), .B1(\us13\/_0102_ ), .C1(\us13\/_0060_ ), .Y(\us13\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1442_ ( .A1(\sa13\[1\] ), .A2(\us13\/_0734_ ), .B1(\us13\/_0109_ ), .C1(\us13\/_0056_ ), .Y(\us13\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1443_ ( .A(\us13\/_0666_ ), .B(\us13\/_0667_ ), .C(\us13\/_0668_ ), .D(\us13\/_0669_ ), .X(\us13\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1444_ ( .A(\us13\/_0650_ ), .B(\us13\/_0658_ ), .C(\us13\/_0665_ ), .D(\us13\/_0670_ ), .X(\us13\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us13/_1445_ ( .A(\us13\/_0641_ ), .B(\us13\/_0174_ ), .C(\us13\/_0671_ ), .Y(\us13\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us13/_1446_ ( .A(\us13\/_0049_ ), .B(\us13\/_0618_ ), .C_N(\us13\/_0052_ ), .Y(\us13\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us13/_1447_ ( .A(\us13\/_0239_ ), .Y(\us13\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1448_ ( .A(\us13\/_0716_ ), .B(\us13\/_0032_ ), .Y(\us13\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1449_ ( .A1(\us13\/_0054_ ), .A2(\us13\/_0732_ ), .B1(\us13\/_0036_ ), .B2(\us13\/_0705_ ), .Y(\us13\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1450_ ( .A1(\us13\/_0304_ ), .A2(\us13\/_0732_ ), .B1(\us13\/_0048_ ), .B2(\us13\/_0750_ ), .Y(\us13\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1451_ ( .A(\us13\/_0674_ ), .B(\us13\/_0675_ ), .C(\us13\/_0676_ ), .D(\us13\/_0677_ ), .X(\us13\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us13/_1452_ ( .A_N(\us13\/_0584_ ), .B(\us13\/_0283_ ), .X(\us13\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1453_ ( .A(\us13\/_0673_ ), .B(\us13\/_0678_ ), .C(\us13\/_0679_ ), .D(\us13\/_0508_ ), .X(\us13\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1454_ ( .A1(\us13\/_0016_ ), .A2(\us13\/_0733_ ), .B1(\us13\/_0355_ ), .B2(\us13\/_0092_ ), .Y(\us13\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1455_ ( .A(\us13\/_0681_ ), .B(\us13\/_0034_ ), .X(\us13\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us13/_1456_ ( .A1(\us13\/_0330_ ), .A2(\us13\/_0139_ ), .B1(\us13\/_0324_ ), .B2(\us13\/_0089_ ), .X(\us13\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1457_ ( .A1(\us13\/_0146_ ), .A2(\us13\/_0147_ ), .B1(\us13\/_0133_ ), .C1(\us13\/_0684_ ), .Y(\us13\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1458_ ( .A(\us13\/_0113_ ), .B(\us13\/_0251_ ), .Y(\us13\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us13/_1459_ ( .A_N(\us13\/_0463_ ), .B(\us13\/_0686_ ), .C(\us13\/_0383_ ), .D(\us13\/_0464_ ), .X(\us13\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1460_ ( .A1(\us13\/_0051_ ), .A2(\us13\/_0293_ ), .B1(\us13\/_0084_ ), .B2(\us13\/_0716_ ), .Y(\us13\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1461_ ( .A1(\us13\/_0018_ ), .A2(\us13\/_0072_ ), .B1(\us13\/_0134_ ), .B2(\us13\/_0078_ ), .Y(\us13\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1462_ ( .A(\us13\/_0687_ ), .B(\us13\/_0236_ ), .C(\us13\/_0688_ ), .D(\us13\/_0689_ ), .X(\us13\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1463_ ( .A(\us13\/_0680_ ), .B(\us13\/_0682_ ), .C(\us13\/_0685_ ), .D(\us13\/_0690_ ), .X(\us13\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us13/_1464_ ( .A1(\us13\/_0532_ ), .A2(\us13\/_0380_ ), .B1(\us13\/_0102_ ), .C1(\us13\/_0355_ ), .X(\us13\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us13/_1465_ ( .A(\us13\/_0692_ ), .B(\us13\/_0338_ ), .C(\us13\/_0644_ ), .Y(\us13\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1466_ ( .A(\us13\/_0016_ ), .B(\us13\/_0020_ ), .Y(\us13\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1467_ ( .A1(\us13\/_0032_ ), .A2(\us13\/_0137_ ), .B1(\us13\/_0279_ ), .B2(\us13\/_0094_ ), .Y(\us13\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1468_ ( .A1(\us13\/_0575_ ), .A2(\us13\/_0153_ ), .B1(\us13\/_0161_ ), .B2(\us13\/_0293_ ), .Y(\us13\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1469_ ( .A(\us13\/_0259_ ), .B(\us13\/_0695_ ), .C(\us13\/_0696_ ), .D(\us13\/_0697_ ), .X(\us13\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us13/_1470_ ( .A1(\us13\/_0255_ ), .A2(\us13\/_0640_ ), .B1(\us13\/_0016_ ), .B2(\us13\/_0193_ ), .X(\us13\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1471_ ( .A1(\us13\/_0060_ ), .A2(\us13\/_0176_ ), .B1(\us13\/_0699_ ), .C1(\us13\/_0177_ ), .Y(\us13\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1472_ ( .A1(\us13\/_0091_ ), .A2(\us13\/_0499_ ), .B1(\us13\/_0092_ ), .B2(\us13\/_0716_ ), .Y(\us13\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us13/_1473_ ( .A1(\us13\/_0716_ ), .A2(\us13\/_0683_ ), .B1(\us13\/_0093_ ), .B2(\us13\/_0114_ ), .Y(\us13\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us13/_1474_ ( .A1(\us13\/_0683_ ), .A2(\us13\/_0084_ ), .B1(\us13\/_0094_ ), .Y(\us13\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us13/_1475_ ( .A1(\us13\/_0543_ ), .A2(\us13\/_0216_ ), .B1(\us13\/_0038_ ), .C1(\us13\/_0056_ ), .Y(\us13\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1476_ ( .A(\us13\/_0701_ ), .B(\us13\/_0702_ ), .C(\us13\/_0703_ ), .D(\us13\/_0704_ ), .X(\us13\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1477_ ( .A(\us13\/_0693_ ), .B(\us13\/_0698_ ), .C(\us13\/_0700_ ), .D(\us13\/_0706_ ), .X(\us13\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us13/_1478_ ( .A1(\us13\/_0113_ ), .A2(\us13\/_0640_ ), .B1(\us13\/_0099_ ), .B2(\us13\/_0058_ ), .X(\us13\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us13/_1479_ ( .A(\us13\/_0407_ ), .B(\us13\/_0708_ ), .C(\us13\/_0529_ ), .Y(\us13\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1480_ ( .A(\us13\/_0568_ ), .B(\us13\/_0175_ ), .Y(\us13\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us13/_1481_ ( .A1(\us13\/_0029_ ), .A2(\us13\/_0114_ ), .A3(\us13\/_0051_ ), .B1(\us13\/_0130_ ), .Y(\us13\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1482_ ( .A(\us13\/_0709_ ), .B(\us13\/_0550_ ), .C(\us13\/_0710_ ), .D(\us13\/_0711_ ), .X(\us13\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us13/_1483_ ( .A1(\us13\/_0114_ ), .A2(\us13\/_0064_ ), .B1(\us13\/_0261_ ), .B2(\us13\/_0089_ ), .X(\us13\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1484_ ( .A1(\us13\/_0355_ ), .A2(\us13\/_0261_ ), .B1(\us13\/_0198_ ), .C1(\us13\/_0713_ ), .Y(\us13\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1485_ ( .A(\us13\/_0586_ ), .B(\us13\/_0478_ ), .Y(\us13\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us13/_1486_ ( .A_N(\us13\/_0541_ ), .B(\us13\/_0267_ ), .C(\us13\/_0715_ ), .D(\us13\/_0320_ ), .X(\us13\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1487_ ( .A(\us13\/_0586_ ), .B(\us13\/_0070_ ), .Y(\us13\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us13/_1488_ ( .A_N(\us13\/_0211_ ), .B(\us13\/_0155_ ), .C(\us13\/_0202_ ), .D(\us13\/_0718_ ), .X(\us13\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us13/_1489_ ( .A(\us13\/_0150_ ), .B(\us13\/_0216_ ), .C(\us13\/_0380_ ), .Y(\us13\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us13/_1490_ ( .A(\us13\/_0411_ ), .B(\us13\/_0720_ ), .X(\us13\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us13/_1491_ ( .A1(\us13\/_0018_ ), .A2(\us13\/_0022_ ), .B1(\us13\/_0078_ ), .X(\us13\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us13/_1492_ ( .A1(\us13\/_0134_ ), .A2(\us13\/_0738_ ), .B1(\us13\/_0101_ ), .C1(\us13\/_0722_ ), .Y(\us13\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1493_ ( .A(\us13\/_0717_ ), .B(\us13\/_0719_ ), .C(\us13\/_0721_ ), .D(\us13\/_0723_ ), .X(\us13\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us13/_1494_ ( .A(\us13\/_0739_ ), .B(\us13\/_0193_ ), .Y(\us13\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1495_ ( .A(\us13\/_0344_ ), .B(\us13\/_0184_ ), .C(\us13\/_0449_ ), .D(\us13\/_0725_ ), .X(\us13\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us13/_1496_ ( .A(\us13\/_0712_ ), .B(\us13\/_0714_ ), .C(\us13\/_0724_ ), .D(\us13\/_0726_ ), .X(\us13\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \us13/_1497_ ( .A(\us13\/_0691_ ), .B(\us13\/_0707_ ), .C(\us13\/_0728_ ), .Y(\us13\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \us20/_0753_ ( .A(\sa20\[2\] ), .B_N(\sa20\[3\] ), .Y(\us20\/_0096_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0754_ ( .A(\sa20\[1\] ), .X(\us20\/_0107_ ) );
sky130_fd_sc_hd__and2_1 \us20/_0755_ ( .A(\us20\/_0107_ ), .B(\sa20\[0\] ), .X(\us20\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us20/_0756_ ( .A(\us20\/_0096_ ), .B(\us20\/_0118_ ), .X(\us20\/_0129_ ) );
sky130_fd_sc_hd__and2_1 \us20/_0757_ ( .A(\sa20\[7\] ), .B(\sa20\[6\] ), .X(\us20\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_0758_ ( .A(\sa20\[4\] ), .B(\sa20\[5\] ), .Y(\us20\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0759_ ( .A(\us20\/_0140_ ), .B(\us20\/_0151_ ), .X(\us20\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0761_ ( .A(\us20\/_0129_ ), .B(\us20\/_0162_ ), .X(\us20\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0762_ ( .A(\us20\/_0096_ ), .X(\us20\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \us20/_0763_ ( .A(\us20\/_0107_ ), .B_N(\sa20\[0\] ), .Y(\us20\/_0205_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0764_ ( .A(\us20\/_0205_ ), .X(\us20\/_0216_ ) );
sky130_fd_sc_hd__and3_1 \us20/_0765_ ( .A(\us20\/_0162_ ), .B(\us20\/_0194_ ), .C(\us20\/_0216_ ), .X(\us20\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us20/_0766_ ( .A(\us20\/_0183_ ), .SLEEP(\us20\/_0227_ ), .X(\us20\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \us20/_0767_ ( .A(\sa20\[0\] ), .B_N(\sa20\[1\] ), .Y(\us20\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_0768_ ( .A(\sa20\[2\] ), .B(\sa20\[3\] ), .Y(\us20\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0769_ ( .A(\us20\/_0249_ ), .B(\us20\/_0260_ ), .X(\us20\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0771_ ( .A(\us20\/_0271_ ), .X(\us20\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0772_ ( .A(\us20\/_0162_ ), .X(\us20\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_0773_ ( .A(\us20\/_0293_ ), .B(\us20\/_0304_ ), .Y(\us20\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us20/_0774_ ( .A(\us20\/_0107_ ), .Y(\us20\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us20/_0776_ ( .A(\sa20\[0\] ), .Y(\us20\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0777_ ( .A(\sa20\[2\] ), .B(\sa20\[3\] ), .X(\us20\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0779_ ( .A(\us20\/_0358_ ), .X(\us20\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_0780_ ( .A1(\us20\/_0325_ ), .A2(\us20\/_0347_ ), .B1(\us20\/_0380_ ), .C1(\us20\/_0304_ ), .Y(\us20\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us20/_0781_ ( .A_N(\us20\/_0238_ ), .B(\us20\/_0314_ ), .C(\us20\/_0391_ ), .X(\us20\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us20/_0782_ ( .A(\sa20\[3\] ), .B_N(\sa20\[2\] ), .Y(\us20\/_0412_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0783_ ( .A(\us20\/_0412_ ), .X(\us20\/_0423_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0784_ ( .A(\us20\/_0423_ ), .B(\us20\/_0205_ ), .X(\us20\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \us20/_0787_ ( .A(\sa20\[5\] ), .B_N(\sa20\[4\] ), .Y(\us20\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0788_ ( .A(\us20\/_0467_ ), .B(\us20\/_0140_ ), .X(\us20\/_0478_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_0791_ ( .A(\us20\/_0134_ ), .B(\us20\/_0218_ ), .Y(\us20\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_0792_ ( .A(\us20\/_0478_ ), .B(\us20\/_0271_ ), .Y(\us20\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0793_ ( .A(\us20\/_0194_ ), .X(\us20\/_0532_ ) );
sky130_fd_sc_hd__buf_2 \us20/_0794_ ( .A(\us20\/_0249_ ), .X(\us20\/_0543_ ) );
sky130_fd_sc_hd__and2_1 \us20/_0795_ ( .A(\us20\/_0543_ ), .B(\us20\/_0358_ ), .X(\us20\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0797_ ( .A(\us20\/_0554_ ), .X(\us20\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us20/_0798_ ( .A(\us20\/_0216_ ), .B(\us20\/_0358_ ), .X(\us20\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0800_ ( .A(\us20\/_0586_ ), .X(\us20\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_0801_ ( .A1(\us20\/_0532_ ), .A2(\us20\/_0575_ ), .A3(\us20\/_0608_ ), .B1(\us20\/_0218_ ), .Y(\us20\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us20/_0802_ ( .A(\us20\/_0401_ ), .B(\us20\/_0510_ ), .C(\us20\/_0521_ ), .D(\us20\/_0619_ ), .X(\us20\/_0629_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0803_ ( .A(\us20\/_0358_ ), .B(\us20\/_0107_ ), .X(\us20\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0805_ ( .A(\us20\/_0205_ ), .B(\us20\/_0260_ ), .X(\us20\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0806_ ( .A(\us20\/_0662_ ), .X(\us20\/_0672_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0807_ ( .A(\us20\/_0672_ ), .X(\us20\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us20/_0808_ ( .A(\sa20\[6\] ), .B_N(\sa20\[7\] ), .Y(\us20\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \us20/_0809_ ( .A(\us20\/_0467_ ), .B(\us20\/_0694_ ), .X(\us20\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0811_ ( .A(\us20\/_0705_ ), .X(\us20\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_0812_ ( .A1(\us20\/_0640_ ), .A2(\us20\/_0293_ ), .A3(\us20\/_0683_ ), .B1(\us20\/_0727_ ), .Y(\us20\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_0813_ ( .A(\us20\/_0107_ ), .B(\sa20\[0\] ), .Y(\us20\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0814_ ( .A(\us20\/_0730_ ), .B(\us20\/_0260_ ), .X(\us20\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0815_ ( .A(\us20\/_0731_ ), .X(\us20\/_0732_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0816_ ( .A(\us20\/_0732_ ), .X(\us20\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0817_ ( .A(\sa20\[0\] ), .X(\us20\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us20/_0818_ ( .A1(\us20\/_0325_ ), .A2(\us20\/_0734_ ), .B1(\us20\/_0423_ ), .X(\us20\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0819_ ( .A(\us20\/_0694_ ), .B(\us20\/_0151_ ), .X(\us20\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0821_ ( .A(\us20\/_0736_ ), .X(\us20\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0822_ ( .A(\us20\/_0738_ ), .X(\us20\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_0823_ ( .A1(\us20\/_0733_ ), .A2(\us20\/_0735_ ), .A3(\us20\/_0293_ ), .B1(\us20\/_0739_ ), .Y(\us20\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us20/_0824_ ( .A(\us20\/_0730_ ), .B_N(\us20\/_0358_ ), .Y(\us20\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_0825_ ( .A(\us20\/_0741_ ), .B(\us20\/_0739_ ), .Y(\us20\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_0827_ ( .A1(\us20\/_0118_ ), .A2(\us20\/_0216_ ), .B1(\us20\/_0532_ ), .C1(\us20\/_0739_ ), .Y(\us20\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us20/_0828_ ( .A(\us20\/_0729_ ), .B(\us20\/_0740_ ), .C(\us20\/_0742_ ), .D(\us20\/_0744_ ), .X(\us20\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0829_ ( .A(\us20\/_0423_ ), .B(\us20\/_0730_ ), .X(\us20\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0831_ ( .A(\us20\/_0746_ ), .X(\us20\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us20/_0832_ ( .A(\sa20\[4\] ), .B_N(\sa20\[5\] ), .Y(\us20\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0833_ ( .A(\us20\/_0749_ ), .B(\us20\/_0694_ ), .X(\us20\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0835_ ( .A(\us20\/_0750_ ), .X(\us20\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0836_ ( .A(\us20\/_0752_ ), .X(\us20\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0837_ ( .A(\us20\/_0118_ ), .B(\us20\/_0358_ ), .X(\us20\/_0017_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0839_ ( .A(\us20\/_0752_ ), .B(\us20\/_0017_ ), .X(\us20\/_0019_ ) );
sky130_fd_sc_hd__and2_1 \us20/_0840_ ( .A(\us20\/_0358_ ), .B(\us20\/_0325_ ), .X(\us20\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0842_ ( .A(\us20\/_0096_ ), .B(\us20\/_0205_ ), .X(\us20\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \us20/_0844_ ( .A1(\us20\/_0020_ ), .A2(\us20\/_0022_ ), .B1(\us20\/_0752_ ), .X(\us20\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_0845_ ( .A1(\us20\/_0748_ ), .A2(\us20\/_0016_ ), .B1(\us20\/_0019_ ), .C1(\us20\/_0024_ ), .Y(\us20\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \us20/_0846_ ( .A(\sa20\[4\] ), .B(\sa20\[5\] ), .X(\us20\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0847_ ( .A(\us20\/_0694_ ), .B(\us20\/_0026_ ), .X(\us20\/_0027_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0850_ ( .A(\us20\/_0358_ ), .B(\us20\/_0730_ ), .X(\us20\/_0030_ ) );
sky130_fd_sc_hd__buf_2 \us20/_0852_ ( .A(\us20\/_0030_ ), .X(\us20\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_0853_ ( .A(\us20\/_0247_ ), .B(\us20\/_0032_ ), .Y(\us20\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_0854_ ( .A(\us20\/_0247_ ), .B(\us20\/_0735_ ), .Y(\us20\/_0034_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0855_ ( .A(\us20\/_0118_ ), .B(\us20\/_0260_ ), .X(\us20\/_0035_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0857_ ( .A(\us20\/_0027_ ), .B(\us20\/_0035_ ), .X(\us20\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0858_ ( .A(\us20\/_0260_ ), .X(\us20\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_0859_ ( .A(\us20\/_0038_ ), .B(\us20\/_0347_ ), .Y(\us20\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us20/_0860_ ( .A_N(\us20\/_0039_ ), .B(\us20\/_0027_ ), .X(\us20\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_0861_ ( .A(\us20\/_0037_ ), .B(\us20\/_0040_ ), .Y(\us20\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us20/_0862_ ( .A(\us20\/_0025_ ), .B(\us20\/_0033_ ), .C(\us20\/_0034_ ), .D(\us20\/_0041_ ), .X(\us20\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0863_ ( .A(\us20\/_0749_ ), .B(\us20\/_0140_ ), .X(\us20\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us20/_0865_ ( .A(\sa20\[0\] ), .B(\sa20\[2\] ), .C(\sa20\[3\] ), .X(\us20\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0866_ ( .A(\us20\/_0043_ ), .B(\us20\/_0045_ ), .X(\us20\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0867_ ( .A(\us20\/_0096_ ), .B(\us20\/_0543_ ), .X(\us20\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0869_ ( .A(\us20\/_0047_ ), .B(\us20\/_0043_ ), .X(\us20\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0870_ ( .A(\us20\/_0730_ ), .X(\us20\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0871_ ( .A(\us20\/_0043_ ), .X(\us20\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_0872_ ( .A1(\us20\/_0118_ ), .A2(\us20\/_0050_ ), .B1(\us20\/_0194_ ), .C1(\us20\/_0051_ ), .Y(\us20\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us20/_0873_ ( .A(\us20\/_0046_ ), .B(\us20\/_0049_ ), .C_N(\us20\/_0052_ ), .Y(\us20\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0874_ ( .A(\us20\/_0026_ ), .B(\us20\/_0140_ ), .X(\us20\/_0054_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_0877_ ( .A1(\us20\/_0532_ ), .A2(\us20\/_0575_ ), .B1(\us20\/_0292_ ), .Y(\us20\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0878_ ( .A(\us20\/_0423_ ), .B(\us20\/_0325_ ), .X(\us20\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0880_ ( .A(\us20\/_0051_ ), .X(\us20\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_0881_ ( .A1(\us20\/_0732_ ), .A2(\us20\/_0035_ ), .A3(\us20\/_0058_ ), .B1(\us20\/_0060_ ), .Y(\us20\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0882_ ( .A(\us20\/_0260_ ), .B(\us20\/_0107_ ), .X(\us20\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0884_ ( .A(\us20\/_0062_ ), .X(\us20\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_0885_ ( .A1(\us20\/_0064_ ), .A2(\us20\/_0748_ ), .A3(\us20\/_0683_ ), .B1(\us20\/_0292_ ), .Y(\us20\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us20/_0886_ ( .A(\us20\/_0053_ ), .B(\us20\/_0057_ ), .C(\us20\/_0061_ ), .D(\us20\/_0065_ ), .X(\us20\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us20/_0887_ ( .A(\us20\/_0629_ ), .B(\us20\/_0745_ ), .C(\us20\/_0042_ ), .D(\us20\/_0066_ ), .X(\us20\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us20/_0889_ ( .A(\sa20\[7\] ), .B_N(\sa20\[6\] ), .Y(\us20\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0890_ ( .A(\us20\/_0069_ ), .B(\us20\/_0151_ ), .X(\us20\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0892_ ( .A(\us20\/_0070_ ), .X(\us20\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_0893_ ( .A1(\us20\/_0129_ ), .A2(\us20\/_0586_ ), .B1(\us20\/_0072_ ), .Y(\us20\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_0894_ ( .A1(\us20\/_0380_ ), .A2(\us20\/_0347_ ), .B1(\us20\/_0194_ ), .B2(\us20\/_0216_ ), .Y(\us20\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us20/_0895_ ( .A(\us20\/_0074_ ), .B_N(\us20\/_0070_ ), .Y(\us20\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us20/_0896_ ( .A(\us20\/_0073_ ), .SLEEP(\us20\/_0075_ ), .X(\us20\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us20/_0897_ ( .A(\us20\/_0467_ ), .B(\us20\/_0069_ ), .X(\us20\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0898_ ( .A(\us20\/_0077_ ), .X(\us20\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0899_ ( .A(\us20\/_0412_ ), .B(\us20\/_0118_ ), .X(\us20\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0901_ ( .A(\us20\/_0078_ ), .B(\us20\/_0079_ ), .X(\us20\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0902_ ( .A(\us20\/_0412_ ), .B(\us20\/_0249_ ), .X(\us20\/_0082_ ) );
sky130_fd_sc_hd__buf_2 \us20/_0904_ ( .A(\us20\/_0082_ ), .X(\us20\/_0084_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0905_ ( .A(\us20\/_0084_ ), .B(\us20\/_0078_ ), .X(\us20\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us20/_0906_ ( .A1(\sa20\[0\] ), .A2(\us20\/_0325_ ), .B1(\us20\/_0260_ ), .Y(\us20\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us20/_0907_ ( .A_N(\us20\/_0086_ ), .B(\us20\/_0078_ ), .X(\us20\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us20/_0908_ ( .A(\us20\/_0081_ ), .B(\us20\/_0085_ ), .C(\us20\/_0087_ ), .Y(\us20\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0909_ ( .A(\us20\/_0072_ ), .X(\us20\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_0910_ ( .A1(\us20\/_0733_ ), .A2(\us20\/_0748_ ), .A3(\us20\/_0683_ ), .B1(\us20\/_0089_ ), .Y(\us20\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0911_ ( .A(\us20\/_0129_ ), .X(\us20\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0912_ ( .A(\us20\/_0017_ ), .X(\us20\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0913_ ( .A(\us20\/_0022_ ), .X(\us20\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0914_ ( .A(\us20\/_0078_ ), .X(\us20\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_0915_ ( .A1(\us20\/_0091_ ), .A2(\us20\/_0092_ ), .A3(\us20\/_0093_ ), .B1(\us20\/_0094_ ), .Y(\us20\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us20/_0916_ ( .A(\us20\/_0076_ ), .B(\us20\/_0088_ ), .C(\us20\/_0090_ ), .D(\us20\/_0095_ ), .X(\us20\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us20/_0917_ ( .A(\us20\/_0069_ ), .B(\us20\/_0026_ ), .X(\us20\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \us20/_0918_ ( .A(\us20\/_0098_ ), .X(\us20\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0919_ ( .A(\us20\/_0434_ ), .B(\us20\/_0099_ ), .X(\us20\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0920_ ( .A(\us20\/_0079_ ), .B(\us20\/_0098_ ), .X(\us20\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0921_ ( .A(\us20\/_0325_ ), .X(\us20\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_0922_ ( .A1(\us20\/_0102_ ), .A2(\us20\/_0734_ ), .B1(\us20\/_0038_ ), .C1(\us20\/_0099_ ), .Y(\us20\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us20/_0923_ ( .A(\us20\/_0100_ ), .B(\us20\/_0101_ ), .C_N(\us20\/_0103_ ), .Y(\us20\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_0924_ ( .A1(\us20\/_0554_ ), .A2(\us20\/_0586_ ), .B1(\us20\/_0099_ ), .Y(\us20\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_0925_ ( .A(\us20\/_0129_ ), .B(\us20\/_0099_ ), .Y(\us20\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0926_ ( .A(\us20\/_0105_ ), .B(\us20\/_0106_ ), .X(\us20\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0927_ ( .A(\us20\/_0423_ ), .X(\us20\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us20/_0928_ ( .A(\us20\/_0260_ ), .B(\sa20\[0\] ), .X(\us20\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0929_ ( .A(\us20\/_0069_ ), .B(\us20\/_0749_ ), .X(\us20\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0931_ ( .A(\us20\/_0111_ ), .X(\us20\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0932_ ( .A(\us20\/_0113_ ), .X(\us20\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_0933_ ( .A1(\us20\/_0109_ ), .A2(\us20\/_0110_ ), .B1(\us20\/_0114_ ), .Y(\us20\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us20/_0934_ ( .A(\us20\/_0022_ ), .Y(\us20\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us20/_0935_ ( .A(\us20\/_0554_ ), .Y(\us20\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us20/_0936_ ( .A1(\us20\/_0050_ ), .A2(\us20\/_0118_ ), .B1(\us20\/_0194_ ), .Y(\us20\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us20/_0937_ ( .A(\us20\/_0113_ ), .Y(\us20\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us20/_0938_ ( .A1(\us20\/_0116_ ), .A2(\us20\/_0117_ ), .A3(\us20\/_0119_ ), .B1(\us20\/_0120_ ), .X(\us20\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us20/_0939_ ( .A(\us20\/_0104_ ), .B(\us20\/_0108_ ), .C(\us20\/_0115_ ), .D(\us20\/_0121_ ), .X(\us20\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_0940_ ( .A(\sa20\[7\] ), .B(\sa20\[6\] ), .Y(\us20\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0941_ ( .A(\us20\/_0749_ ), .B(\us20\/_0123_ ), .X(\us20\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0943_ ( .A(\us20\/_0082_ ), .B(\us20\/_0124_ ), .X(\us20\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_0944_ ( .A(\us20\/_0271_ ), .B(\us20\/_0124_ ), .Y(\us20\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0945_ ( .A(\us20\/_0124_ ), .X(\us20\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0946_ ( .A(\us20\/_0260_ ), .B(\us20\/_0325_ ), .X(\us20\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_0948_ ( .A(\us20\/_0128_ ), .B(\us20\/_0130_ ), .Y(\us20\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_0949_ ( .A(\us20\/_0127_ ), .B(\us20\/_0132_ ), .Y(\us20\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us20/_0950_ ( .A(\us20\/_0434_ ), .X(\us20\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_0951_ ( .A(\us20\/_0134_ ), .B(\us20\/_0128_ ), .Y(\us20\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us20/_0952_ ( .A(\us20\/_0126_ ), .B(\us20\/_0133_ ), .C_N(\us20\/_0135_ ), .Y(\us20\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us20/_0953_ ( .A(\us20\/_0026_ ), .B(\us20\/_0123_ ), .X(\us20\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0955_ ( .A(\us20\/_0137_ ), .X(\us20\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_0956_ ( .A1(\us20\/_0110_ ), .A2(\us20\/_0293_ ), .A3(\us20\/_0084_ ), .B1(\us20\/_0139_ ), .Y(\us20\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0957_ ( .A(\us20\/_0096_ ), .B(\us20\/_0730_ ), .X(\us20\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0959_ ( .A(\us20\/_0142_ ), .X(\us20\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_0960_ ( .A1(\us20\/_0020_ ), .A2(\us20\/_0144_ ), .A3(\us20\/_0017_ ), .B1(\us20\/_0139_ ), .Y(\us20\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \us20/_0961_ ( .A(\sa20\[2\] ), .B(\us20\/_0050_ ), .C_N(\sa20\[3\] ), .Y(\us20\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0962_ ( .A(\us20\/_0128_ ), .X(\us20\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_0963_ ( .A1(\us20\/_0146_ ), .A2(\us20\/_0032_ ), .A3(\us20\/_0640_ ), .B1(\us20\/_0147_ ), .Y(\us20\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us20/_0964_ ( .A(\us20\/_0136_ ), .B(\us20\/_0141_ ), .C(\us20\/_0145_ ), .D(\us20\/_0148_ ), .X(\us20\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0965_ ( .A(\us20\/_0123_ ), .B(\us20\/_0151_ ), .X(\us20\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0967_ ( .A(\us20\/_0150_ ), .X(\us20\/_0153_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0968_ ( .A(\us20\/_0150_ ), .B(\us20\/_0062_ ), .X(\us20\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_0969_ ( .A(\us20\/_0079_ ), .B(\us20\/_0150_ ), .Y(\us20\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us20/_0970_ ( .A(\us20\/_0150_ ), .B(\us20\/_0423_ ), .C(\us20\/_0543_ ), .Y(\us20\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_0971_ ( .A(\us20\/_0155_ ), .B(\us20\/_0156_ ), .Y(\us20\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_0972_ ( .A1(\us20\/_0153_ ), .A2(\us20\/_0134_ ), .B1(\us20\/_0154_ ), .C1(\us20\/_0157_ ), .Y(\us20\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0973_ ( .A(\us20\/_0467_ ), .B(\us20\/_0123_ ), .X(\us20\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_0975_ ( .A(\us20\/_0159_ ), .X(\us20\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us20/_0976_ ( .A_N(\us20\/_0119_ ), .B(\us20\/_0161_ ), .X(\us20\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us20/_0977_ ( .A(\us20\/_0163_ ), .Y(\us20\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_0978_ ( .A1(\us20\/_0146_ ), .A2(\us20\/_0575_ ), .A3(\us20\/_0608_ ), .B1(\us20\/_0153_ ), .Y(\us20\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_0979_ ( .A1(\us20\/_0062_ ), .A2(\us20\/_0084_ ), .A3(\us20\/_0134_ ), .B1(\us20\/_0161_ ), .Y(\us20\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us20/_0980_ ( .A(\us20\/_0158_ ), .B(\us20\/_0164_ ), .C(\us20\/_0165_ ), .D(\us20\/_0166_ ), .X(\us20\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us20/_0981_ ( .A(\us20\/_0097_ ), .B(\us20\/_0122_ ), .C(\us20\/_0149_ ), .D(\us20\/_0167_ ), .X(\us20\/_0168_ ) );
sky130_fd_sc_hd__and2_1 \us20/_0982_ ( .A(\us20\/_0672_ ), .B(\us20\/_0150_ ), .X(\us20\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_0983_ ( .A(\us20\/_0154_ ), .B(\us20\/_0169_ ), .Y(\us20\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us20/_0984_ ( .A(\us20\/_0123_ ), .B(\us20\/_0151_ ), .C(\us20\/_0038_ ), .X(\us20\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0985_ ( .A(\us20\/_0170_ ), .B(\us20\/_0171_ ), .X(\us20\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \us20/_0986_ ( .A(\us20\/_0172_ ), .Y(\us20\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \us20/_0987_ ( .A(\us20\/_0067_ ), .B(\us20\/_0168_ ), .C(\us20\/_0174_ ), .Y(\us20\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us20/_0988_ ( .A(\us20\/_0107_ ), .B(\sa20\[0\] ), .Y(\us20\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us20/_0989_ ( .A(\us20\/_0175_ ), .B(\us20\/_0358_ ), .X(\us20\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0990_ ( .A(\us20\/_0176_ ), .B(\us20\/_0478_ ), .X(\us20\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_0991_ ( .A(\us20\/_0084_ ), .B(\us20\/_0113_ ), .Y(\us20\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0992_ ( .A(\us20\/_0111_ ), .B(\us20\/_0062_ ), .X(\us20\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0993_ ( .A(\us20\/_0111_ ), .B(\us20\/_0672_ ), .X(\us20\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_0994_ ( .A(\us20\/_0179_ ), .B(\us20\/_0180_ ), .Y(\us20\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0995_ ( .A(\us20\/_0054_ ), .B(\us20\/_0058_ ), .X(\us20\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us20/_0996_ ( .A(\us20\/_0182_ ), .Y(\us20\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us20/_0997_ ( .A_N(\us20\/_0177_ ), .B(\us20\/_0178_ ), .C(\us20\/_0181_ ), .D(\us20\/_0184_ ), .X(\us20\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0998_ ( .A(\us20\/_0098_ ), .B(\us20\/_0741_ ), .X(\us20\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us20/_0999_ ( .A(\us20\/_0047_ ), .B(\us20\/_0098_ ), .X(\us20\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us20/_1000_ ( .A(\us20\/_0186_ ), .B(\us20\/_0187_ ), .X(\us20\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1001_ ( .A(\us20\/_0188_ ), .Y(\us20\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1002_ ( .A(\us20\/_0738_ ), .B(\us20\/_0735_ ), .X(\us20\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1003_ ( .A(\us20\/_0271_ ), .B(\us20\/_0736_ ), .X(\us20\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_1004_ ( .A(\us20\/_0190_ ), .B(\us20\/_0191_ ), .Y(\us20\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us20/_1005_ ( .A(\us20\/_0096_ ), .B(\us20\/_0325_ ), .X(\us20\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1006_ ( .A1(\us20\/_0193_ ), .A2(\us20\/_0176_ ), .B1(\us20\/_0043_ ), .Y(\us20\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1007_ ( .A(\us20\/_0185_ ), .B(\us20\/_0189_ ), .C(\us20\/_0192_ ), .D(\us20\/_0195_ ), .X(\us20\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us20/_1008_ ( .A_N(\sa20\[3\] ), .B(\us20\/_0734_ ), .C(\sa20\[2\] ), .X(\us20\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1009_ ( .A(\us20\/_0137_ ), .B(\us20\/_0197_ ), .X(\us20\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_1010_ ( .A(\us20\/_0198_ ), .B(\us20\/_0040_ ), .Y(\us20\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1011_ ( .A(\us20\/_0293_ ), .B(\us20\/_0137_ ), .X(\us20\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1012_ ( .A(\us20\/_0200_ ), .Y(\us20\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1013_ ( .A(\us20\/_0137_ ), .B(\us20\/_0110_ ), .Y(\us20\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1014_ ( .A(\us20\/_0139_ ), .B(\us20\/_0020_ ), .Y(\us20\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1015_ ( .A(\us20\/_0199_ ), .B(\us20\/_0201_ ), .C(\us20\/_0202_ ), .D(\us20\/_0203_ ), .X(\us20\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us20/_1016_ ( .A1(\us20\/_0532_ ), .A2(\us20\/_0109_ ), .B1(\us20\/_0102_ ), .C1(\us20\/_0727_ ), .X(\us20\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1017_ ( .A(\us20\/_0022_ ), .B(\us20\/_0078_ ), .Y(\us20\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1018_ ( .A(\us20\/_0078_ ), .B(\us20\/_0142_ ), .Y(\us20\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1019_ ( .A(\us20\/_0207_ ), .B(\us20\/_0208_ ), .Y(\us20\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1020_ ( .A1(\us20\/_0094_ ), .A2(\us20\/_0176_ ), .B1(\us20\/_0206_ ), .C1(\us20\/_0209_ ), .Y(\us20\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1021_ ( .A(\us20\/_0662_ ), .B(\us20\/_0070_ ), .X(\us20\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us20/_1022_ ( .A(\us20\/_0732_ ), .B(\us20\/_0123_ ), .C(\us20\/_0749_ ), .Y(\us20\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us20/_1023_ ( .A(\us20\/_0732_ ), .B(\us20\/_0467_ ), .C(\us20\/_0069_ ), .Y(\us20\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us20/_1024_ ( .A_N(\us20\/_0211_ ), .B(\us20\/_0127_ ), .C(\us20\/_0212_ ), .D(\us20\/_0213_ ), .X(\us20\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1025_ ( .A(\us20\/_0137_ ), .Y(\us20\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1026_ ( .A(\us20\/_0128_ ), .B(\us20\/_0035_ ), .Y(\us20\/_0217_ ) );
sky130_fd_sc_hd__buf_2 \us20/_1027_ ( .A(\us20\/_0478_ ), .X(\us20\/_0218_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1028_ ( .A1(\us20\/_0159_ ), .A2(\us20\/_0746_ ), .B1(\us20\/_0434_ ), .B2(\us20\/_0218_ ), .Y(\us20\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us20/_1029_ ( .A1(\us20\/_0116_ ), .A2(\us20\/_0215_ ), .B1(\us20\/_0217_ ), .C1(\us20\/_0219_ ), .X(\us20\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1030_ ( .A(\us20\/_0113_ ), .B(\us20\/_0746_ ), .X(\us20\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us20/_1031_ ( .A1(\us20\/_0098_ ), .A2(\us20\/_0746_ ), .B1(\us20\/_0434_ ), .B2(\us20\/_0750_ ), .X(\us20\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1032_ ( .A1(\us20\/_0047_ ), .A2(\us20\/_0113_ ), .B1(\us20\/_0221_ ), .C1(\us20\/_0222_ ), .Y(\us20\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us20/_1033_ ( .A1(\us20\/_0129_ ), .A2(\us20\/_0162_ ), .B1(\us20\/_0271_ ), .B2(\us20\/_0705_ ), .X(\us20\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1034_ ( .A1(\us20\/_0093_ ), .A2(\us20\/_0738_ ), .B1(\us20\/_0081_ ), .C1(\us20\/_0224_ ), .Y(\us20\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1035_ ( .A(\us20\/_0214_ ), .B(\us20\/_0220_ ), .C(\us20\/_0223_ ), .D(\us20\/_0225_ ), .X(\us20\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1036_ ( .A(\us20\/_0196_ ), .B(\us20\/_0204_ ), .C(\us20\/_0210_ ), .D(\us20\/_0226_ ), .X(\us20\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1037_ ( .A(\us20\/_0111_ ), .B(\us20\/_0554_ ), .X(\us20\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1038_ ( .A(\us20\/_0229_ ), .Y(\us20\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1039_ ( .A(\us20\/_0111_ ), .B(\us20\/_0129_ ), .Y(\us20\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1040_ ( .A(\us20\/_0017_ ), .B(\us20\/_0738_ ), .Y(\us20\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1041_ ( .A(\us20\/_0030_ ), .B(\us20\/_0304_ ), .Y(\us20\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1042_ ( .A(\us20\/_0230_ ), .B(\us20\/_0231_ ), .C(\us20\/_0232_ ), .D(\us20\/_0233_ ), .X(\us20\/_0234_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1043_ ( .A(\us20\/_0047_ ), .B(\us20\/_0478_ ), .X(\us20\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1044_ ( .A1(\us20\/_0129_ ), .A2(\us20\/_0554_ ), .B1(\us20\/_0137_ ), .Y(\us20\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us20/_1045_ ( .A(\us20\/_0235_ ), .B(\us20\/_0049_ ), .C_N(\us20\/_0236_ ), .Y(\us20\/_0237_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1046_ ( .A(\us20\/_0047_ ), .B(\us20\/_0077_ ), .X(\us20\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1047_ ( .A(\us20\/_0070_ ), .B(\us20\/_0035_ ), .X(\us20\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us20/_1048_ ( .A1(\us20\/_0047_ ), .A2(\us20\/_0736_ ), .B1(\us20\/_0022_ ), .B2(\us20\/_0099_ ), .X(\us20\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us20/_1049_ ( .A(\us20\/_0239_ ), .B(\us20\/_0240_ ), .C(\us20\/_0241_ ), .Y(\us20\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1050_ ( .A(\us20\/_0554_ ), .B(\us20\/_0072_ ), .X(\us20\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us20/_1051_ ( .A1(\us20\/_0142_ ), .A2(\us20\/_0137_ ), .B1(\us20\/_0159_ ), .B2(\us20\/_0082_ ), .X(\us20\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1052_ ( .A1(\us20\/_0608_ ), .A2(\us20\/_0072_ ), .B1(\us20\/_0243_ ), .C1(\us20\/_0244_ ), .Y(\us20\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1053_ ( .A(\us20\/_0234_ ), .B(\us20\/_0237_ ), .C(\us20\/_0242_ ), .D(\us20\/_0245_ ), .X(\us20\/_0246_ ) );
sky130_fd_sc_hd__buf_2 \us20/_1054_ ( .A(\us20\/_0027_ ), .X(\us20\/_0247_ ) );
sky130_fd_sc_hd__o21a_1 \us20/_1055_ ( .A1(\us20\/_0554_ ), .A2(\us20\/_0586_ ), .B1(\us20\/_0247_ ), .X(\us20\/_0248_ ) );
sky130_fd_sc_hd__and2_1 \us20/_1056_ ( .A(\us20\/_0082_ ), .B(\us20\/_0478_ ), .X(\us20\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_1057_ ( .A(\us20\/_0079_ ), .X(\us20\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1058_ ( .A(\us20\/_0251_ ), .B(\us20\/_0478_ ), .X(\us20\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_1059_ ( .A(\us20\/_0250_ ), .B(\us20\/_0252_ ), .Y(\us20\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1060_ ( .A(\us20\/_0016_ ), .B(\us20\/_0064_ ), .Y(\us20\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_1061_ ( .A(\us20\/_0304_ ), .X(\us20\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1062_ ( .A(\us20\/_0255_ ), .B(\us20\/_0640_ ), .Y(\us20\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us20/_1063_ ( .A_N(\us20\/_0248_ ), .B(\us20\/_0253_ ), .C(\us20\/_0254_ ), .D(\us20\/_0256_ ), .X(\us20\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1064_ ( .A(\us20\/_0099_ ), .B(\us20\/_0110_ ), .X(\us20\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us20/_1065_ ( .A1(\us20\/_0161_ ), .A2(\us20\/_0130_ ), .B1(\us20\/_0258_ ), .Y(\us20\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1066_ ( .A(\us20\/_0194_ ), .B(\us20\/_0107_ ), .X(\us20\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1068_ ( .A(\us20\/_0261_ ), .B(\us20\/_0153_ ), .Y(\us20\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us20/_1069_ ( .A_N(\us20\/_0154_ ), .B(\us20\/_0259_ ), .C(\us20\/_0263_ ), .X(\us20\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1070_ ( .A(\us20\/_0246_ ), .B(\us20\/_0174_ ), .C(\us20\/_0257_ ), .D(\us20\/_0264_ ), .X(\us20\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us20/_1071_ ( .A1(\us20\/_0261_ ), .A2(\us20\/_0554_ ), .B1(\us20\/_0159_ ), .X(\us20\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1072_ ( .A(\us20\/_0746_ ), .B(\us20\/_0150_ ), .Y(\us20\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1073_ ( .A(\us20\/_0175_ ), .Y(\us20\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us20/_1074_ ( .A(\us20\/_0423_ ), .B(\us20\/_0123_ ), .C(\us20\/_0151_ ), .X(\us20\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1075_ ( .A(\us20\/_0268_ ), .B(\us20\/_0269_ ), .Y(\us20\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us20/_1076_ ( .A_N(\us20\/_0266_ ), .B(\us20\/_0267_ ), .C(\us20\/_0270_ ), .X(\us20\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1077_ ( .A(\us20\/_0554_ ), .B(\us20\/_0150_ ), .X(\us20\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1078_ ( .A(\us20\/_0273_ ), .Y(\us20\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1079_ ( .A1(\us20\/_0734_ ), .A2(\us20\/_0325_ ), .B1(\us20\/_0380_ ), .Y(\us20\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1080_ ( .A(\us20\/_0275_ ), .Y(\us20\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1081_ ( .A(\us20\/_0276_ ), .B(\us20\/_0153_ ), .Y(\us20\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us20/_1082_ ( .A(\us20\/_0272_ ), .B(\us20\/_0274_ ), .C(\us20\/_0277_ ), .X(\us20\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_1083_ ( .A(\us20\/_0035_ ), .X(\us20\/_0279_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1085_ ( .A1(\us20\/_0218_ ), .A2(\us20\/_0279_ ), .B1(\us20\/_0084_ ), .B2(\us20\/_0060_ ), .Y(\us20\/_0281_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1086_ ( .A1(\us20\/_0251_ ), .A2(\us20\/_0434_ ), .B1(\us20\/_0304_ ), .Y(\us20\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1087_ ( .A(\us20\/_0091_ ), .B(\us20\/_0292_ ), .Y(\us20\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1088_ ( .A1(\us20\/_0118_ ), .A2(\us20\/_0050_ ), .B1(\us20\/_0038_ ), .C1(\us20\/_0255_ ), .Y(\us20\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1089_ ( .A(\us20\/_0281_ ), .B(\us20\/_0283_ ), .C(\us20\/_0284_ ), .D(\us20\/_0285_ ), .X(\us20\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1090_ ( .A(\us20\/_0082_ ), .B(\us20\/_0027_ ), .X(\us20\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1091_ ( .A(\us20\/_0129_ ), .B(\us20\/_0027_ ), .X(\us20\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_1092_ ( .A(\us20\/_0287_ ), .B(\us20\/_0288_ ), .Y(\us20\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1093_ ( .A1(\us20\/_0752_ ), .A2(\us20\/_0683_ ), .B1(\us20\/_0093_ ), .B2(\us20\/_0247_ ), .Y(\us20\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1094_ ( .A1(\us20\/_0092_ ), .A2(\us20\/_0575_ ), .B1(\us20\/_0292_ ), .Y(\us20\/_0291_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_1095_ ( .A(\us20\/_0054_ ), .X(\us20\/_0292_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1096_ ( .A1(\us20\/_0218_ ), .A2(\us20\/_0672_ ), .B1(\us20\/_0084_ ), .B2(\us20\/_0292_ ), .Y(\us20\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1097_ ( .A(\us20\/_0289_ ), .B(\us20\/_0290_ ), .C(\us20\/_0291_ ), .D(\us20\/_0294_ ), .X(\us20\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1098_ ( .A(\us20\/_0750_ ), .B(\us20\/_0193_ ), .X(\us20\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1099_ ( .A(\us20\/_0705_ ), .B(\us20\/_0380_ ), .X(\us20\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1100_ ( .A(\us20\/_0752_ ), .B(\us20\/_0129_ ), .Y(\us20\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us20/_1101_ ( .A(\us20\/_0296_ ), .B(\us20\/_0297_ ), .C_N(\us20\/_0298_ ), .Y(\us20\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1102_ ( .A(\us20\/_0089_ ), .B(\us20\/_0532_ ), .Y(\us20\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1103_ ( .A(\sa20\[2\] ), .Y(\us20\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \us20/_1104_ ( .A(\us20\/_0301_ ), .B(\sa20\[3\] ), .C(\us20\/_0118_ ), .Y(\us20\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1105_ ( .A(\us20\/_0072_ ), .B(\us20\/_0302_ ), .X(\us20\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1106_ ( .A(\us20\/_0303_ ), .Y(\us20\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1107_ ( .A(\us20\/_0147_ ), .B(\us20\/_0302_ ), .Y(\us20\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1108_ ( .A(\us20\/_0299_ ), .B(\us20\/_0300_ ), .C(\us20\/_0305_ ), .D(\us20\/_0306_ ), .X(\us20\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1109_ ( .A(\us20\/_0278_ ), .B(\us20\/_0286_ ), .C(\us20\/_0295_ ), .D(\us20\/_0307_ ), .X(\us20\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us20/_1110_ ( .A(\us20\/_0228_ ), .B(\us20\/_0265_ ), .C(\us20\/_0308_ ), .Y(\us20\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1111_ ( .A(\us20\/_0235_ ), .Y(\us20\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1112_ ( .A(\us20\/_0478_ ), .B(\us20\/_0640_ ), .X(\us20\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1113_ ( .A(\us20\/_0310_ ), .Y(\us20\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1114_ ( .A(\us20\/_0022_ ), .B(\us20\/_0218_ ), .Y(\us20\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1115_ ( .A(\us20\/_0218_ ), .B(\us20\/_0032_ ), .Y(\us20\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1116_ ( .A(\us20\/_0309_ ), .B(\us20\/_0311_ ), .C(\us20\/_0312_ ), .D(\us20\/_0313_ ), .X(\us20\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1117_ ( .A(\us20\/_0218_ ), .B(\us20\/_0064_ ), .Y(\us20\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1118_ ( .A(\us20\/_0218_ ), .B(\us20\/_0683_ ), .Y(\us20\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1119_ ( .A(\us20\/_0315_ ), .B(\us20\/_0316_ ), .C(\us20\/_0317_ ), .D(\us20\/_0253_ ), .X(\us20\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1120_ ( .A(\us20\/_0047_ ), .B(\us20\/_0304_ ), .Y(\us20\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1121_ ( .A(\us20\/_0586_ ), .B(\us20\/_0162_ ), .Y(\us20\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1122_ ( .A(\us20\/_0319_ ), .B(\us20\/_0320_ ), .Y(\us20\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_1123_ ( .A(\us20\/_0321_ ), .B(\us20\/_0238_ ), .Y(\us20\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1124_ ( .A(\us20\/_0304_ ), .B(\us20\/_0062_ ), .Y(\us20\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_1125_ ( .A(\us20\/_0251_ ), .X(\us20\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1126_ ( .A1(\us20\/_0324_ ), .A2(\us20\/_0084_ ), .B1(\us20\/_0255_ ), .Y(\us20\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1127_ ( .A1(\us20\/_0050_ ), .A2(\us20\/_0216_ ), .B1(\us20\/_0109_ ), .C1(\us20\/_0255_ ), .Y(\us20\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1128_ ( .A(\us20\/_0322_ ), .B(\us20\/_0323_ ), .C(\us20\/_0326_ ), .D(\us20\/_0327_ ), .X(\us20\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1129_ ( .A1(\us20\/_0733_ ), .A2(\us20\/_0279_ ), .A3(\us20\/_0058_ ), .B1(\us20\/_0292_ ), .Y(\us20\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_1130_ ( .A(\us20\/_0047_ ), .X(\us20\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1131_ ( .A(\us20\/_0330_ ), .B(\us20\/_0292_ ), .Y(\us20\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1132_ ( .A(\us20\/_0054_ ), .B(\us20\/_0045_ ), .Y(\us20\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1133_ ( .A(\us20\/_0329_ ), .B(\us20\/_0331_ ), .C(\us20\/_0284_ ), .D(\us20\/_0332_ ), .X(\us20\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us20/_1134_ ( .A1(\us20\/_0543_ ), .A2(\us20\/_0216_ ), .B1(\us20\/_0532_ ), .C1(\us20\/_0060_ ), .X(\us20\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1135_ ( .A(\us20\/_0084_ ), .B(\us20\/_0060_ ), .Y(\us20\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1136_ ( .A(\us20\/_0324_ ), .B(\us20\/_0060_ ), .Y(\us20\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1137_ ( .A(\us20\/_0335_ ), .B(\us20\/_0337_ ), .Y(\us20\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1138_ ( .A1(\us20\/_0276_ ), .A2(\us20\/_0060_ ), .B1(\us20\/_0334_ ), .C1(\us20\/_0338_ ), .Y(\us20\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1139_ ( .A(\us20\/_0318_ ), .B(\us20\/_0328_ ), .C(\us20\/_0333_ ), .D(\us20\/_0339_ ), .X(\us20\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us20/_1140_ ( .A1(\us20\/_0746_ ), .A2(\us20\/_0134_ ), .B1(\us20\/_0128_ ), .X(\us20\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us20/_1141_ ( .A_N(\us20\/_0086_ ), .B(\us20\/_0128_ ), .X(\us20\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1142_ ( .A(\us20\/_0079_ ), .B(\us20\/_0124_ ), .X(\us20\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_1143_ ( .A(\us20\/_0126_ ), .B(\us20\/_0343_ ), .Y(\us20\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us20/_1144_ ( .A(\us20\/_0341_ ), .B(\us20\/_0342_ ), .C_N(\us20\/_0344_ ), .Y(\us20\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1146_ ( .A1(\us20\/_0193_ ), .A2(\us20\/_0092_ ), .A3(\us20\/_0330_ ), .B1(\us20\/_0147_ ), .Y(\us20\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1147_ ( .A1(\us20\/_0130_ ), .A2(\us20\/_0084_ ), .A3(\us20\/_0134_ ), .B1(\us20\/_0139_ ), .Y(\us20\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1148_ ( .A1(\us20\/_0144_ ), .A2(\us20\/_0608_ ), .A3(\us20\/_0092_ ), .B1(\us20\/_0139_ ), .Y(\us20\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1149_ ( .A(\us20\/_0345_ ), .B(\us20\/_0348_ ), .C(\us20\/_0349_ ), .D(\us20\/_0350_ ), .X(\us20\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us20/_1150_ ( .A(\us20\/_0150_ ), .B(\us20\/_0194_ ), .C(\us20\/_0543_ ), .X(\us20\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us20/_1151_ ( .A(\us20\/_0277_ ), .SLEEP(\us20\/_0352_ ), .X(\us20\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us20/_1152_ ( .A1(\us20\/_0268_ ), .A2(\us20\/_0171_ ), .B1(\us20\/_0157_ ), .Y(\us20\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us20/_1153_ ( .A(\us20\/_0161_ ), .X(\us20\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1154_ ( .A1(\us20\/_0279_ ), .A2(\us20\/_0084_ ), .B1(\us20\/_0355_ ), .Y(\us20\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1155_ ( .A1(\us20\/_0020_ ), .A2(\us20\/_0193_ ), .A3(\us20\/_0091_ ), .B1(\us20\/_0355_ ), .Y(\us20\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1156_ ( .A(\us20\/_0353_ ), .B(\us20\/_0354_ ), .C(\us20\/_0356_ ), .D(\us20\/_0357_ ), .X(\us20\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1157_ ( .A(\us20\/_0111_ ), .B(\us20\/_0586_ ), .X(\us20\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1158_ ( .A(\us20\/_0360_ ), .Y(\us20\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us20/_1159_ ( .A1(\us20\/_0119_ ), .A2(\us20\/_0120_ ), .B1(\us20\/_0230_ ), .C1(\us20\/_0361_ ), .X(\us20\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1160_ ( .A1(\us20\/_0672_ ), .A2(\us20\/_0251_ ), .A3(\us20\/_0134_ ), .B1(\us20\/_0114_ ), .Y(\us20\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1162_ ( .A1(\us20\/_0035_ ), .A2(\us20\/_0251_ ), .A3(\us20\/_0134_ ), .B1(\us20\/_0099_ ), .Y(\us20\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1163_ ( .A1(\us20\/_0193_ ), .A2(\us20\/_0608_ ), .B1(\us20\/_0099_ ), .Y(\us20\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1164_ ( .A(\us20\/_0362_ ), .B(\us20\/_0363_ ), .C(\us20\/_0365_ ), .D(\us20\/_0366_ ), .X(\us20\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1165_ ( .A1(\us20\/_0575_ ), .A2(\us20\/_0092_ ), .A3(\us20\/_0330_ ), .B1(\us20\/_0089_ ), .Y(\us20\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1166_ ( .A1(\us20\/_0586_ ), .A2(\us20\/_0017_ ), .A3(\us20\/_0330_ ), .B1(\us20\/_0094_ ), .Y(\us20\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \us20/_1167_ ( .A1(\us20\/_0293_ ), .A2(\us20\/_0134_ ), .B1(\us20\/_0089_ ), .Y(\us20\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1168_ ( .A1(\us20\/_0279_ ), .A2(\us20\/_0134_ ), .B1(\us20\/_0094_ ), .Y(\us20\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1169_ ( .A(\us20\/_0368_ ), .B(\us20\/_0370_ ), .C(\us20\/_0371_ ), .D(\us20\/_0372_ ), .X(\us20\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1170_ ( .A(\us20\/_0351_ ), .B(\us20\/_0359_ ), .C(\us20\/_0367_ ), .D(\us20\/_0373_ ), .X(\us20\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1171_ ( .A1(\us20\/_0102_ ), .A2(\us20\/_0347_ ), .B1(\us20\/_0109_ ), .C1(\us20\/_0247_ ), .Y(\us20\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1172_ ( .A1(\us20\/_0102_ ), .A2(\us20\/_0347_ ), .B1(\us20\/_0532_ ), .C1(\us20\/_0247_ ), .Y(\us20\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1173_ ( .A1(\us20\/_0050_ ), .A2(\us20\/_0543_ ), .B1(\us20\/_0380_ ), .C1(\us20\/_0247_ ), .Y(\us20\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1174_ ( .A(\us20\/_0041_ ), .B(\us20\/_0375_ ), .C(\us20\/_0376_ ), .D(\us20\/_0377_ ), .X(\us20\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1175_ ( .A(\us20\/_0047_ ), .B(\us20\/_0750_ ), .X(\us20\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1176_ ( .A(\us20\/_0379_ ), .Y(\us20\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1177_ ( .A(\us20\/_0016_ ), .B(\us20\/_0608_ ), .Y(\us20\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1178_ ( .A(\us20\/_0752_ ), .B(\us20\/_0554_ ), .Y(\us20\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1179_ ( .A1(\us20\/_0107_ ), .A2(\us20\/_0734_ ), .B1(\us20\/_0109_ ), .C1(\us20\/_0016_ ), .Y(\us20\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1180_ ( .A(\us20\/_0381_ ), .B(\us20\/_0382_ ), .C(\us20\/_0383_ ), .D(\us20\/_0384_ ), .X(\us20\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us20/_1181_ ( .A(\us20\/_0086_ ), .B_N(\us20\/_0736_ ), .X(\us20\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1182_ ( .A1(\us20\/_0748_ ), .A2(\us20\/_0134_ ), .B1(\us20\/_0739_ ), .Y(\us20\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1183_ ( .A1(\us20\/_0118_ ), .A2(\us20\/_0543_ ), .B1(\us20\/_0109_ ), .C1(\us20\/_0739_ ), .Y(\us20\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1184_ ( .A1(\us20\/_0102_ ), .A2(\us20\/_0301_ ), .B1(\sa20\[3\] ), .C1(\us20\/_0739_ ), .Y(\us20\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1185_ ( .A(\us20\/_0386_ ), .B(\us20\/_0387_ ), .C(\us20\/_0388_ ), .D(\us20\/_0389_ ), .X(\us20\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1186_ ( .A(\us20\/_0020_ ), .Y(\us20\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1187_ ( .A(\us20\/_0727_ ), .Y(\us20\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1188_ ( .A(\us20\/_0727_ ), .B(\us20\/_0064_ ), .Y(\us20\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1189_ ( .A1(\us20\/_0102_ ), .A2(\us20\/_0734_ ), .B1(\us20\/_0532_ ), .C1(\us20\/_0727_ ), .Y(\us20\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us20/_1190_ ( .A1(\us20\/_0392_ ), .A2(\us20\/_0393_ ), .B1(\us20\/_0394_ ), .C1(\us20\/_0395_ ), .X(\us20\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1191_ ( .A(\us20\/_0378_ ), .B(\us20\/_0385_ ), .C(\us20\/_0390_ ), .D(\us20\/_0396_ ), .X(\us20\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us20/_1192_ ( .A(\us20\/_0340_ ), .B(\us20\/_0374_ ), .C(\us20\/_0397_ ), .Y(\us20\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1193_ ( .A(\us20\/_0077_ ), .B(\us20\/_0129_ ), .X(\us20\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_1194_ ( .A(\us20\/_0398_ ), .B(\us20\/_0239_ ), .Y(\us20\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1195_ ( .A(\us20\/_0022_ ), .B(\us20\/_0111_ ), .X(\us20\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us20/_1196_ ( .A_N(\us20\/_0400_ ), .B(\us20\/_0231_ ), .Y(\us20\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us20/_1197_ ( .A(\us20\/_0399_ ), .SLEEP(\us20\/_0402_ ), .X(\us20\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_1198_ ( .A(\us20\/_0746_ ), .B(\us20\/_0251_ ), .Y(\us20\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us20/_1199_ ( .A_N(\us20\/_0404_ ), .B(\us20\/_0752_ ), .Y(\us20\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us20/_1200_ ( .A(\us20\/_0467_ ), .B(\us20\/_0194_ ), .C(\us20\/_0694_ ), .X(\us20\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us20/_1201_ ( .A_N(\us20\/_0175_ ), .B(\us20\/_0406_ ), .X(\us20\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1202_ ( .A(\us20\/_0407_ ), .Y(\us20\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1203_ ( .A1(\us20\/_0094_ ), .A2(\us20\/_0197_ ), .B1(\us20\/_0114_ ), .B2(\us20\/_0640_ ), .Y(\us20\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1204_ ( .A(\us20\/_0403_ ), .B(\us20\/_0405_ ), .C(\us20\/_0408_ ), .D(\us20\/_0409_ ), .X(\us20\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1205_ ( .A(\us20\/_0030_ ), .B(\us20\/_0150_ ), .Y(\us20\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us20/_1206_ ( .A_N(\us20\/_0169_ ), .B(\us20\/_0289_ ), .C(\us20\/_0411_ ), .X(\us20\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us20/_1207_ ( .A1(\us20\/_0467_ ), .A2(\us20\/_0151_ ), .B1(\us20\/_0140_ ), .C1(\us20\/_0129_ ), .X(\us20\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1208_ ( .A1(\us20\/_0608_ ), .A2(\us20\/_0099_ ), .B1(\us20\/_0037_ ), .C1(\us20\/_0414_ ), .Y(\us20\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1209_ ( .A(\us20\/_0738_ ), .Y(\us20\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1210_ ( .A(\us20\/_0586_ ), .B(\us20\/_0736_ ), .Y(\us20\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1211_ ( .A1(\us20\/_0194_ ), .A2(\us20\/_0038_ ), .B1(\us20\/_0118_ ), .C1(\us20\/_0153_ ), .Y(\us20\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us20/_1212_ ( .A1(\us20\/_0416_ ), .A2(\us20\/_0117_ ), .B1(\us20\/_0417_ ), .C1(\us20\/_0418_ ), .X(\us20\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1213_ ( .A(\us20\/_0077_ ), .B(\us20\/_0035_ ), .X(\us20\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1214_ ( .A(\us20\/_0672_ ), .B(\us20\/_0124_ ), .Y(\us20\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1215_ ( .A(\us20\/_0030_ ), .B(\us20\/_0137_ ), .Y(\us20\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1216_ ( .A(\us20\/_0072_ ), .B(\us20\/_0732_ ), .Y(\us20\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us20/_1217_ ( .A_N(\us20\/_0420_ ), .B(\us20\/_0421_ ), .C(\us20\/_0422_ ), .D(\us20\/_0424_ ), .X(\us20\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1218_ ( .A(\us20\/_0413_ ), .B(\us20\/_0415_ ), .C(\us20\/_0419_ ), .D(\us20\/_0425_ ), .X(\us20\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us20/_1219_ ( .A(\us20\/_0355_ ), .B(\us20\/_0102_ ), .C(\us20\/_0109_ ), .Y(\us20\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1220_ ( .A(\us20\/_0077_ ), .B(\us20\/_0017_ ), .X(\us20\/_0428_ ) );
sky130_fd_sc_hd__and2_1 \us20/_1221_ ( .A(\us20\/_0077_ ), .B(\us20\/_0554_ ), .X(\us20\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us20/_1222_ ( .A1(\us20\/_0050_ ), .A2(\us20\/_0216_ ), .B1(\us20\/_0380_ ), .C1(\us20\/_0078_ ), .X(\us20\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us20/_1223_ ( .A(\us20\/_0428_ ), .B(\us20\/_0429_ ), .C(\us20\/_0430_ ), .Y(\us20\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us20/_1224_ ( .A_N(\us20\/_0209_ ), .B(\us20\/_0431_ ), .X(\us20\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us20/_1225_ ( .A1(\us20\/_0215_ ), .A2(\us20\/_0404_ ), .B1(\us20\/_0427_ ), .C1(\us20\/_0432_ ), .X(\us20\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1226_ ( .A(\us20\/_0043_ ), .B(\us20\/_0058_ ), .Y(\us20\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1227_ ( .A(\us20\/_0195_ ), .B(\us20\/_0233_ ), .C(\us20\/_0320_ ), .D(\us20\/_0435_ ), .X(\us20\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1228_ ( .A(\us20\/_0261_ ), .B(\us20\/_0738_ ), .Y(\us20\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1229_ ( .A1(\us20\/_0218_ ), .A2(\us20\/_0640_ ), .B1(\us20\/_0261_ ), .B2(\us20\/_0292_ ), .Y(\us20\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1230_ ( .A(\us20\/_0436_ ), .B(\us20\/_0394_ ), .C(\us20\/_0437_ ), .D(\us20\/_0438_ ), .X(\us20\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1231_ ( .A(\us20\/_0410_ ), .B(\us20\/_0426_ ), .C(\us20\/_0433_ ), .D(\us20\/_0439_ ), .X(\us20\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us20/_1232_ ( .A(\us20\/_0135_ ), .SLEEP(\us20\/_0273_ ), .X(\us20\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1233_ ( .A1(\us20\/_0279_ ), .A2(\us20\/_0134_ ), .B1(\us20\/_0099_ ), .Y(\us20\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1234_ ( .A(\us20\/_0441_ ), .B(\us20\/_0164_ ), .C(\us20\/_0270_ ), .D(\us20\/_0442_ ), .X(\us20\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1235_ ( .A(\us20\/_0051_ ), .B(\us20\/_0672_ ), .Y(\us20\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1236_ ( .A(\us20\/_0051_ ), .B(\us20\/_0271_ ), .Y(\us20\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1237_ ( .A(\us20\/_0444_ ), .B(\us20\/_0446_ ), .X(\us20\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1238_ ( .A(\us20\/_0193_ ), .B(\us20\/_0304_ ), .X(\us20\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1239_ ( .A(\us20\/_0448_ ), .Y(\us20\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1240_ ( .A(\us20\/_0162_ ), .B(\us20\/_0130_ ), .X(\us20\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1241_ ( .A(\us20\/_0450_ ), .Y(\us20\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1242_ ( .A1(\us20\/_0129_ ), .A2(\us20\/_0554_ ), .B1(\us20\/_0043_ ), .Y(\us20\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1243_ ( .A(\us20\/_0447_ ), .B(\us20\/_0449_ ), .C(\us20\/_0451_ ), .D(\us20\/_0452_ ), .X(\us20\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1244_ ( .A(\us20\/_0292_ ), .B(\us20\/_0064_ ), .Y(\us20\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us20/_1245_ ( .A_N(\us20\/_0248_ ), .B(\us20\/_0454_ ), .C(\us20\/_0254_ ), .D(\us20\/_0256_ ), .X(\us20\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1246_ ( .A1(\us20\/_0330_ ), .A2(\us20\/_0099_ ), .B1(\us20\/_0134_ ), .B2(\us20\/_0705_ ), .Y(\us20\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1247_ ( .A1(\us20\/_0748_ ), .A2(\us20\/_0738_ ), .B1(\us20\/_0092_ ), .B2(\us20\/_0752_ ), .Y(\us20\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1248_ ( .A1(\us20\/_0072_ ), .A2(\us20\/_0035_ ), .B1(\us20\/_0748_ ), .B2(\us20\/_0292_ ), .Y(\us20\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1249_ ( .A1(\us20\/_0748_ ), .A2(\us20\/_0251_ ), .B1(\us20\/_0247_ ), .Y(\us20\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1250_ ( .A(\us20\/_0457_ ), .B(\us20\/_0458_ ), .C(\us20\/_0459_ ), .D(\us20\/_0460_ ), .X(\us20\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1251_ ( .A(\us20\/_0443_ ), .B(\us20\/_0453_ ), .C(\us20\/_0455_ ), .D(\us20\/_0461_ ), .X(\us20\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1252_ ( .A(\us20\/_0705_ ), .B(\us20\/_0079_ ), .X(\us20\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1253_ ( .A(\us20\/_0586_ ), .B(\us20\/_0124_ ), .Y(\us20\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1254_ ( .A(\us20\/_0218_ ), .B(\us20\/_0746_ ), .Y(\us20\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us20/_1255_ ( .A_N(\us20\/_0463_ ), .B(\us20\/_0464_ ), .C(\us20\/_0465_ ), .X(\us20\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us20/_1256_ ( .A1(\us20\/_0271_ ), .A2(\us20\/_0072_ ), .B1(\us20\/_0142_ ), .B2(\us20\/_0027_ ), .X(\us20\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1257_ ( .A1(\us20\/_0144_ ), .A2(\us20\/_0099_ ), .B1(\us20\/_0360_ ), .C1(\us20\/_0468_ ), .Y(\us20\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us20/_1258_ ( .A1(\us20\/_0672_ ), .A2(\us20\/_0251_ ), .B1(\us20\/_0218_ ), .X(\us20\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1259_ ( .A1(\us20\/_0575_ ), .A2(\us20\/_0292_ ), .B1(\us20\/_0379_ ), .C1(\us20\/_0470_ ), .Y(\us20\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1260_ ( .A(\us20\/_0466_ ), .B(\us20\/_0469_ ), .C(\us20\/_0471_ ), .D(\us20\/_0305_ ), .X(\us20\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us20/_1261_ ( .A1(\us20\/_0247_ ), .A2(\us20\/_0683_ ), .B1(\us20\/_0324_ ), .B2(\us20\/_0292_ ), .X(\us20\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1262_ ( .A(\us20\/_0084_ ), .B(\us20\/_0099_ ), .X(\us20\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us20/_1263_ ( .A1(\us20\/_0092_ ), .A2(\us20\/_0247_ ), .B1(\us20\/_0474_ ), .X(\us20\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us20/_1264_ ( .A(\us20\/_0075_ ), .B(\us20\/_0473_ ), .C(\us20\/_0475_ ), .Y(\us20\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1265_ ( .A1(\us20\/_0279_ ), .A2(\us20\/_0255_ ), .B1(\us20\/_0084_ ), .B2(\us20\/_0060_ ), .Y(\us20\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1266_ ( .A1(\us20\/_0093_ ), .A2(\us20\/_0292_ ), .B1(\us20\/_0134_ ), .B2(\us20\/_0114_ ), .Y(\us20\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1267_ ( .A1(\us20\/_0161_ ), .A2(\us20\/_0032_ ), .B1(\us20\/_0324_ ), .B2(\us20\/_0147_ ), .Y(\us20\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1268_ ( .A1(\us20\/_0054_ ), .A2(\us20\/_0732_ ), .B1(\us20\/_0748_ ), .B2(\us20\/_0304_ ), .Y(\us20\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1269_ ( .A(\us20\/_0477_ ), .B(\us20\/_0479_ ), .C(\us20\/_0480_ ), .D(\us20\/_0481_ ), .X(\us20\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1270_ ( .A(\us20\/_0161_ ), .B(\us20\/_0064_ ), .Y(\us20\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us20/_1271_ ( .A(\us20\/_0732_ ), .B(\us20\/_0123_ ), .C(\us20\/_0467_ ), .Y(\us20\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1272_ ( .A(\us20\/_0483_ ), .B(\us20\/_0484_ ), .Y(\us20\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1273_ ( .A(\us20\/_0297_ ), .Y(\us20\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us20/_1274_ ( .A_N(\us20\/_0485_ ), .B(\us20\/_0181_ ), .C(\us20\/_0486_ ), .D(\us20\/_0386_ ), .X(\us20\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1275_ ( .A(\us20\/_0472_ ), .B(\us20\/_0476_ ), .C(\us20\/_0482_ ), .D(\us20\/_0487_ ), .X(\us20\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \us20/_1276_ ( .A(\us20\/_0440_ ), .B(\us20\/_0462_ ), .C(\us20\/_0488_ ), .Y(\us20\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1277_ ( .A(\us20\/_0403_ ), .B(\us20\/_0230_ ), .C(\us20\/_0451_ ), .D(\us20\/_0361_ ), .X(\us20\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1278_ ( .A1(\us20\/_0118_ ), .A2(\us20\/_0050_ ), .B1(\us20\/_0109_ ), .C1(\us20\/_0139_ ), .Y(\us20\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1279_ ( .A(\us20\/_0447_ ), .B(\us20\/_0437_ ), .C(\us20\/_0491_ ), .D(\us20\/_0427_ ), .X(\us20\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1280_ ( .A1(\us20\/_0084_ ), .A2(\us20\/_0255_ ), .B1(\us20\/_0608_ ), .B2(\us20\/_0247_ ), .Y(\us20\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1281_ ( .A1(\us20\/_0144_ ), .A2(\us20\/_0147_ ), .B1(\us20\/_0355_ ), .B2(\us20\/_0093_ ), .Y(\us20\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1282_ ( .A1(\us20\/_0705_ ), .A2(\us20\/_0279_ ), .B1(\us20\/_0330_ ), .B2(\us20\/_0247_ ), .Y(\us20\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1283_ ( .A1(\us20\/_0279_ ), .A2(\us20\/_0084_ ), .B1(\us20\/_0114_ ), .Y(\us20\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1284_ ( .A(\us20\/_0493_ ), .B(\us20\/_0494_ ), .C(\us20\/_0495_ ), .D(\us20\/_0496_ ), .X(\us20\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1285_ ( .A1(\us20\/_0134_ ), .A2(\us20\/_0137_ ), .B1(\us20\/_0355_ ), .B2(\us20\/_0575_ ), .Y(\us20\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1286_ ( .A1(\us20\/_0099_ ), .A2(\us20\/_0733_ ), .B1(\us20\/_0093_ ), .B2(\us20\/_0218_ ), .Y(\us20\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1287_ ( .A(\us20\/_0147_ ), .B(\us20\/_0640_ ), .Y(\us20\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1288_ ( .A1(\us20\/_0153_ ), .A2(\us20\/_0292_ ), .B1(\us20\/_0748_ ), .Y(\us20\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1289_ ( .A(\us20\/_0498_ ), .B(\us20\/_0500_ ), .C(\us20\/_0501_ ), .D(\us20\/_0502_ ), .X(\us20\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1290_ ( .A(\us20\/_0490_ ), .B(\us20\/_0492_ ), .C(\us20\/_0497_ ), .D(\us20\/_0503_ ), .X(\us20\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us20/_1291_ ( .A_N(\us20\/_0275_ ), .B(\us20\/_0705_ ), .X(\us20\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1292_ ( .A(\us20\/_0505_ ), .Y(\us20\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1293_ ( .A(\us20\/_0380_ ), .B(\us20\/_0347_ ), .X(\us20\/_0507_ ) );
sky130_fd_sc_hd__o21ai_1 \us20/_1294_ ( .A1(\us20\/_0507_ ), .A2(\us20\/_0093_ ), .B1(\us20\/_0292_ ), .Y(\us20\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1295_ ( .A(\us20\/_0322_ ), .B(\us20\/_0277_ ), .C(\us20\/_0506_ ), .D(\us20\/_0508_ ), .X(\us20\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1296_ ( .A(\us20\/_0084_ ), .B(\us20\/_0705_ ), .X(\us20\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1297_ ( .A1(\us20\/_0733_ ), .A2(\us20\/_0114_ ), .B1(\us20\/_0429_ ), .C1(\us20\/_0511_ ), .Y(\us20\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_1298_ ( .A(\us20\/_0019_ ), .B(\us20\/_0024_ ), .Y(\us20\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1299_ ( .A(\us20\/_0512_ ), .B(\us20\/_0513_ ), .C(\us20\/_0742_ ), .D(\us20\/_0306_ ), .X(\us20\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1300_ ( .A1(\us20\/_0532_ ), .A2(\us20\/_0089_ ), .B1(\us20\/_0154_ ), .C1(\us20\/_0169_ ), .Y(\us20\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us20/_1301_ ( .A1(\us20\/_0749_ ), .A2(\us20\/_0026_ ), .B1(\us20\/_0069_ ), .C1(\us20\/_0032_ ), .X(\us20\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us20/_1302_ ( .A1(\us20\/_0324_ ), .A2(\us20\/_0355_ ), .B1(\us20\/_0330_ ), .B2(\us20\/_0727_ ), .X(\us20\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us20/_1303_ ( .A(\us20\/_0133_ ), .B(\us20\/_0516_ ), .C(\us20\/_0517_ ), .Y(\us20\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1304_ ( .A(\us20\/_0509_ ), .B(\us20\/_0514_ ), .C(\us20\/_0515_ ), .D(\us20\/_0518_ ), .X(\us20\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1305_ ( .A(\us20\/_0746_ ), .B(\us20\/_0072_ ), .Y(\us20\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1306_ ( .A1(\us20\/_0082_ ), .A2(\us20\/_0070_ ), .B1(\us20\/_0043_ ), .B2(\us20\/_0193_ ), .Y(\us20\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1307_ ( .A(\us20\/_0311_ ), .B(\us20\/_0520_ ), .C(\us20\/_0332_ ), .D(\us20\/_0522_ ), .X(\us20\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1308_ ( .A(\us20\/_0129_ ), .B(\us20\/_0218_ ), .X(\us20\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_1309_ ( .A(\us20\/_0235_ ), .B(\us20\/_0524_ ), .Y(\us20\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us20/_1310_ ( .A(\us20\/_0081_ ), .B(\us20\/_0085_ ), .Y(\us20\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1311_ ( .A1(\us20\/_0051_ ), .A2(\us20\/_0045_ ), .B1(\us20\/_0130_ ), .B2(\us20\/_0094_ ), .Y(\us20\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1312_ ( .A(\us20\/_0523_ ), .B(\us20\/_0525_ ), .C(\us20\/_0526_ ), .D(\us20\/_0527_ ), .X(\us20\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us20/_1313_ ( .A_N(\us20\/_0250_ ), .B(\us20\/_0521_ ), .Y(\us20\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1314_ ( .A(\us20\/_0128_ ), .B(\us20\/_0020_ ), .X(\us20\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1315_ ( .A(\us20\/_0530_ ), .Y(\us20\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1316_ ( .A(\us20\/_0099_ ), .B(\us20\/_0058_ ), .X(\us20\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1317_ ( .A(\us20\/_0533_ ), .Y(\us20\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us20/_1318_ ( .A_N(\us20\/_0529_ ), .B(\us20\/_0531_ ), .C(\us20\/_0534_ ), .D(\us20\/_0192_ ), .X(\us20\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1319_ ( .A(\us20\/_0434_ ), .B(\us20\/_0078_ ), .X(\us20\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us20/_1320_ ( .A1(\us20\/_0750_ ), .A2(\us20\/_0079_ ), .B1(\us20\/_0129_ ), .B2(\us20\/_0705_ ), .X(\us20\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1321_ ( .A1(\us20\/_0161_ ), .A2(\us20\/_0032_ ), .B1(\us20\/_0536_ ), .C1(\us20\/_0537_ ), .Y(\us20\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us20/_1322_ ( .A1(\us20\/_0746_ ), .A2(\us20\/_0162_ ), .B1(\us20\/_0079_ ), .B2(\us20\/_0043_ ), .X(\us20\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1323_ ( .A1(\us20\/_0093_ ), .A2(\us20\/_0247_ ), .B1(\us20\/_0240_ ), .C1(\us20\/_0539_ ), .Y(\us20\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1324_ ( .A(\us20\/_0434_ ), .B(\us20\/_0043_ ), .X(\us20\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us20/_1325_ ( .A1(\us20\/_0142_ ), .A2(\us20\/_0150_ ), .B1(\us20\/_0022_ ), .B2(\us20\/_0137_ ), .X(\us20\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1326_ ( .A1(\us20\/_0279_ ), .A2(\us20\/_0051_ ), .B1(\us20\/_0541_ ), .C1(\us20\/_0542_ ), .Y(\us20\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1327_ ( .A(\us20\/_0159_ ), .B(\us20\/_0035_ ), .X(\us20\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us20/_1328_ ( .A1(\us20\/_0271_ ), .A2(\us20\/_0434_ ), .B1(\us20\/_0027_ ), .X(\us20\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1329_ ( .A1(\us20\/_0091_ ), .A2(\us20\/_0128_ ), .B1(\us20\/_0545_ ), .C1(\us20\/_0546_ ), .Y(\us20\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1330_ ( .A(\us20\/_0538_ ), .B(\us20\/_0540_ ), .C(\us20\/_0544_ ), .D(\us20\/_0547_ ), .X(\us20\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1331_ ( .A(\us20\/_0099_ ), .B(\us20\/_0193_ ), .X(\us20\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us20/_1332_ ( .A(\us20\/_0549_ ), .B(\us20\/_0186_ ), .C(\us20\/_0187_ ), .Y(\us20\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1333_ ( .A(\us20\/_0062_ ), .B(\us20\/_0347_ ), .C(\us20\/_0749_ ), .D(\us20\/_0694_ ), .X(\us20\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1334_ ( .A1(\us20\/_0130_ ), .A2(\us20\/_0218_ ), .B1(\us20\/_0551_ ), .C1(\us20\/_0101_ ), .Y(\us20\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1335_ ( .A(\us20\/_0139_ ), .B(\us20\/_0640_ ), .Y(\us20\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1336_ ( .A1(\us20\/_0752_ ), .A2(\us20\/_0672_ ), .B1(\us20\/_0084_ ), .B2(\us20\/_0099_ ), .Y(\us20\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1337_ ( .A(\us20\/_0550_ ), .B(\us20\/_0552_ ), .C(\us20\/_0553_ ), .D(\us20\/_0555_ ), .X(\us20\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1338_ ( .A(\us20\/_0528_ ), .B(\us20\/_0535_ ), .C(\us20\/_0548_ ), .D(\us20\/_0556_ ), .X(\us20\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us20/_1339_ ( .A(\us20\/_0504_ ), .B(\us20\/_0519_ ), .C(\us20\/_0557_ ), .Y(\us20\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1340_ ( .A(\us20\/_0054_ ), .B(\us20\/_0507_ ), .X(\us20\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us20/_1341_ ( .A_N(\us20\/_0558_ ), .B(\us20\/_0408_ ), .C(\us20\/_0451_ ), .D(\us20\/_0452_ ), .X(\us20\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1342_ ( .A(\us20\/_0549_ ), .Y(\us20\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1343_ ( .A(\us20\/_0559_ ), .B(\us20\/_0403_ ), .C(\us20\/_0560_ ), .D(\us20\/_0371_ ), .X(\us20\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1344_ ( .A(\us20\/_0181_ ), .B(\us20\/_0178_ ), .X(\us20\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1345_ ( .A(\us20\/_0562_ ), .B(\us20\/_0552_ ), .C(\us20\/_0553_ ), .D(\us20\/_0555_ ), .X(\us20\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1346_ ( .A(\us20\/_0247_ ), .B(\us20\/_0020_ ), .Y(\us20\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1347_ ( .A(\us20\/_0051_ ), .B(\us20\/_0130_ ), .X(\us20\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1348_ ( .A(\us20\/_0566_ ), .Y(\us20\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1349_ ( .A(\us20\/_0159_ ), .B(\us20\/_0423_ ), .X(\us20\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1350_ ( .A1(\us20\/_0752_ ), .A2(\us20\/_0640_ ), .B1(\us20\/_0568_ ), .B2(\us20\/_0175_ ), .Y(\us20\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1351_ ( .A(\us20\/_0076_ ), .B(\us20\/_0565_ ), .C(\us20\/_0567_ ), .D(\us20\/_0569_ ), .X(\us20\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us20/_1352_ ( .A1(\us20\/_0035_ ), .A2(\us20\/_0142_ ), .B1(\us20\/_0161_ ), .X(\us20\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1353_ ( .A(\us20\/_0099_ ), .B(\us20\/_0672_ ), .Y(\us20\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us20/_1354_ ( .A(\us20\/_0420_ ), .B(\us20\/_0571_ ), .C_N(\us20\/_0572_ ), .Y(\us20\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1355_ ( .A(\us20\/_0051_ ), .B(\us20\/_0746_ ), .Y(\us20\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1356_ ( .A(\us20\/_0574_ ), .B(\us20\/_0319_ ), .C(\us20\/_0320_ ), .D(\us20\/_0411_ ), .X(\us20\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1357_ ( .A(\us20\/_0736_ ), .B(\us20\/_0035_ ), .Y(\us20\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1358_ ( .A(\us20\/_0736_ ), .B(\us20\/_0030_ ), .Y(\us20\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1359_ ( .A(\us20\/_0298_ ), .B(\us20\/_0208_ ), .C(\us20\/_0577_ ), .D(\us20\/_0578_ ), .X(\us20\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1360_ ( .A1(\us20\/_0020_ ), .A2(\us20\/_0137_ ), .B1(\us20\/_0261_ ), .B2(\us20\/_0128_ ), .Y(\us20\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1361_ ( .A(\us20\/_0573_ ), .B(\us20\/_0576_ ), .C(\us20\/_0579_ ), .D(\us20\/_0580_ ), .X(\us20\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1362_ ( .A(\us20\/_0561_ ), .B(\us20\/_0563_ ), .C(\us20\/_0570_ ), .D(\us20\/_0581_ ), .X(\us20\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1363_ ( .A(\us20\/_0128_ ), .B(\us20\/_0193_ ), .X(\us20\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1364_ ( .A(\us20\/_0082_ ), .B(\us20\/_0162_ ), .X(\us20\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us20/_1365_ ( .A(\us20\/_0583_ ), .B(\us20\/_0584_ ), .C_N(\us20\/_0437_ ), .Y(\us20\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us20/_1366_ ( .A(\us20\/_0150_ ), .B(\us20\/_0118_ ), .C(\us20\/_0380_ ), .Y(\us20\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us20/_1367_ ( .A_N(\us20\/_0182_ ), .B(\us20\/_0587_ ), .C(\us20\/_0323_ ), .X(\us20\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1368_ ( .A1(\us20\/_0575_ ), .A2(\us20\/_0153_ ), .B1(\us20\/_0727_ ), .B2(\us20\/_0058_ ), .Y(\us20\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1369_ ( .A1(\us20\/_0218_ ), .A2(\us20\/_0064_ ), .B1(\us20\/_0134_ ), .B2(\us20\/_0255_ ), .Y(\us20\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1370_ ( .A(\us20\/_0585_ ), .B(\us20\/_0588_ ), .C(\us20\/_0589_ ), .D(\us20\/_0590_ ), .X(\us20\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us20/_1371_ ( .A1(\us20\/_0091_ ), .A2(\us20\/_0139_ ), .B1(\us20\/_0250_ ), .Y(\us20\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1372_ ( .A1(\us20\/_0092_ ), .A2(\us20\/_0739_ ), .B1(\us20\/_0324_ ), .B2(\us20\/_0247_ ), .Y(\us20\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1373_ ( .A1(\us20\/_0144_ ), .A2(\us20\/_0153_ ), .B1(\us20\/_0683_ ), .B2(\us20\/_0292_ ), .Y(\us20\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1374_ ( .A1(\us20\/_0091_ ), .A2(\us20\/_0218_ ), .B1(\us20\/_0330_ ), .B2(\us20\/_0292_ ), .Y(\us20\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1375_ ( .A(\us20\/_0592_ ), .B(\us20\/_0593_ ), .C(\us20\/_0594_ ), .D(\us20\/_0595_ ), .X(\us20\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1376_ ( .A(\us20\/_0218_ ), .B(\us20\/_0144_ ), .Y(\us20\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1377_ ( .A(\us20\/_0312_ ), .B(\us20\/_0598_ ), .Y(\us20\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1378_ ( .A(\us20\/_0575_ ), .B(\us20\/_0147_ ), .Y(\us20\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1379_ ( .A1(\us20\/_0293_ ), .A2(\us20\/_0137_ ), .B1(\us20\/_0093_ ), .B2(\us20\/_0739_ ), .Y(\us20\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1380_ ( .A1(\us20\/_0734_ ), .A2(\us20\/_0531_ ), .B1(\us20\/_0600_ ), .C1(\us20\/_0601_ ), .Y(\us20\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1381_ ( .A1(\us20\/_0153_ ), .A2(\us20\/_0261_ ), .B1(\us20\/_0599_ ), .C1(\us20\/_0602_ ), .Y(\us20\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1382_ ( .A(\us20\/_0591_ ), .B(\us20\/_0596_ ), .C(\us20\/_0174_ ), .D(\us20\/_0603_ ), .X(\us20\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1383_ ( .A(\us20\/_0247_ ), .B(\us20\/_0144_ ), .Y(\us20\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1384_ ( .A(\us20\/_0113_ ), .B(\us20\/_0017_ ), .Y(\us20\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1385_ ( .A(\us20\/_0381_ ), .B(\us20\/_0605_ ), .C(\us20\/_0361_ ), .D(\us20\/_0606_ ), .X(\us20\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1386_ ( .A1(\us20\/_0016_ ), .A2(\us20\/_0727_ ), .B1(\us20\/_0733_ ), .Y(\us20\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1387_ ( .A1(\us20\/_0586_ ), .A2(\us20\/_0159_ ), .B1(\us20\/_0082_ ), .B2(\us20\/_0750_ ), .Y(\us20\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1388_ ( .A1(\us20\/_0142_ ), .A2(\us20\/_0162_ ), .B1(\us20\/_0079_ ), .B2(\us20\/_0054_ ), .Y(\us20\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1389_ ( .A(\us20\/_0610_ ), .B(\us20\/_0611_ ), .C(\us20\/_0105_ ), .D(\us20\/_0106_ ), .X(\us20\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1390_ ( .A1(\us20\/_0094_ ), .A2(\us20\/_0302_ ), .B1(\us20\/_0324_ ), .B2(\us20\/_0089_ ), .Y(\us20\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1391_ ( .A(\us20\/_0607_ ), .B(\us20\/_0609_ ), .C(\us20\/_0612_ ), .D(\us20\/_0613_ ), .X(\us20\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1392_ ( .A(\us20\/_0041_ ), .B(\us20\/_0170_ ), .X(\us20\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1393_ ( .A(\us20\/_0554_ ), .B(\us20\/_0027_ ), .X(\us20\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1394_ ( .A(\us20\/_0027_ ), .B(\us20\/_0261_ ), .Y(\us20\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us20/_1395_ ( .A_N(\us20\/_0616_ ), .B(\us20\/_0617_ ), .Y(\us20\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1396_ ( .A1(\us20\/_0147_ ), .A2(\us20\/_0302_ ), .B1(\us20\/_0342_ ), .C1(\us20\/_0618_ ), .Y(\us20\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1397_ ( .A(\us20\/_0614_ ), .B(\us20\/_0272_ ), .C(\us20\/_0615_ ), .D(\us20\/_0620_ ), .X(\us20\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us20/_1398_ ( .A(\us20\/_0582_ ), .B(\us20\/_0604_ ), .C(\us20\/_0621_ ), .Y(\us20\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1399_ ( .A1(\us20\/_0084_ ), .A2(\us20\/_0134_ ), .B1(\us20\/_0089_ ), .Y(\us20\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1400_ ( .A1(\us20\/_0144_ ), .A2(\us20\/_0608_ ), .A3(\us20\/_0330_ ), .B1(\us20\/_0089_ ), .Y(\us20\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1401_ ( .A1(\us20\/_0197_ ), .A2(\us20\/_0130_ ), .A3(\us20\/_0110_ ), .B1(\us20\/_0094_ ), .Y(\us20\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1402_ ( .A(\us20\/_0432_ ), .B(\us20\/_0622_ ), .C(\us20\/_0623_ ), .D(\us20\/_0624_ ), .X(\us20\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us20/_1403_ ( .A1(\us20\/_0554_ ), .A2(\us20\/_0017_ ), .A3(\us20\/_0022_ ), .B1(\us20\/_0161_ ), .X(\us20\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us20/_1404_ ( .A_N(\us20\/_0269_ ), .B(\us20\/_0170_ ), .X(\us20\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1405_ ( .A1(\us20\/_0109_ ), .A2(\us20\/_0064_ ), .A3(\us20\/_0733_ ), .B1(\us20\/_0355_ ), .Y(\us20\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us20/_1406_ ( .A_N(\us20\/_0626_ ), .B(\us20\/_0627_ ), .C(\us20\/_0353_ ), .D(\us20\/_0628_ ), .X(\us20\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1407_ ( .A1(\us20\/_0091_ ), .A2(\us20\/_0110_ ), .A3(\us20\/_0176_ ), .B1(\us20\/_0139_ ), .Y(\us20\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1408_ ( .A1(\us20\/_0020_ ), .A2(\us20\/_0261_ ), .B1(\us20\/_0147_ ), .Y(\us20\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1409_ ( .A(\us20\/_0631_ ), .B(\us20\/_0344_ ), .C(\us20\/_0421_ ), .D(\us20\/_0632_ ), .X(\us20\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us20/_1410_ ( .A1(\us20\/_0325_ ), .A2(\us20\/_0734_ ), .B1(\us20\/_0038_ ), .C1(\us20\/_0113_ ), .X(\us20\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1411_ ( .A1(\us20\/_0134_ ), .A2(\us20\/_0114_ ), .B1(\us20\/_0221_ ), .C1(\us20\/_0634_ ), .Y(\us20\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us20/_1412_ ( .A(\us20\/_0119_ ), .B_N(\us20\/_0111_ ), .Y(\us20\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1413_ ( .A1(\us20\/_0032_ ), .A2(\us20\/_0113_ ), .B1(\us20\/_0636_ ), .C1(\us20\/_0400_ ), .Y(\us20\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1414_ ( .A1(\us20\/_0732_ ), .A2(\us20\/_0293_ ), .A3(\us20\/_0251_ ), .B1(\us20\/_0099_ ), .Y(\us20\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1415_ ( .A(\us20\/_0189_ ), .B(\us20\/_0635_ ), .C(\us20\/_0637_ ), .D(\us20\/_0638_ ), .X(\us20\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1416_ ( .A(\us20\/_0625_ ), .B(\us20\/_0630_ ), .C(\us20\/_0633_ ), .D(\us20\/_0639_ ), .X(\us20\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1417_ ( .A(\us20\/_0746_ ), .B(\us20\/_0738_ ), .X(\us20\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1418_ ( .A(\us20\/_0736_ ), .B(\us20\/_0731_ ), .X(\us20\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us20/_1419_ ( .A_N(\us20\/_0643_ ), .B(\us20\/_0577_ ), .Y(\us20\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1420_ ( .A1(\us20\/_0084_ ), .A2(\us20\/_0739_ ), .B1(\us20\/_0642_ ), .C1(\us20\/_0644_ ), .Y(\us20\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1421_ ( .A1(\us20\/_0050_ ), .A2(\us20\/_0543_ ), .B1(\us20\/_0194_ ), .C1(\us20\/_0738_ ), .Y(\us20\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1422_ ( .A(\us20\/_0646_ ), .B(\us20\/_0232_ ), .C(\us20\/_0417_ ), .D(\us20\/_0578_ ), .X(\us20\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1423_ ( .A1(\us20\/_0064_ ), .A2(\us20\/_0733_ ), .B1(\us20\/_0727_ ), .Y(\us20\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1424_ ( .A1(\us20\/_0193_ ), .A2(\us20\/_0276_ ), .B1(\us20\/_0727_ ), .Y(\us20\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1425_ ( .A(\us20\/_0645_ ), .B(\us20\/_0647_ ), .C(\us20\/_0648_ ), .D(\us20\/_0649_ ), .X(\us20\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1426_ ( .A1(\us20\/_0325_ ), .A2(\us20\/_0734_ ), .B1(\us20\/_0038_ ), .C1(\us20\/_0247_ ), .Y(\us20\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1427_ ( .A1(\us20\/_0543_ ), .A2(\us20\/_0216_ ), .B1(\us20\/_0423_ ), .C1(\us20\/_0247_ ), .Y(\us20\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1428_ ( .A(\us20\/_0652_ ), .B(\us20\/_0653_ ), .X(\us20\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1429_ ( .A1(\us20\/_0733_ ), .A2(\us20\/_0748_ ), .A3(\us20\/_0324_ ), .B1(\us20\/_0016_ ), .Y(\us20\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1430_ ( .A1(\us20\/_0640_ ), .A2(\us20\/_0193_ ), .A3(\us20\/_0091_ ), .B1(\us20\/_0016_ ), .Y(\us20\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1431_ ( .A1(\us20\/_0102_ ), .A2(\us20\/_0301_ ), .B1(\sa20\[3\] ), .C1(\us20\/_0247_ ), .Y(\us20\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1432_ ( .A(\us20\/_0654_ ), .B(\us20\/_0655_ ), .C(\us20\/_0656_ ), .D(\us20\/_0657_ ), .X(\us20\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1433_ ( .A1(\us20\/_0118_ ), .A2(\us20\/_0050_ ), .B1(\us20\/_0038_ ), .C1(\us20\/_0478_ ), .Y(\us20\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us20/_1434_ ( .A_N(\us20\/_0250_ ), .B(\us20\/_0465_ ), .C(\us20\/_0659_ ), .X(\us20\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1435_ ( .A1(\us20\/_0683_ ), .A2(\us20\/_0324_ ), .B1(\us20\/_0255_ ), .Y(\us20\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1436_ ( .A1(\us20\/_0032_ ), .A2(\us20\/_0193_ ), .A3(\us20\/_0047_ ), .B1(\us20\/_0255_ ), .Y(\us20\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1437_ ( .A1(\us20\/_0144_ ), .A2(\us20\/_0586_ ), .A3(\us20\/_0047_ ), .B1(\us20\/_0218_ ), .Y(\us20\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1438_ ( .A(\us20\/_0660_ ), .B(\us20\/_0661_ ), .C(\us20\/_0663_ ), .D(\us20\/_0664_ ), .X(\us20\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1439_ ( .A1(\us20\/_0091_ ), .A2(\us20\/_0276_ ), .B1(\us20\/_0060_ ), .Y(\us20\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1440_ ( .A1(\us20\/_0144_ ), .A2(\us20\/_0608_ ), .B1(\us20\/_0292_ ), .Y(\us20\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1441_ ( .A1(\us20\/_0423_ ), .A2(\us20\/_0038_ ), .B1(\us20\/_0102_ ), .C1(\us20\/_0060_ ), .Y(\us20\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1442_ ( .A1(\us20\/_0107_ ), .A2(\us20\/_0734_ ), .B1(\us20\/_0109_ ), .C1(\us20\/_0292_ ), .Y(\us20\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1443_ ( .A(\us20\/_0666_ ), .B(\us20\/_0667_ ), .C(\us20\/_0668_ ), .D(\us20\/_0669_ ), .X(\us20\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1444_ ( .A(\us20\/_0650_ ), .B(\us20\/_0658_ ), .C(\us20\/_0665_ ), .D(\us20\/_0670_ ), .X(\us20\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us20/_1445_ ( .A(\us20\/_0641_ ), .B(\us20\/_0174_ ), .C(\us20\/_0671_ ), .Y(\us20\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us20/_1446_ ( .A(\us20\/_0049_ ), .B(\us20\/_0618_ ), .C_N(\us20\/_0052_ ), .Y(\us20\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us20/_1447_ ( .A(\us20\/_0239_ ), .Y(\us20\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1448_ ( .A(\us20\/_0705_ ), .B(\us20\/_0032_ ), .Y(\us20\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1449_ ( .A1(\us20\/_0054_ ), .A2(\us20\/_0732_ ), .B1(\us20\/_0035_ ), .B2(\us20\/_0705_ ), .Y(\us20\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1450_ ( .A1(\us20\/_0304_ ), .A2(\us20\/_0732_ ), .B1(\us20\/_0047_ ), .B2(\us20\/_0750_ ), .Y(\us20\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1451_ ( .A(\us20\/_0674_ ), .B(\us20\/_0675_ ), .C(\us20\/_0676_ ), .D(\us20\/_0677_ ), .X(\us20\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us20/_1452_ ( .A_N(\us20\/_0584_ ), .B(\us20\/_0283_ ), .X(\us20\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1453_ ( .A(\us20\/_0673_ ), .B(\us20\/_0678_ ), .C(\us20\/_0679_ ), .D(\us20\/_0508_ ), .X(\us20\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1454_ ( .A1(\us20\/_0016_ ), .A2(\us20\/_0733_ ), .B1(\us20\/_0355_ ), .B2(\us20\/_0092_ ), .Y(\us20\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1455_ ( .A(\us20\/_0681_ ), .B(\us20\/_0034_ ), .X(\us20\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us20/_1456_ ( .A1(\us20\/_0330_ ), .A2(\us20\/_0139_ ), .B1(\us20\/_0324_ ), .B2(\us20\/_0089_ ), .X(\us20\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1457_ ( .A1(\us20\/_0146_ ), .A2(\us20\/_0147_ ), .B1(\us20\/_0133_ ), .C1(\us20\/_0684_ ), .Y(\us20\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1458_ ( .A(\us20\/_0113_ ), .B(\us20\/_0251_ ), .Y(\us20\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us20/_1459_ ( .A_N(\us20\/_0463_ ), .B(\us20\/_0686_ ), .C(\us20\/_0383_ ), .D(\us20\/_0464_ ), .X(\us20\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1460_ ( .A1(\us20\/_0051_ ), .A2(\us20\/_0293_ ), .B1(\us20\/_0084_ ), .B2(\us20\/_0705_ ), .Y(\us20\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1461_ ( .A1(\us20\/_0017_ ), .A2(\us20\/_0072_ ), .B1(\us20\/_0134_ ), .B2(\us20\/_0078_ ), .Y(\us20\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1462_ ( .A(\us20\/_0687_ ), .B(\us20\/_0236_ ), .C(\us20\/_0688_ ), .D(\us20\/_0689_ ), .X(\us20\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1463_ ( .A(\us20\/_0680_ ), .B(\us20\/_0682_ ), .C(\us20\/_0685_ ), .D(\us20\/_0690_ ), .X(\us20\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us20/_1464_ ( .A1(\us20\/_0532_ ), .A2(\us20\/_0380_ ), .B1(\us20\/_0102_ ), .C1(\us20\/_0355_ ), .X(\us20\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us20/_1465_ ( .A(\us20\/_0692_ ), .B(\us20\/_0338_ ), .C(\us20\/_0644_ ), .Y(\us20\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1466_ ( .A(\us20\/_0016_ ), .B(\us20\/_0020_ ), .Y(\us20\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1467_ ( .A1(\us20\/_0032_ ), .A2(\us20\/_0137_ ), .B1(\us20\/_0279_ ), .B2(\us20\/_0094_ ), .Y(\us20\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1468_ ( .A1(\us20\/_0575_ ), .A2(\us20\/_0153_ ), .B1(\us20\/_0161_ ), .B2(\us20\/_0293_ ), .Y(\us20\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1469_ ( .A(\us20\/_0259_ ), .B(\us20\/_0695_ ), .C(\us20\/_0696_ ), .D(\us20\/_0697_ ), .X(\us20\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us20/_1470_ ( .A1(\us20\/_0255_ ), .A2(\us20\/_0640_ ), .B1(\us20\/_0016_ ), .B2(\us20\/_0193_ ), .X(\us20\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1471_ ( .A1(\us20\/_0060_ ), .A2(\us20\/_0176_ ), .B1(\us20\/_0699_ ), .C1(\us20\/_0177_ ), .Y(\us20\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1472_ ( .A1(\us20\/_0091_ ), .A2(\us20\/_0218_ ), .B1(\us20\/_0092_ ), .B2(\us20\/_0705_ ), .Y(\us20\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us20/_1473_ ( .A1(\us20\/_0705_ ), .A2(\us20\/_0683_ ), .B1(\us20\/_0093_ ), .B2(\us20\/_0114_ ), .Y(\us20\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us20/_1474_ ( .A1(\us20\/_0683_ ), .A2(\us20\/_0084_ ), .B1(\us20\/_0094_ ), .Y(\us20\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us20/_1475_ ( .A1(\us20\/_0543_ ), .A2(\us20\/_0216_ ), .B1(\us20\/_0038_ ), .C1(\us20\/_0292_ ), .Y(\us20\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1476_ ( .A(\us20\/_0701_ ), .B(\us20\/_0702_ ), .C(\us20\/_0703_ ), .D(\us20\/_0704_ ), .X(\us20\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1477_ ( .A(\us20\/_0693_ ), .B(\us20\/_0698_ ), .C(\us20\/_0700_ ), .D(\us20\/_0706_ ), .X(\us20\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us20/_1478_ ( .A1(\us20\/_0113_ ), .A2(\us20\/_0640_ ), .B1(\us20\/_0099_ ), .B2(\us20\/_0058_ ), .X(\us20\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us20/_1479_ ( .A(\us20\/_0407_ ), .B(\us20\/_0708_ ), .C(\us20\/_0529_ ), .Y(\us20\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1480_ ( .A(\us20\/_0568_ ), .B(\us20\/_0175_ ), .Y(\us20\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us20/_1481_ ( .A1(\us20\/_0247_ ), .A2(\us20\/_0114_ ), .A3(\us20\/_0051_ ), .B1(\us20\/_0130_ ), .Y(\us20\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1482_ ( .A(\us20\/_0709_ ), .B(\us20\/_0550_ ), .C(\us20\/_0710_ ), .D(\us20\/_0711_ ), .X(\us20\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us20/_1483_ ( .A1(\us20\/_0114_ ), .A2(\us20\/_0064_ ), .B1(\us20\/_0261_ ), .B2(\us20\/_0089_ ), .X(\us20\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1484_ ( .A1(\us20\/_0355_ ), .A2(\us20\/_0261_ ), .B1(\us20\/_0198_ ), .C1(\us20\/_0713_ ), .Y(\us20\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1485_ ( .A(\us20\/_0586_ ), .B(\us20\/_0478_ ), .Y(\us20\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us20/_1486_ ( .A_N(\us20\/_0541_ ), .B(\us20\/_0267_ ), .C(\us20\/_0715_ ), .D(\us20\/_0320_ ), .X(\us20\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1487_ ( .A(\us20\/_0586_ ), .B(\us20\/_0070_ ), .Y(\us20\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us20/_1488_ ( .A_N(\us20\/_0211_ ), .B(\us20\/_0155_ ), .C(\us20\/_0202_ ), .D(\us20\/_0718_ ), .X(\us20\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us20/_1489_ ( .A(\us20\/_0150_ ), .B(\us20\/_0216_ ), .C(\us20\/_0380_ ), .Y(\us20\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us20/_1490_ ( .A(\us20\/_0411_ ), .B(\us20\/_0720_ ), .X(\us20\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us20/_1491_ ( .A1(\us20\/_0017_ ), .A2(\us20\/_0022_ ), .B1(\us20\/_0078_ ), .X(\us20\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us20/_1492_ ( .A1(\us20\/_0134_ ), .A2(\us20\/_0738_ ), .B1(\us20\/_0101_ ), .C1(\us20\/_0722_ ), .Y(\us20\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1493_ ( .A(\us20\/_0717_ ), .B(\us20\/_0719_ ), .C(\us20\/_0721_ ), .D(\us20\/_0723_ ), .X(\us20\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us20/_1494_ ( .A(\us20\/_0739_ ), .B(\us20\/_0193_ ), .Y(\us20\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1495_ ( .A(\us20\/_0344_ ), .B(\us20\/_0184_ ), .C(\us20\/_0449_ ), .D(\us20\/_0725_ ), .X(\us20\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us20/_1496_ ( .A(\us20\/_0712_ ), .B(\us20\/_0714_ ), .C(\us20\/_0724_ ), .D(\us20\/_0726_ ), .X(\us20\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \us20/_1497_ ( .A(\us20\/_0691_ ), .B(\us20\/_0707_ ), .C(\us20\/_0728_ ), .Y(\us20\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \us21/_0753_ ( .A(\sa21\[2\] ), .B_N(\sa21\[3\] ), .Y(\us21\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \us21/_0755_ ( .A(\sa21\[1\] ), .B(\sa21\[0\] ), .X(\us21\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us21/_0756_ ( .A(\us21\/_0096_ ), .B(\us21\/_0118_ ), .X(\us21\/_0129_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0757_ ( .A(\sa21\[7\] ), .B(\sa21\[6\] ), .X(\us21\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_0758_ ( .A(\sa21\[4\] ), .B(\sa21\[5\] ), .Y(\us21\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0759_ ( .A(\us21\/_0140_ ), .B(\us21\/_0151_ ), .X(\us21\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0761_ ( .A(\us21\/_0129_ ), .B(\us21\/_0162_ ), .X(\us21\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0762_ ( .A(\us21\/_0096_ ), .X(\us21\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \us21/_0763_ ( .A(\sa21\[1\] ), .B_N(\sa21\[0\] ), .Y(\us21\/_0205_ ) );
sky130_fd_sc_hd__and3_1 \us21/_0765_ ( .A(\us21\/_0162_ ), .B(\us21\/_0194_ ), .C(\us21\/_0205_ ), .X(\us21\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us21/_0766_ ( .A(\us21\/_0183_ ), .SLEEP(\us21\/_0227_ ), .X(\us21\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \us21/_0767_ ( .A(\sa21\[0\] ), .B_N(\sa21\[1\] ), .Y(\us21\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_0768_ ( .A(\sa21\[2\] ), .B(\sa21\[3\] ), .Y(\us21\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0769_ ( .A(\us21\/_0249_ ), .B(\us21\/_0260_ ), .X(\us21\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0771_ ( .A(\us21\/_0271_ ), .X(\us21\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0772_ ( .A(\us21\/_0162_ ), .X(\us21\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_0773_ ( .A(\us21\/_0293_ ), .B(\us21\/_0304_ ), .Y(\us21\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us21/_0774_ ( .A(\sa21\[1\] ), .Y(\us21\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us21/_0776_ ( .A(\sa21\[0\] ), .Y(\us21\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0777_ ( .A(\sa21\[2\] ), .B(\sa21\[3\] ), .X(\us21\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0779_ ( .A(\us21\/_0358_ ), .X(\us21\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_0780_ ( .A1(\us21\/_0325_ ), .A2(\us21\/_0347_ ), .B1(\us21\/_0380_ ), .C1(\us21\/_0304_ ), .Y(\us21\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us21/_0781_ ( .A_N(\us21\/_0238_ ), .B(\us21\/_0314_ ), .C(\us21\/_0391_ ), .X(\us21\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us21/_0782_ ( .A(\sa21\[3\] ), .B_N(\sa21\[2\] ), .Y(\us21\/_0412_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0784_ ( .A(\us21\/_0412_ ), .B(\us21\/_0205_ ), .X(\us21\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \us21/_0787_ ( .A(\sa21\[5\] ), .B_N(\sa21\[4\] ), .Y(\us21\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0788_ ( .A(\us21\/_0467_ ), .B(\us21\/_0140_ ), .X(\us21\/_0478_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_0791_ ( .A(\us21\/_0134_ ), .B(\us21\/_0218_ ), .Y(\us21\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_0792_ ( .A(\us21\/_0478_ ), .B(\us21\/_0271_ ), .Y(\us21\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0793_ ( .A(\us21\/_0194_ ), .X(\us21\/_0532_ ) );
sky130_fd_sc_hd__and2_1 \us21/_0795_ ( .A(\us21\/_0249_ ), .B(\us21\/_0358_ ), .X(\us21\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0797_ ( .A(\us21\/_0554_ ), .X(\us21\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us21/_0798_ ( .A(\us21\/_0205_ ), .B(\us21\/_0358_ ), .X(\us21\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0800_ ( .A(\us21\/_0586_ ), .X(\us21\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_0801_ ( .A1(\us21\/_0532_ ), .A2(\us21\/_0575_ ), .A3(\us21\/_0608_ ), .B1(\us21\/_0218_ ), .Y(\us21\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us21/_0802_ ( .A(\us21\/_0401_ ), .B(\us21\/_0510_ ), .C(\us21\/_0521_ ), .D(\us21\/_0619_ ), .X(\us21\/_0629_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0803_ ( .A(\us21\/_0358_ ), .B(\sa21\[1\] ), .X(\us21\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0805_ ( .A(\us21\/_0205_ ), .B(\us21\/_0260_ ), .X(\us21\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0807_ ( .A(\us21\/_0662_ ), .X(\us21\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us21/_0808_ ( .A(\sa21\[6\] ), .B_N(\sa21\[7\] ), .Y(\us21\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \us21/_0809_ ( .A(\us21\/_0467_ ), .B(\us21\/_0694_ ), .X(\us21\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0811_ ( .A(\us21\/_0705_ ), .X(\us21\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_0812_ ( .A1(\us21\/_0640_ ), .A2(\us21\/_0293_ ), .A3(\us21\/_0683_ ), .B1(\us21\/_0727_ ), .Y(\us21\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_0813_ ( .A(\sa21\[1\] ), .B(\sa21\[0\] ), .Y(\us21\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0814_ ( .A(\us21\/_0730_ ), .B(\us21\/_0260_ ), .X(\us21\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0816_ ( .A(\us21\/_0731_ ), .X(\us21\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0817_ ( .A(\sa21\[0\] ), .X(\us21\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us21/_0818_ ( .A1(\us21\/_0325_ ), .A2(\us21\/_0734_ ), .B1(\us21\/_0412_ ), .X(\us21\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0819_ ( .A(\us21\/_0694_ ), .B(\us21\/_0151_ ), .X(\us21\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0821_ ( .A(\us21\/_0736_ ), .X(\us21\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0822_ ( .A(\us21\/_0738_ ), .X(\us21\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_0823_ ( .A1(\us21\/_0733_ ), .A2(\us21\/_0735_ ), .A3(\us21\/_0293_ ), .B1(\us21\/_0739_ ), .Y(\us21\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us21/_0824_ ( .A(\us21\/_0730_ ), .B_N(\us21\/_0358_ ), .Y(\us21\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_0825_ ( .A(\us21\/_0741_ ), .B(\us21\/_0739_ ), .Y(\us21\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_0827_ ( .A1(\us21\/_0118_ ), .A2(\us21\/_0205_ ), .B1(\us21\/_0532_ ), .C1(\us21\/_0739_ ), .Y(\us21\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us21/_0828_ ( .A(\us21\/_0729_ ), .B(\us21\/_0740_ ), .C(\us21\/_0742_ ), .D(\us21\/_0744_ ), .X(\us21\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0829_ ( .A(\us21\/_0412_ ), .B(\us21\/_0730_ ), .X(\us21\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0830_ ( .A(\us21\/_0746_ ), .X(\us21\/_0747_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0831_ ( .A(\us21\/_0747_ ), .X(\us21\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us21/_0832_ ( .A(\sa21\[4\] ), .B_N(\sa21\[5\] ), .Y(\us21\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0833_ ( .A(\us21\/_0749_ ), .B(\us21\/_0694_ ), .X(\us21\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0835_ ( .A(\us21\/_0750_ ), .X(\us21\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0836_ ( .A(\us21\/_0752_ ), .X(\us21\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0837_ ( .A(\us21\/_0118_ ), .B(\us21\/_0358_ ), .X(\us21\/_0017_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0839_ ( .A(\us21\/_0752_ ), .B(\us21\/_0017_ ), .X(\us21\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0840_ ( .A(\us21\/_0358_ ), .B(\us21\/_0325_ ), .X(\us21\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0842_ ( .A(\us21\/_0096_ ), .B(\us21\/_0205_ ), .X(\us21\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \us21/_0844_ ( .A1(\us21\/_0020_ ), .A2(\us21\/_0022_ ), .B1(\us21\/_0752_ ), .X(\us21\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_0845_ ( .A1(\us21\/_0748_ ), .A2(\us21\/_0016_ ), .B1(\us21\/_0019_ ), .C1(\us21\/_0024_ ), .Y(\us21\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \us21/_0846_ ( .A(\sa21\[4\] ), .B(\sa21\[5\] ), .X(\us21\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0847_ ( .A(\us21\/_0694_ ), .B(\us21\/_0026_ ), .X(\us21\/_0027_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0850_ ( .A(\us21\/_0358_ ), .B(\us21\/_0730_ ), .X(\us21\/_0030_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0852_ ( .A(\us21\/_0030_ ), .X(\us21\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_0853_ ( .A(\us21\/_0247_ ), .B(\us21\/_0032_ ), .Y(\us21\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_0854_ ( .A(\us21\/_0247_ ), .B(\us21\/_0735_ ), .Y(\us21\/_0034_ ) );
sky130_fd_sc_hd__and2_1 \us21/_0855_ ( .A(\us21\/_0118_ ), .B(\us21\/_0260_ ), .X(\us21\/_0035_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0857_ ( .A(\us21\/_0027_ ), .B(\us21\/_0035_ ), .X(\us21\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0858_ ( .A(\us21\/_0260_ ), .X(\us21\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_0859_ ( .A(\us21\/_0038_ ), .B(\us21\/_0347_ ), .Y(\us21\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us21/_0860_ ( .A_N(\us21\/_0039_ ), .B(\us21\/_0027_ ), .X(\us21\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_0861_ ( .A(\us21\/_0037_ ), .B(\us21\/_0040_ ), .Y(\us21\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us21/_0862_ ( .A(\us21\/_0025_ ), .B(\us21\/_0033_ ), .C(\us21\/_0034_ ), .D(\us21\/_0041_ ), .X(\us21\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0863_ ( .A(\us21\/_0749_ ), .B(\us21\/_0140_ ), .X(\us21\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us21/_0865_ ( .A(\sa21\[0\] ), .B(\sa21\[2\] ), .C(\sa21\[3\] ), .X(\us21\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0866_ ( .A(\us21\/_0043_ ), .B(\us21\/_0045_ ), .X(\us21\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0867_ ( .A(\us21\/_0096_ ), .B(\us21\/_0249_ ), .X(\us21\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0869_ ( .A(\us21\/_0047_ ), .B(\us21\/_0043_ ), .X(\us21\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0870_ ( .A(\us21\/_0730_ ), .X(\us21\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0871_ ( .A(\us21\/_0043_ ), .X(\us21\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_0872_ ( .A1(\us21\/_0118_ ), .A2(\us21\/_0050_ ), .B1(\us21\/_0194_ ), .C1(\us21\/_0051_ ), .Y(\us21\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us21/_0873_ ( .A(\us21\/_0046_ ), .B(\us21\/_0049_ ), .C_N(\us21\/_0052_ ), .Y(\us21\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0874_ ( .A(\us21\/_0026_ ), .B(\us21\/_0140_ ), .X(\us21\/_0054_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0876_ ( .A(\us21\/_0054_ ), .X(\us21\/_0056_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_0877_ ( .A1(\us21\/_0532_ ), .A2(\us21\/_0575_ ), .B1(\us21\/_0056_ ), .Y(\us21\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0878_ ( .A(\us21\/_0412_ ), .B(\us21\/_0325_ ), .X(\us21\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0880_ ( .A(\us21\/_0051_ ), .X(\us21\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_0881_ ( .A1(\us21\/_0731_ ), .A2(\us21\/_0035_ ), .A3(\us21\/_0058_ ), .B1(\us21\/_0060_ ), .Y(\us21\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0882_ ( .A(\us21\/_0260_ ), .B(\sa21\[1\] ), .X(\us21\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0884_ ( .A(\us21\/_0062_ ), .X(\us21\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_0885_ ( .A1(\us21\/_0064_ ), .A2(\us21\/_0748_ ), .A3(\us21\/_0683_ ), .B1(\us21\/_0056_ ), .Y(\us21\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us21/_0886_ ( .A(\us21\/_0053_ ), .B(\us21\/_0057_ ), .C(\us21\/_0061_ ), .D(\us21\/_0065_ ), .X(\us21\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us21/_0887_ ( .A(\us21\/_0629_ ), .B(\us21\/_0745_ ), .C(\us21\/_0042_ ), .D(\us21\/_0066_ ), .X(\us21\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us21/_0889_ ( .A(\sa21\[7\] ), .B_N(\sa21\[6\] ), .Y(\us21\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0890_ ( .A(\us21\/_0069_ ), .B(\us21\/_0151_ ), .X(\us21\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0892_ ( .A(\us21\/_0070_ ), .X(\us21\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_0893_ ( .A1(\us21\/_0129_ ), .A2(\us21\/_0586_ ), .B1(\us21\/_0072_ ), .Y(\us21\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_0894_ ( .A1(\us21\/_0380_ ), .A2(\us21\/_0347_ ), .B1(\us21\/_0194_ ), .B2(\us21\/_0205_ ), .Y(\us21\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us21/_0895_ ( .A(\us21\/_0074_ ), .B_N(\us21\/_0070_ ), .Y(\us21\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us21/_0896_ ( .A(\us21\/_0073_ ), .SLEEP(\us21\/_0075_ ), .X(\us21\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us21/_0897_ ( .A(\us21\/_0467_ ), .B(\us21\/_0069_ ), .X(\us21\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0898_ ( .A(\us21\/_0077_ ), .X(\us21\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0899_ ( .A(\us21\/_0412_ ), .B(\us21\/_0118_ ), .X(\us21\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0901_ ( .A(\us21\/_0078_ ), .B(\us21\/_0079_ ), .X(\us21\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0902_ ( .A(\us21\/_0412_ ), .B(\us21\/_0249_ ), .X(\us21\/_0082_ ) );
sky130_fd_sc_hd__buf_2 \us21/_0904_ ( .A(\us21\/_0082_ ), .X(\us21\/_0084_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0905_ ( .A(\us21\/_0084_ ), .B(\us21\/_0078_ ), .X(\us21\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us21/_0906_ ( .A1(\sa21\[0\] ), .A2(\us21\/_0325_ ), .B1(\us21\/_0260_ ), .Y(\us21\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us21/_0907_ ( .A_N(\us21\/_0086_ ), .B(\us21\/_0078_ ), .X(\us21\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us21/_0908_ ( .A(\us21\/_0081_ ), .B(\us21\/_0085_ ), .C(\us21\/_0087_ ), .Y(\us21\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0909_ ( .A(\us21\/_0072_ ), .X(\us21\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_0910_ ( .A1(\us21\/_0733_ ), .A2(\us21\/_0748_ ), .A3(\us21\/_0683_ ), .B1(\us21\/_0089_ ), .Y(\us21\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0911_ ( .A(\us21\/_0129_ ), .X(\us21\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0912_ ( .A(\us21\/_0017_ ), .X(\us21\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0913_ ( .A(\us21\/_0022_ ), .X(\us21\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0914_ ( .A(\us21\/_0078_ ), .X(\us21\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_0915_ ( .A1(\us21\/_0091_ ), .A2(\us21\/_0092_ ), .A3(\us21\/_0093_ ), .B1(\us21\/_0094_ ), .Y(\us21\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us21/_0916_ ( .A(\us21\/_0076_ ), .B(\us21\/_0088_ ), .C(\us21\/_0090_ ), .D(\us21\/_0095_ ), .X(\us21\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us21/_0917_ ( .A(\us21\/_0069_ ), .B(\us21\/_0026_ ), .X(\us21\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \us21/_0918_ ( .A(\us21\/_0098_ ), .X(\us21\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0919_ ( .A(\us21\/_0434_ ), .B(\us21\/_0099_ ), .X(\us21\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0920_ ( .A(\us21\/_0079_ ), .B(\us21\/_0098_ ), .X(\us21\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0921_ ( .A(\us21\/_0325_ ), .X(\us21\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_0922_ ( .A1(\us21\/_0102_ ), .A2(\us21\/_0734_ ), .B1(\us21\/_0038_ ), .C1(\us21\/_0099_ ), .Y(\us21\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us21/_0923_ ( .A(\us21\/_0100_ ), .B(\us21\/_0101_ ), .C_N(\us21\/_0103_ ), .Y(\us21\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_0924_ ( .A1(\us21\/_0554_ ), .A2(\us21\/_0586_ ), .B1(\us21\/_0099_ ), .Y(\us21\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_0925_ ( .A(\us21\/_0129_ ), .B(\us21\/_0099_ ), .Y(\us21\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0926_ ( .A(\us21\/_0105_ ), .B(\us21\/_0106_ ), .X(\us21\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0927_ ( .A(\us21\/_0412_ ), .X(\us21\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us21/_0928_ ( .A(\us21\/_0260_ ), .B(\sa21\[0\] ), .X(\us21\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0929_ ( .A(\us21\/_0069_ ), .B(\us21\/_0749_ ), .X(\us21\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0931_ ( .A(\us21\/_0111_ ), .X(\us21\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0932_ ( .A(\us21\/_0113_ ), .X(\us21\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_0933_ ( .A1(\us21\/_0109_ ), .A2(\us21\/_0110_ ), .B1(\us21\/_0114_ ), .Y(\us21\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us21/_0934_ ( .A(\us21\/_0022_ ), .Y(\us21\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us21/_0935_ ( .A(\us21\/_0554_ ), .Y(\us21\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us21/_0936_ ( .A1(\us21\/_0050_ ), .A2(\us21\/_0118_ ), .B1(\us21\/_0194_ ), .Y(\us21\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us21/_0937_ ( .A(\us21\/_0113_ ), .Y(\us21\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us21/_0938_ ( .A1(\us21\/_0116_ ), .A2(\us21\/_0117_ ), .A3(\us21\/_0119_ ), .B1(\us21\/_0120_ ), .X(\us21\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us21/_0939_ ( .A(\us21\/_0104_ ), .B(\us21\/_0108_ ), .C(\us21\/_0115_ ), .D(\us21\/_0121_ ), .X(\us21\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_0940_ ( .A(\sa21\[7\] ), .B(\sa21\[6\] ), .Y(\us21\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0941_ ( .A(\us21\/_0749_ ), .B(\us21\/_0123_ ), .X(\us21\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0943_ ( .A(\us21\/_0082_ ), .B(\us21\/_0124_ ), .X(\us21\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_0944_ ( .A(\us21\/_0271_ ), .B(\us21\/_0124_ ), .Y(\us21\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0945_ ( .A(\us21\/_0124_ ), .X(\us21\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0946_ ( .A(\us21\/_0260_ ), .B(\us21\/_0325_ ), .X(\us21\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_0948_ ( .A(\us21\/_0128_ ), .B(\us21\/_0130_ ), .Y(\us21\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_0949_ ( .A(\us21\/_0127_ ), .B(\us21\/_0132_ ), .Y(\us21\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us21/_0950_ ( .A(\us21\/_0434_ ), .X(\us21\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_0951_ ( .A(\us21\/_0134_ ), .B(\us21\/_0128_ ), .Y(\us21\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us21/_0952_ ( .A(\us21\/_0126_ ), .B(\us21\/_0133_ ), .C_N(\us21\/_0135_ ), .Y(\us21\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us21/_0953_ ( .A(\us21\/_0026_ ), .B(\us21\/_0123_ ), .X(\us21\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0955_ ( .A(\us21\/_0137_ ), .X(\us21\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_0956_ ( .A1(\us21\/_0110_ ), .A2(\us21\/_0293_ ), .A3(\us21\/_0084_ ), .B1(\us21\/_0139_ ), .Y(\us21\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0957_ ( .A(\us21\/_0096_ ), .B(\us21\/_0730_ ), .X(\us21\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0959_ ( .A(\us21\/_0142_ ), .X(\us21\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_0960_ ( .A1(\us21\/_0020_ ), .A2(\us21\/_0144_ ), .A3(\us21\/_0017_ ), .B1(\us21\/_0139_ ), .Y(\us21\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \us21/_0961_ ( .A(\sa21\[2\] ), .B(\us21\/_0050_ ), .C_N(\sa21\[3\] ), .Y(\us21\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0962_ ( .A(\us21\/_0128_ ), .X(\us21\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_0963_ ( .A1(\us21\/_0146_ ), .A2(\us21\/_0032_ ), .A3(\us21\/_0640_ ), .B1(\us21\/_0147_ ), .Y(\us21\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us21/_0964_ ( .A(\us21\/_0136_ ), .B(\us21\/_0141_ ), .C(\us21\/_0145_ ), .D(\us21\/_0148_ ), .X(\us21\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0965_ ( .A(\us21\/_0123_ ), .B(\us21\/_0151_ ), .X(\us21\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0967_ ( .A(\us21\/_0150_ ), .X(\us21\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \us21/_0968_ ( .A(\us21\/_0150_ ), .B(\us21\/_0062_ ), .X(\us21\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_0969_ ( .A(\us21\/_0079_ ), .B(\us21\/_0150_ ), .Y(\us21\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us21/_0970_ ( .A(\us21\/_0150_ ), .B(\us21\/_0412_ ), .C(\us21\/_0249_ ), .Y(\us21\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_0971_ ( .A(\us21\/_0155_ ), .B(\us21\/_0156_ ), .Y(\us21\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_0972_ ( .A1(\us21\/_0153_ ), .A2(\us21\/_0134_ ), .B1(\us21\/_0154_ ), .C1(\us21\/_0157_ ), .Y(\us21\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0973_ ( .A(\us21\/_0467_ ), .B(\us21\/_0123_ ), .X(\us21\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_0975_ ( .A(\us21\/_0159_ ), .X(\us21\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us21/_0976_ ( .A_N(\us21\/_0119_ ), .B(\us21\/_0161_ ), .X(\us21\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us21/_0977_ ( .A(\us21\/_0163_ ), .Y(\us21\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_0978_ ( .A1(\us21\/_0146_ ), .A2(\us21\/_0575_ ), .A3(\us21\/_0608_ ), .B1(\us21\/_0153_ ), .Y(\us21\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_0979_ ( .A1(\us21\/_0062_ ), .A2(\us21\/_0084_ ), .A3(\us21\/_0134_ ), .B1(\us21\/_0161_ ), .Y(\us21\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us21/_0980_ ( .A(\us21\/_0158_ ), .B(\us21\/_0164_ ), .C(\us21\/_0165_ ), .D(\us21\/_0166_ ), .X(\us21\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us21/_0981_ ( .A(\us21\/_0097_ ), .B(\us21\/_0122_ ), .C(\us21\/_0149_ ), .D(\us21\/_0167_ ), .X(\us21\/_0168_ ) );
sky130_fd_sc_hd__and2_1 \us21/_0982_ ( .A(\us21\/_0662_ ), .B(\us21\/_0150_ ), .X(\us21\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_0983_ ( .A(\us21\/_0154_ ), .B(\us21\/_0169_ ), .Y(\us21\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us21/_0984_ ( .A(\us21\/_0123_ ), .B(\us21\/_0151_ ), .C(\us21\/_0038_ ), .X(\us21\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0985_ ( .A(\us21\/_0170_ ), .B(\us21\/_0171_ ), .X(\us21\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \us21/_0986_ ( .A(\us21\/_0172_ ), .Y(\us21\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \us21/_0987_ ( .A(\us21\/_0067_ ), .B(\us21\/_0168_ ), .C(\us21\/_0174_ ), .Y(\us21\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us21/_0988_ ( .A(\sa21\[1\] ), .B(\sa21\[0\] ), .Y(\us21\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us21/_0989_ ( .A(\us21\/_0175_ ), .B(\us21\/_0358_ ), .X(\us21\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0990_ ( .A(\us21\/_0176_ ), .B(\us21\/_0478_ ), .X(\us21\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_0991_ ( .A(\us21\/_0084_ ), .B(\us21\/_0113_ ), .Y(\us21\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0992_ ( .A(\us21\/_0111_ ), .B(\us21\/_0062_ ), .X(\us21\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0993_ ( .A(\us21\/_0111_ ), .B(\us21\/_0662_ ), .X(\us21\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_0994_ ( .A(\us21\/_0179_ ), .B(\us21\/_0180_ ), .Y(\us21\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0995_ ( .A(\us21\/_0054_ ), .B(\us21\/_0058_ ), .X(\us21\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us21/_0996_ ( .A(\us21\/_0182_ ), .Y(\us21\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us21/_0997_ ( .A_N(\us21\/_0177_ ), .B(\us21\/_0178_ ), .C(\us21\/_0181_ ), .D(\us21\/_0184_ ), .X(\us21\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0998_ ( .A(\us21\/_0098_ ), .B(\us21\/_0741_ ), .X(\us21\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us21/_0999_ ( .A(\us21\/_0047_ ), .B(\us21\/_0098_ ), .X(\us21\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us21/_1000_ ( .A(\us21\/_0186_ ), .B(\us21\/_0187_ ), .X(\us21\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1001_ ( .A(\us21\/_0188_ ), .Y(\us21\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1002_ ( .A(\us21\/_0738_ ), .B(\us21\/_0735_ ), .X(\us21\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1003_ ( .A(\us21\/_0271_ ), .B(\us21\/_0736_ ), .X(\us21\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_1004_ ( .A(\us21\/_0190_ ), .B(\us21\/_0191_ ), .Y(\us21\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us21/_1005_ ( .A(\us21\/_0096_ ), .B(\us21\/_0325_ ), .X(\us21\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1006_ ( .A1(\us21\/_0193_ ), .A2(\us21\/_0176_ ), .B1(\us21\/_0043_ ), .Y(\us21\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1007_ ( .A(\us21\/_0185_ ), .B(\us21\/_0189_ ), .C(\us21\/_0192_ ), .D(\us21\/_0195_ ), .X(\us21\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us21/_1008_ ( .A_N(\sa21\[3\] ), .B(\us21\/_0734_ ), .C(\sa21\[2\] ), .X(\us21\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1009_ ( .A(\us21\/_0137_ ), .B(\us21\/_0197_ ), .X(\us21\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_1010_ ( .A(\us21\/_0198_ ), .B(\us21\/_0040_ ), .Y(\us21\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1011_ ( .A(\us21\/_0293_ ), .B(\us21\/_0137_ ), .X(\us21\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1012_ ( .A(\us21\/_0200_ ), .Y(\us21\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1013_ ( .A(\us21\/_0137_ ), .B(\us21\/_0110_ ), .Y(\us21\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1014_ ( .A(\us21\/_0139_ ), .B(\us21\/_0020_ ), .Y(\us21\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1015_ ( .A(\us21\/_0199_ ), .B(\us21\/_0201_ ), .C(\us21\/_0202_ ), .D(\us21\/_0203_ ), .X(\us21\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us21/_1016_ ( .A1(\us21\/_0532_ ), .A2(\us21\/_0109_ ), .B1(\us21\/_0102_ ), .C1(\us21\/_0727_ ), .X(\us21\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1017_ ( .A(\us21\/_0022_ ), .B(\us21\/_0078_ ), .Y(\us21\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1018_ ( .A(\us21\/_0078_ ), .B(\us21\/_0142_ ), .Y(\us21\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1019_ ( .A(\us21\/_0207_ ), .B(\us21\/_0208_ ), .Y(\us21\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1020_ ( .A1(\us21\/_0094_ ), .A2(\us21\/_0176_ ), .B1(\us21\/_0206_ ), .C1(\us21\/_0209_ ), .Y(\us21\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1021_ ( .A(\us21\/_0662_ ), .B(\us21\/_0070_ ), .X(\us21\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us21/_1022_ ( .A(\us21\/_0731_ ), .B(\us21\/_0123_ ), .C(\us21\/_0749_ ), .Y(\us21\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us21/_1023_ ( .A(\us21\/_0731_ ), .B(\us21\/_0467_ ), .C(\us21\/_0069_ ), .Y(\us21\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us21/_1024_ ( .A_N(\us21\/_0211_ ), .B(\us21\/_0127_ ), .C(\us21\/_0212_ ), .D(\us21\/_0213_ ), .X(\us21\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1025_ ( .A(\us21\/_0137_ ), .Y(\us21\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1026_ ( .A(\us21\/_0128_ ), .B(\us21\/_0035_ ), .Y(\us21\/_0217_ ) );
sky130_fd_sc_hd__buf_2 \us21/_1027_ ( .A(\us21\/_0478_ ), .X(\us21\/_0218_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1028_ ( .A1(\us21\/_0159_ ), .A2(\us21\/_0747_ ), .B1(\us21\/_0434_ ), .B2(\us21\/_0218_ ), .Y(\us21\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us21/_1029_ ( .A1(\us21\/_0116_ ), .A2(\us21\/_0215_ ), .B1(\us21\/_0217_ ), .C1(\us21\/_0219_ ), .X(\us21\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1030_ ( .A(\us21\/_0113_ ), .B(\us21\/_0746_ ), .X(\us21\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us21/_1031_ ( .A1(\us21\/_0098_ ), .A2(\us21\/_0746_ ), .B1(\us21\/_0434_ ), .B2(\us21\/_0750_ ), .X(\us21\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1032_ ( .A1(\us21\/_0047_ ), .A2(\us21\/_0113_ ), .B1(\us21\/_0221_ ), .C1(\us21\/_0222_ ), .Y(\us21\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us21/_1033_ ( .A1(\us21\/_0129_ ), .A2(\us21\/_0162_ ), .B1(\us21\/_0271_ ), .B2(\us21\/_0705_ ), .X(\us21\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1034_ ( .A1(\us21\/_0093_ ), .A2(\us21\/_0738_ ), .B1(\us21\/_0081_ ), .C1(\us21\/_0224_ ), .Y(\us21\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1035_ ( .A(\us21\/_0214_ ), .B(\us21\/_0220_ ), .C(\us21\/_0223_ ), .D(\us21\/_0225_ ), .X(\us21\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1036_ ( .A(\us21\/_0196_ ), .B(\us21\/_0204_ ), .C(\us21\/_0210_ ), .D(\us21\/_0226_ ), .X(\us21\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1037_ ( .A(\us21\/_0111_ ), .B(\us21\/_0554_ ), .X(\us21\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1038_ ( .A(\us21\/_0229_ ), .Y(\us21\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1039_ ( .A(\us21\/_0111_ ), .B(\us21\/_0129_ ), .Y(\us21\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1040_ ( .A(\us21\/_0017_ ), .B(\us21\/_0738_ ), .Y(\us21\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1041_ ( .A(\us21\/_0030_ ), .B(\us21\/_0304_ ), .Y(\us21\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1042_ ( .A(\us21\/_0230_ ), .B(\us21\/_0231_ ), .C(\us21\/_0232_ ), .D(\us21\/_0233_ ), .X(\us21\/_0234_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1043_ ( .A(\us21\/_0047_ ), .B(\us21\/_0478_ ), .X(\us21\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1044_ ( .A1(\us21\/_0129_ ), .A2(\us21\/_0554_ ), .B1(\us21\/_0137_ ), .Y(\us21\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us21/_1045_ ( .A(\us21\/_0235_ ), .B(\us21\/_0049_ ), .C_N(\us21\/_0236_ ), .Y(\us21\/_0237_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1046_ ( .A(\us21\/_0047_ ), .B(\us21\/_0077_ ), .X(\us21\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1047_ ( .A(\us21\/_0070_ ), .B(\us21\/_0035_ ), .X(\us21\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us21/_1048_ ( .A1(\us21\/_0047_ ), .A2(\us21\/_0736_ ), .B1(\us21\/_0022_ ), .B2(\us21\/_0099_ ), .X(\us21\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us21/_1049_ ( .A(\us21\/_0239_ ), .B(\us21\/_0240_ ), .C(\us21\/_0241_ ), .Y(\us21\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1050_ ( .A(\us21\/_0554_ ), .B(\us21\/_0072_ ), .X(\us21\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us21/_1051_ ( .A1(\us21\/_0142_ ), .A2(\us21\/_0137_ ), .B1(\us21\/_0159_ ), .B2(\us21\/_0082_ ), .X(\us21\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1052_ ( .A1(\us21\/_0608_ ), .A2(\us21\/_0072_ ), .B1(\us21\/_0243_ ), .C1(\us21\/_0244_ ), .Y(\us21\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1053_ ( .A(\us21\/_0234_ ), .B(\us21\/_0237_ ), .C(\us21\/_0242_ ), .D(\us21\/_0245_ ), .X(\us21\/_0246_ ) );
sky130_fd_sc_hd__buf_2 \us21/_1054_ ( .A(\us21\/_0027_ ), .X(\us21\/_0247_ ) );
sky130_fd_sc_hd__o21a_1 \us21/_1055_ ( .A1(\us21\/_0554_ ), .A2(\us21\/_0586_ ), .B1(\us21\/_0247_ ), .X(\us21\/_0248_ ) );
sky130_fd_sc_hd__and2_1 \us21/_1056_ ( .A(\us21\/_0082_ ), .B(\us21\/_0478_ ), .X(\us21\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_1057_ ( .A(\us21\/_0079_ ), .X(\us21\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1058_ ( .A(\us21\/_0251_ ), .B(\us21\/_0478_ ), .X(\us21\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_1059_ ( .A(\us21\/_0250_ ), .B(\us21\/_0252_ ), .Y(\us21\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1060_ ( .A(\us21\/_0016_ ), .B(\us21\/_0064_ ), .Y(\us21\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_1061_ ( .A(\us21\/_0304_ ), .X(\us21\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1062_ ( .A(\us21\/_0255_ ), .B(\us21\/_0640_ ), .Y(\us21\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us21/_1063_ ( .A_N(\us21\/_0248_ ), .B(\us21\/_0253_ ), .C(\us21\/_0254_ ), .D(\us21\/_0256_ ), .X(\us21\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1064_ ( .A(\us21\/_0099_ ), .B(\us21\/_0110_ ), .X(\us21\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us21/_1065_ ( .A1(\us21\/_0161_ ), .A2(\us21\/_0130_ ), .B1(\us21\/_0258_ ), .Y(\us21\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1066_ ( .A(\us21\/_0194_ ), .B(\sa21\[1\] ), .X(\us21\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1068_ ( .A(\us21\/_0261_ ), .B(\us21\/_0153_ ), .Y(\us21\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us21/_1069_ ( .A_N(\us21\/_0154_ ), .B(\us21\/_0259_ ), .C(\us21\/_0263_ ), .X(\us21\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1070_ ( .A(\us21\/_0246_ ), .B(\us21\/_0174_ ), .C(\us21\/_0257_ ), .D(\us21\/_0264_ ), .X(\us21\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us21/_1071_ ( .A1(\us21\/_0261_ ), .A2(\us21\/_0554_ ), .B1(\us21\/_0159_ ), .X(\us21\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1072_ ( .A(\us21\/_0747_ ), .B(\us21\/_0150_ ), .Y(\us21\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1073_ ( .A(\us21\/_0175_ ), .Y(\us21\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us21/_1074_ ( .A(\us21\/_0412_ ), .B(\us21\/_0123_ ), .C(\us21\/_0151_ ), .X(\us21\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1075_ ( .A(\us21\/_0268_ ), .B(\us21\/_0269_ ), .Y(\us21\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us21/_1076_ ( .A_N(\us21\/_0266_ ), .B(\us21\/_0267_ ), .C(\us21\/_0270_ ), .X(\us21\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1077_ ( .A(\us21\/_0554_ ), .B(\us21\/_0150_ ), .X(\us21\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1078_ ( .A(\us21\/_0273_ ), .Y(\us21\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1079_ ( .A1(\us21\/_0734_ ), .A2(\us21\/_0325_ ), .B1(\us21\/_0380_ ), .Y(\us21\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1080_ ( .A(\us21\/_0275_ ), .Y(\us21\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1081_ ( .A(\us21\/_0276_ ), .B(\us21\/_0153_ ), .Y(\us21\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us21/_1082_ ( .A(\us21\/_0272_ ), .B(\us21\/_0274_ ), .C(\us21\/_0277_ ), .X(\us21\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_1083_ ( .A(\us21\/_0035_ ), .X(\us21\/_0279_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1085_ ( .A1(\us21\/_0218_ ), .A2(\us21\/_0279_ ), .B1(\us21\/_0084_ ), .B2(\us21\/_0060_ ), .Y(\us21\/_0281_ ) );
sky130_fd_sc_hd__o21ai_1 \us21/_1086_ ( .A1(\us21\/_0251_ ), .A2(\us21\/_0434_ ), .B1(\us21\/_0304_ ), .Y(\us21\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1087_ ( .A(\us21\/_0091_ ), .B(\us21\/_0056_ ), .Y(\us21\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1088_ ( .A1(\us21\/_0118_ ), .A2(\us21\/_0050_ ), .B1(\us21\/_0038_ ), .C1(\us21\/_0255_ ), .Y(\us21\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1089_ ( .A(\us21\/_0281_ ), .B(\us21\/_0283_ ), .C(\us21\/_0284_ ), .D(\us21\/_0285_ ), .X(\us21\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1090_ ( .A(\us21\/_0082_ ), .B(\us21\/_0027_ ), .X(\us21\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1091_ ( .A(\us21\/_0129_ ), .B(\us21\/_0027_ ), .X(\us21\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_1092_ ( .A(\us21\/_0287_ ), .B(\us21\/_0288_ ), .Y(\us21\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1093_ ( .A1(\us21\/_0752_ ), .A2(\us21\/_0683_ ), .B1(\us21\/_0093_ ), .B2(\us21\/_0247_ ), .Y(\us21\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1094_ ( .A1(\us21\/_0092_ ), .A2(\us21\/_0575_ ), .B1(\us21\/_0056_ ), .Y(\us21\/_0291_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1096_ ( .A1(\us21\/_0218_ ), .A2(\us21\/_0662_ ), .B1(\us21\/_0084_ ), .B2(\us21\/_0056_ ), .Y(\us21\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1097_ ( .A(\us21\/_0289_ ), .B(\us21\/_0290_ ), .C(\us21\/_0291_ ), .D(\us21\/_0294_ ), .X(\us21\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1098_ ( .A(\us21\/_0750_ ), .B(\us21\/_0193_ ), .X(\us21\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1099_ ( .A(\us21\/_0705_ ), .B(\us21\/_0380_ ), .X(\us21\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1100_ ( .A(\us21\/_0752_ ), .B(\us21\/_0129_ ), .Y(\us21\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us21/_1101_ ( .A(\us21\/_0296_ ), .B(\us21\/_0297_ ), .C_N(\us21\/_0298_ ), .Y(\us21\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1102_ ( .A(\us21\/_0089_ ), .B(\us21\/_0532_ ), .Y(\us21\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1103_ ( .A(\sa21\[2\] ), .Y(\us21\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \us21/_1104_ ( .A(\us21\/_0301_ ), .B(\sa21\[3\] ), .C(\us21\/_0118_ ), .Y(\us21\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1105_ ( .A(\us21\/_0072_ ), .B(\us21\/_0302_ ), .X(\us21\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1106_ ( .A(\us21\/_0303_ ), .Y(\us21\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1107_ ( .A(\us21\/_0147_ ), .B(\us21\/_0302_ ), .Y(\us21\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1108_ ( .A(\us21\/_0299_ ), .B(\us21\/_0300_ ), .C(\us21\/_0305_ ), .D(\us21\/_0306_ ), .X(\us21\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1109_ ( .A(\us21\/_0278_ ), .B(\us21\/_0286_ ), .C(\us21\/_0295_ ), .D(\us21\/_0307_ ), .X(\us21\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us21/_1110_ ( .A(\us21\/_0228_ ), .B(\us21\/_0265_ ), .C(\us21\/_0308_ ), .Y(\us21\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1111_ ( .A(\us21\/_0235_ ), .Y(\us21\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1112_ ( .A(\us21\/_0478_ ), .B(\us21\/_0640_ ), .X(\us21\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1113_ ( .A(\us21\/_0310_ ), .Y(\us21\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1114_ ( .A(\us21\/_0022_ ), .B(\us21\/_0218_ ), .Y(\us21\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1115_ ( .A(\us21\/_0218_ ), .B(\us21\/_0032_ ), .Y(\us21\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1116_ ( .A(\us21\/_0309_ ), .B(\us21\/_0311_ ), .C(\us21\/_0312_ ), .D(\us21\/_0313_ ), .X(\us21\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1117_ ( .A(\us21\/_0218_ ), .B(\us21\/_0064_ ), .Y(\us21\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1118_ ( .A(\us21\/_0218_ ), .B(\us21\/_0683_ ), .Y(\us21\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1119_ ( .A(\us21\/_0315_ ), .B(\us21\/_0316_ ), .C(\us21\/_0317_ ), .D(\us21\/_0253_ ), .X(\us21\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1120_ ( .A(\us21\/_0047_ ), .B(\us21\/_0304_ ), .Y(\us21\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1121_ ( .A(\us21\/_0586_ ), .B(\us21\/_0162_ ), .Y(\us21\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1122_ ( .A(\us21\/_0319_ ), .B(\us21\/_0320_ ), .Y(\us21\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_1123_ ( .A(\us21\/_0321_ ), .B(\us21\/_0238_ ), .Y(\us21\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1124_ ( .A(\us21\/_0304_ ), .B(\us21\/_0062_ ), .Y(\us21\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_1125_ ( .A(\us21\/_0251_ ), .X(\us21\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1126_ ( .A1(\us21\/_0324_ ), .A2(\us21\/_0084_ ), .B1(\us21\/_0255_ ), .Y(\us21\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1127_ ( .A1(\us21\/_0050_ ), .A2(\us21\/_0205_ ), .B1(\us21\/_0109_ ), .C1(\us21\/_0255_ ), .Y(\us21\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1128_ ( .A(\us21\/_0322_ ), .B(\us21\/_0323_ ), .C(\us21\/_0326_ ), .D(\us21\/_0327_ ), .X(\us21\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1129_ ( .A1(\us21\/_0733_ ), .A2(\us21\/_0279_ ), .A3(\us21\/_0058_ ), .B1(\us21\/_0056_ ), .Y(\us21\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_1130_ ( .A(\us21\/_0047_ ), .X(\us21\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1131_ ( .A(\us21\/_0330_ ), .B(\us21\/_0056_ ), .Y(\us21\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1132_ ( .A(\us21\/_0054_ ), .B(\us21\/_0045_ ), .Y(\us21\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1133_ ( .A(\us21\/_0329_ ), .B(\us21\/_0331_ ), .C(\us21\/_0284_ ), .D(\us21\/_0332_ ), .X(\us21\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us21/_1134_ ( .A1(\us21\/_0249_ ), .A2(\us21\/_0205_ ), .B1(\us21\/_0532_ ), .C1(\us21\/_0060_ ), .X(\us21\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1135_ ( .A(\us21\/_0084_ ), .B(\us21\/_0060_ ), .Y(\us21\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1136_ ( .A(\us21\/_0324_ ), .B(\us21\/_0060_ ), .Y(\us21\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1137_ ( .A(\us21\/_0335_ ), .B(\us21\/_0337_ ), .Y(\us21\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1138_ ( .A1(\us21\/_0276_ ), .A2(\us21\/_0060_ ), .B1(\us21\/_0334_ ), .C1(\us21\/_0338_ ), .Y(\us21\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1139_ ( .A(\us21\/_0318_ ), .B(\us21\/_0328_ ), .C(\us21\/_0333_ ), .D(\us21\/_0339_ ), .X(\us21\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us21/_1140_ ( .A1(\us21\/_0747_ ), .A2(\us21\/_0134_ ), .B1(\us21\/_0128_ ), .X(\us21\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us21/_1141_ ( .A_N(\us21\/_0086_ ), .B(\us21\/_0128_ ), .X(\us21\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1142_ ( .A(\us21\/_0079_ ), .B(\us21\/_0124_ ), .X(\us21\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_1143_ ( .A(\us21\/_0126_ ), .B(\us21\/_0343_ ), .Y(\us21\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us21/_1144_ ( .A(\us21\/_0341_ ), .B(\us21\/_0342_ ), .C_N(\us21\/_0344_ ), .Y(\us21\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1146_ ( .A1(\us21\/_0193_ ), .A2(\us21\/_0092_ ), .A3(\us21\/_0330_ ), .B1(\us21\/_0147_ ), .Y(\us21\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1147_ ( .A1(\us21\/_0130_ ), .A2(\us21\/_0084_ ), .A3(\us21\/_0134_ ), .B1(\us21\/_0139_ ), .Y(\us21\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1148_ ( .A1(\us21\/_0144_ ), .A2(\us21\/_0608_ ), .A3(\us21\/_0092_ ), .B1(\us21\/_0139_ ), .Y(\us21\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1149_ ( .A(\us21\/_0345_ ), .B(\us21\/_0348_ ), .C(\us21\/_0349_ ), .D(\us21\/_0350_ ), .X(\us21\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us21/_1150_ ( .A(\us21\/_0150_ ), .B(\us21\/_0194_ ), .C(\us21\/_0249_ ), .X(\us21\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us21/_1151_ ( .A(\us21\/_0277_ ), .SLEEP(\us21\/_0352_ ), .X(\us21\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us21/_1152_ ( .A1(\us21\/_0268_ ), .A2(\us21\/_0171_ ), .B1(\us21\/_0157_ ), .Y(\us21\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us21/_1153_ ( .A(\us21\/_0161_ ), .X(\us21\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1154_ ( .A1(\us21\/_0279_ ), .A2(\us21\/_0084_ ), .B1(\us21\/_0355_ ), .Y(\us21\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1155_ ( .A1(\us21\/_0020_ ), .A2(\us21\/_0193_ ), .A3(\us21\/_0091_ ), .B1(\us21\/_0355_ ), .Y(\us21\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1156_ ( .A(\us21\/_0353_ ), .B(\us21\/_0354_ ), .C(\us21\/_0356_ ), .D(\us21\/_0357_ ), .X(\us21\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1157_ ( .A(\us21\/_0111_ ), .B(\us21\/_0586_ ), .X(\us21\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1158_ ( .A(\us21\/_0360_ ), .Y(\us21\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us21/_1159_ ( .A1(\us21\/_0119_ ), .A2(\us21\/_0120_ ), .B1(\us21\/_0230_ ), .C1(\us21\/_0361_ ), .X(\us21\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1160_ ( .A1(\us21\/_0662_ ), .A2(\us21\/_0251_ ), .A3(\us21\/_0134_ ), .B1(\us21\/_0114_ ), .Y(\us21\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1162_ ( .A1(\us21\/_0035_ ), .A2(\us21\/_0251_ ), .A3(\us21\/_0134_ ), .B1(\us21\/_0099_ ), .Y(\us21\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1163_ ( .A1(\us21\/_0193_ ), .A2(\us21\/_0608_ ), .B1(\us21\/_0099_ ), .Y(\us21\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1164_ ( .A(\us21\/_0362_ ), .B(\us21\/_0363_ ), .C(\us21\/_0365_ ), .D(\us21\/_0366_ ), .X(\us21\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1165_ ( .A1(\us21\/_0575_ ), .A2(\us21\/_0092_ ), .A3(\us21\/_0330_ ), .B1(\us21\/_0089_ ), .Y(\us21\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1166_ ( .A1(\us21\/_0586_ ), .A2(\us21\/_0017_ ), .A3(\us21\/_0330_ ), .B1(\us21\/_0094_ ), .Y(\us21\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \us21/_1167_ ( .A1(\us21\/_0293_ ), .A2(\us21\/_0134_ ), .B1(\us21\/_0089_ ), .Y(\us21\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1168_ ( .A1(\us21\/_0279_ ), .A2(\us21\/_0134_ ), .B1(\us21\/_0094_ ), .Y(\us21\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1169_ ( .A(\us21\/_0368_ ), .B(\us21\/_0370_ ), .C(\us21\/_0371_ ), .D(\us21\/_0372_ ), .X(\us21\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1170_ ( .A(\us21\/_0351_ ), .B(\us21\/_0359_ ), .C(\us21\/_0367_ ), .D(\us21\/_0373_ ), .X(\us21\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1171_ ( .A1(\us21\/_0102_ ), .A2(\us21\/_0347_ ), .B1(\us21\/_0109_ ), .C1(\us21\/_0247_ ), .Y(\us21\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1172_ ( .A1(\us21\/_0102_ ), .A2(\us21\/_0347_ ), .B1(\us21\/_0532_ ), .C1(\us21\/_0247_ ), .Y(\us21\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1173_ ( .A1(\us21\/_0050_ ), .A2(\us21\/_0249_ ), .B1(\us21\/_0380_ ), .C1(\us21\/_0247_ ), .Y(\us21\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1174_ ( .A(\us21\/_0041_ ), .B(\us21\/_0375_ ), .C(\us21\/_0376_ ), .D(\us21\/_0377_ ), .X(\us21\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1175_ ( .A(\us21\/_0047_ ), .B(\us21\/_0750_ ), .X(\us21\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1176_ ( .A(\us21\/_0379_ ), .Y(\us21\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1177_ ( .A(\us21\/_0016_ ), .B(\us21\/_0608_ ), .Y(\us21\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1178_ ( .A(\us21\/_0752_ ), .B(\us21\/_0554_ ), .Y(\us21\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1179_ ( .A1(\sa21\[1\] ), .A2(\us21\/_0734_ ), .B1(\us21\/_0109_ ), .C1(\us21\/_0016_ ), .Y(\us21\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1180_ ( .A(\us21\/_0381_ ), .B(\us21\/_0382_ ), .C(\us21\/_0383_ ), .D(\us21\/_0384_ ), .X(\us21\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us21/_1181_ ( .A(\us21\/_0086_ ), .B_N(\us21\/_0736_ ), .X(\us21\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1182_ ( .A1(\us21\/_0748_ ), .A2(\us21\/_0134_ ), .B1(\us21\/_0739_ ), .Y(\us21\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1183_ ( .A1(\us21\/_0118_ ), .A2(\us21\/_0249_ ), .B1(\us21\/_0109_ ), .C1(\us21\/_0739_ ), .Y(\us21\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1184_ ( .A1(\us21\/_0102_ ), .A2(\us21\/_0301_ ), .B1(\sa21\[3\] ), .C1(\us21\/_0739_ ), .Y(\us21\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1185_ ( .A(\us21\/_0386_ ), .B(\us21\/_0387_ ), .C(\us21\/_0388_ ), .D(\us21\/_0389_ ), .X(\us21\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1186_ ( .A(\us21\/_0020_ ), .Y(\us21\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1187_ ( .A(\us21\/_0727_ ), .Y(\us21\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1188_ ( .A(\us21\/_0727_ ), .B(\us21\/_0064_ ), .Y(\us21\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1189_ ( .A1(\us21\/_0102_ ), .A2(\us21\/_0734_ ), .B1(\us21\/_0532_ ), .C1(\us21\/_0727_ ), .Y(\us21\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us21/_1190_ ( .A1(\us21\/_0392_ ), .A2(\us21\/_0393_ ), .B1(\us21\/_0394_ ), .C1(\us21\/_0395_ ), .X(\us21\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1191_ ( .A(\us21\/_0378_ ), .B(\us21\/_0385_ ), .C(\us21\/_0390_ ), .D(\us21\/_0396_ ), .X(\us21\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us21/_1192_ ( .A(\us21\/_0340_ ), .B(\us21\/_0374_ ), .C(\us21\/_0397_ ), .Y(\us21\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1193_ ( .A(\us21\/_0077_ ), .B(\us21\/_0129_ ), .X(\us21\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_1194_ ( .A(\us21\/_0398_ ), .B(\us21\/_0239_ ), .Y(\us21\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1195_ ( .A(\us21\/_0022_ ), .B(\us21\/_0111_ ), .X(\us21\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us21/_1196_ ( .A_N(\us21\/_0400_ ), .B(\us21\/_0231_ ), .Y(\us21\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us21/_1197_ ( .A(\us21\/_0399_ ), .SLEEP(\us21\/_0402_ ), .X(\us21\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_1198_ ( .A(\us21\/_0747_ ), .B(\us21\/_0251_ ), .Y(\us21\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us21/_1199_ ( .A_N(\us21\/_0404_ ), .B(\us21\/_0752_ ), .Y(\us21\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us21/_1200_ ( .A(\us21\/_0467_ ), .B(\us21\/_0194_ ), .C(\us21\/_0694_ ), .X(\us21\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us21/_1201_ ( .A_N(\us21\/_0175_ ), .B(\us21\/_0406_ ), .X(\us21\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1202_ ( .A(\us21\/_0407_ ), .Y(\us21\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1203_ ( .A1(\us21\/_0094_ ), .A2(\us21\/_0197_ ), .B1(\us21\/_0114_ ), .B2(\us21\/_0640_ ), .Y(\us21\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1204_ ( .A(\us21\/_0403_ ), .B(\us21\/_0405_ ), .C(\us21\/_0408_ ), .D(\us21\/_0409_ ), .X(\us21\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1205_ ( .A(\us21\/_0030_ ), .B(\us21\/_0150_ ), .Y(\us21\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us21/_1206_ ( .A_N(\us21\/_0169_ ), .B(\us21\/_0289_ ), .C(\us21\/_0411_ ), .X(\us21\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us21/_1207_ ( .A1(\us21\/_0467_ ), .A2(\us21\/_0151_ ), .B1(\us21\/_0140_ ), .C1(\us21\/_0129_ ), .X(\us21\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1208_ ( .A1(\us21\/_0608_ ), .A2(\us21\/_0099_ ), .B1(\us21\/_0037_ ), .C1(\us21\/_0414_ ), .Y(\us21\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1209_ ( .A(\us21\/_0738_ ), .Y(\us21\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1210_ ( .A(\us21\/_0586_ ), .B(\us21\/_0736_ ), .Y(\us21\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1211_ ( .A1(\us21\/_0194_ ), .A2(\us21\/_0038_ ), .B1(\us21\/_0118_ ), .C1(\us21\/_0153_ ), .Y(\us21\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us21/_1212_ ( .A1(\us21\/_0416_ ), .A2(\us21\/_0117_ ), .B1(\us21\/_0417_ ), .C1(\us21\/_0418_ ), .X(\us21\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1213_ ( .A(\us21\/_0077_ ), .B(\us21\/_0035_ ), .X(\us21\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1214_ ( .A(\us21\/_0662_ ), .B(\us21\/_0124_ ), .Y(\us21\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1215_ ( .A(\us21\/_0030_ ), .B(\us21\/_0137_ ), .Y(\us21\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1216_ ( .A(\us21\/_0072_ ), .B(\us21\/_0731_ ), .Y(\us21\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us21/_1217_ ( .A_N(\us21\/_0420_ ), .B(\us21\/_0421_ ), .C(\us21\/_0422_ ), .D(\us21\/_0424_ ), .X(\us21\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1218_ ( .A(\us21\/_0413_ ), .B(\us21\/_0415_ ), .C(\us21\/_0419_ ), .D(\us21\/_0425_ ), .X(\us21\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us21/_1219_ ( .A(\us21\/_0355_ ), .B(\us21\/_0102_ ), .C(\us21\/_0109_ ), .Y(\us21\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1220_ ( .A(\us21\/_0077_ ), .B(\us21\/_0017_ ), .X(\us21\/_0428_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1221_ ( .A(\us21\/_0077_ ), .B(\us21\/_0554_ ), .X(\us21\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us21/_1222_ ( .A1(\us21\/_0050_ ), .A2(\us21\/_0205_ ), .B1(\us21\/_0380_ ), .C1(\us21\/_0078_ ), .X(\us21\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us21/_1223_ ( .A(\us21\/_0428_ ), .B(\us21\/_0429_ ), .C(\us21\/_0430_ ), .Y(\us21\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us21/_1224_ ( .A_N(\us21\/_0209_ ), .B(\us21\/_0431_ ), .X(\us21\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us21/_1225_ ( .A1(\us21\/_0215_ ), .A2(\us21\/_0404_ ), .B1(\us21\/_0427_ ), .C1(\us21\/_0432_ ), .X(\us21\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1226_ ( .A(\us21\/_0043_ ), .B(\us21\/_0058_ ), .Y(\us21\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1227_ ( .A(\us21\/_0195_ ), .B(\us21\/_0233_ ), .C(\us21\/_0320_ ), .D(\us21\/_0435_ ), .X(\us21\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1228_ ( .A(\us21\/_0261_ ), .B(\us21\/_0738_ ), .Y(\us21\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1229_ ( .A1(\us21\/_0218_ ), .A2(\us21\/_0640_ ), .B1(\us21\/_0261_ ), .B2(\us21\/_0056_ ), .Y(\us21\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1230_ ( .A(\us21\/_0436_ ), .B(\us21\/_0394_ ), .C(\us21\/_0437_ ), .D(\us21\/_0438_ ), .X(\us21\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1231_ ( .A(\us21\/_0410_ ), .B(\us21\/_0426_ ), .C(\us21\/_0433_ ), .D(\us21\/_0439_ ), .X(\us21\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us21/_1232_ ( .A(\us21\/_0135_ ), .SLEEP(\us21\/_0273_ ), .X(\us21\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1233_ ( .A1(\us21\/_0279_ ), .A2(\us21\/_0134_ ), .B1(\us21\/_0099_ ), .Y(\us21\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1234_ ( .A(\us21\/_0441_ ), .B(\us21\/_0164_ ), .C(\us21\/_0270_ ), .D(\us21\/_0442_ ), .X(\us21\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1235_ ( .A(\us21\/_0051_ ), .B(\us21\/_0662_ ), .Y(\us21\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1236_ ( .A(\us21\/_0051_ ), .B(\us21\/_0271_ ), .Y(\us21\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1237_ ( .A(\us21\/_0444_ ), .B(\us21\/_0446_ ), .X(\us21\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1238_ ( .A(\us21\/_0193_ ), .B(\us21\/_0304_ ), .X(\us21\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1239_ ( .A(\us21\/_0448_ ), .Y(\us21\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1240_ ( .A(\us21\/_0162_ ), .B(\us21\/_0130_ ), .X(\us21\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1241_ ( .A(\us21\/_0450_ ), .Y(\us21\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1242_ ( .A1(\us21\/_0129_ ), .A2(\us21\/_0554_ ), .B1(\us21\/_0043_ ), .Y(\us21\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1243_ ( .A(\us21\/_0447_ ), .B(\us21\/_0449_ ), .C(\us21\/_0451_ ), .D(\us21\/_0452_ ), .X(\us21\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1244_ ( .A(\us21\/_0056_ ), .B(\us21\/_0064_ ), .Y(\us21\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us21/_1245_ ( .A_N(\us21\/_0248_ ), .B(\us21\/_0454_ ), .C(\us21\/_0254_ ), .D(\us21\/_0256_ ), .X(\us21\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1246_ ( .A1(\us21\/_0330_ ), .A2(\us21\/_0099_ ), .B1(\us21\/_0134_ ), .B2(\us21\/_0705_ ), .Y(\us21\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1247_ ( .A1(\us21\/_0748_ ), .A2(\us21\/_0738_ ), .B1(\us21\/_0092_ ), .B2(\us21\/_0752_ ), .Y(\us21\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1248_ ( .A1(\us21\/_0072_ ), .A2(\us21\/_0035_ ), .B1(\us21\/_0748_ ), .B2(\us21\/_0056_ ), .Y(\us21\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1249_ ( .A1(\us21\/_0748_ ), .A2(\us21\/_0251_ ), .B1(\us21\/_0247_ ), .Y(\us21\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1250_ ( .A(\us21\/_0457_ ), .B(\us21\/_0458_ ), .C(\us21\/_0459_ ), .D(\us21\/_0460_ ), .X(\us21\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1251_ ( .A(\us21\/_0443_ ), .B(\us21\/_0453_ ), .C(\us21\/_0455_ ), .D(\us21\/_0461_ ), .X(\us21\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1252_ ( .A(\us21\/_0705_ ), .B(\us21\/_0079_ ), .X(\us21\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1253_ ( .A(\us21\/_0586_ ), .B(\us21\/_0124_ ), .Y(\us21\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1254_ ( .A(\us21\/_0218_ ), .B(\us21\/_0747_ ), .Y(\us21\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us21/_1255_ ( .A_N(\us21\/_0463_ ), .B(\us21\/_0464_ ), .C(\us21\/_0465_ ), .X(\us21\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us21/_1256_ ( .A1(\us21\/_0271_ ), .A2(\us21\/_0072_ ), .B1(\us21\/_0142_ ), .B2(\us21\/_0027_ ), .X(\us21\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1257_ ( .A1(\us21\/_0144_ ), .A2(\us21\/_0099_ ), .B1(\us21\/_0360_ ), .C1(\us21\/_0468_ ), .Y(\us21\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us21/_1258_ ( .A1(\us21\/_0662_ ), .A2(\us21\/_0251_ ), .B1(\us21\/_0218_ ), .X(\us21\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1259_ ( .A1(\us21\/_0575_ ), .A2(\us21\/_0056_ ), .B1(\us21\/_0379_ ), .C1(\us21\/_0470_ ), .Y(\us21\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1260_ ( .A(\us21\/_0466_ ), .B(\us21\/_0469_ ), .C(\us21\/_0471_ ), .D(\us21\/_0305_ ), .X(\us21\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us21/_1261_ ( .A1(\us21\/_0247_ ), .A2(\us21\/_0683_ ), .B1(\us21\/_0324_ ), .B2(\us21\/_0056_ ), .X(\us21\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1262_ ( .A(\us21\/_0084_ ), .B(\us21\/_0099_ ), .X(\us21\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us21/_1263_ ( .A1(\us21\/_0092_ ), .A2(\us21\/_0247_ ), .B1(\us21\/_0474_ ), .X(\us21\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us21/_1264_ ( .A(\us21\/_0075_ ), .B(\us21\/_0473_ ), .C(\us21\/_0475_ ), .Y(\us21\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1265_ ( .A1(\us21\/_0279_ ), .A2(\us21\/_0255_ ), .B1(\us21\/_0084_ ), .B2(\us21\/_0060_ ), .Y(\us21\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1266_ ( .A1(\us21\/_0093_ ), .A2(\us21\/_0056_ ), .B1(\us21\/_0134_ ), .B2(\us21\/_0114_ ), .Y(\us21\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1267_ ( .A1(\us21\/_0161_ ), .A2(\us21\/_0032_ ), .B1(\us21\/_0324_ ), .B2(\us21\/_0147_ ), .Y(\us21\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1268_ ( .A1(\us21\/_0054_ ), .A2(\us21\/_0731_ ), .B1(\us21\/_0748_ ), .B2(\us21\/_0304_ ), .Y(\us21\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1269_ ( .A(\us21\/_0477_ ), .B(\us21\/_0479_ ), .C(\us21\/_0480_ ), .D(\us21\/_0481_ ), .X(\us21\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1270_ ( .A(\us21\/_0161_ ), .B(\us21\/_0064_ ), .Y(\us21\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us21/_1271_ ( .A(\us21\/_0731_ ), .B(\us21\/_0123_ ), .C(\us21\/_0467_ ), .Y(\us21\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1272_ ( .A(\us21\/_0483_ ), .B(\us21\/_0484_ ), .Y(\us21\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1273_ ( .A(\us21\/_0297_ ), .Y(\us21\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us21/_1274_ ( .A_N(\us21\/_0485_ ), .B(\us21\/_0181_ ), .C(\us21\/_0486_ ), .D(\us21\/_0386_ ), .X(\us21\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1275_ ( .A(\us21\/_0472_ ), .B(\us21\/_0476_ ), .C(\us21\/_0482_ ), .D(\us21\/_0487_ ), .X(\us21\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \us21/_1276_ ( .A(\us21\/_0440_ ), .B(\us21\/_0462_ ), .C(\us21\/_0488_ ), .Y(\us21\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1277_ ( .A(\us21\/_0403_ ), .B(\us21\/_0230_ ), .C(\us21\/_0451_ ), .D(\us21\/_0361_ ), .X(\us21\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1278_ ( .A1(\us21\/_0118_ ), .A2(\us21\/_0050_ ), .B1(\us21\/_0109_ ), .C1(\us21\/_0139_ ), .Y(\us21\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1279_ ( .A(\us21\/_0447_ ), .B(\us21\/_0437_ ), .C(\us21\/_0491_ ), .D(\us21\/_0427_ ), .X(\us21\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1280_ ( .A1(\us21\/_0084_ ), .A2(\us21\/_0255_ ), .B1(\us21\/_0608_ ), .B2(\us21\/_0247_ ), .Y(\us21\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1281_ ( .A1(\us21\/_0144_ ), .A2(\us21\/_0147_ ), .B1(\us21\/_0355_ ), .B2(\us21\/_0093_ ), .Y(\us21\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1282_ ( .A1(\us21\/_0705_ ), .A2(\us21\/_0279_ ), .B1(\us21\/_0330_ ), .B2(\us21\/_0247_ ), .Y(\us21\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1283_ ( .A1(\us21\/_0279_ ), .A2(\us21\/_0084_ ), .B1(\us21\/_0114_ ), .Y(\us21\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1284_ ( .A(\us21\/_0493_ ), .B(\us21\/_0494_ ), .C(\us21\/_0495_ ), .D(\us21\/_0496_ ), .X(\us21\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1285_ ( .A1(\us21\/_0134_ ), .A2(\us21\/_0137_ ), .B1(\us21\/_0355_ ), .B2(\us21\/_0575_ ), .Y(\us21\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1286_ ( .A1(\us21\/_0099_ ), .A2(\us21\/_0733_ ), .B1(\us21\/_0093_ ), .B2(\us21\/_0218_ ), .Y(\us21\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1287_ ( .A(\us21\/_0147_ ), .B(\us21\/_0640_ ), .Y(\us21\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1288_ ( .A1(\us21\/_0153_ ), .A2(\us21\/_0056_ ), .B1(\us21\/_0748_ ), .Y(\us21\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1289_ ( .A(\us21\/_0498_ ), .B(\us21\/_0500_ ), .C(\us21\/_0501_ ), .D(\us21\/_0502_ ), .X(\us21\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1290_ ( .A(\us21\/_0490_ ), .B(\us21\/_0492_ ), .C(\us21\/_0497_ ), .D(\us21\/_0503_ ), .X(\us21\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us21/_1291_ ( .A_N(\us21\/_0275_ ), .B(\us21\/_0705_ ), .X(\us21\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1292_ ( .A(\us21\/_0505_ ), .Y(\us21\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1293_ ( .A(\us21\/_0380_ ), .B(\us21\/_0347_ ), .X(\us21\/_0507_ ) );
sky130_fd_sc_hd__o21ai_1 \us21/_1294_ ( .A1(\us21\/_0507_ ), .A2(\us21\/_0093_ ), .B1(\us21\/_0056_ ), .Y(\us21\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1295_ ( .A(\us21\/_0322_ ), .B(\us21\/_0277_ ), .C(\us21\/_0506_ ), .D(\us21\/_0508_ ), .X(\us21\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1296_ ( .A(\us21\/_0084_ ), .B(\us21\/_0705_ ), .X(\us21\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1297_ ( .A1(\us21\/_0733_ ), .A2(\us21\/_0114_ ), .B1(\us21\/_0429_ ), .C1(\us21\/_0511_ ), .Y(\us21\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_1298_ ( .A(\us21\/_0019_ ), .B(\us21\/_0024_ ), .Y(\us21\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1299_ ( .A(\us21\/_0512_ ), .B(\us21\/_0513_ ), .C(\us21\/_0742_ ), .D(\us21\/_0306_ ), .X(\us21\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1300_ ( .A1(\us21\/_0532_ ), .A2(\us21\/_0089_ ), .B1(\us21\/_0154_ ), .C1(\us21\/_0169_ ), .Y(\us21\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us21/_1301_ ( .A1(\us21\/_0749_ ), .A2(\us21\/_0026_ ), .B1(\us21\/_0069_ ), .C1(\us21\/_0032_ ), .X(\us21\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us21/_1302_ ( .A1(\us21\/_0324_ ), .A2(\us21\/_0355_ ), .B1(\us21\/_0330_ ), .B2(\us21\/_0727_ ), .X(\us21\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us21/_1303_ ( .A(\us21\/_0133_ ), .B(\us21\/_0516_ ), .C(\us21\/_0517_ ), .Y(\us21\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1304_ ( .A(\us21\/_0509_ ), .B(\us21\/_0514_ ), .C(\us21\/_0515_ ), .D(\us21\/_0518_ ), .X(\us21\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1305_ ( .A(\us21\/_0747_ ), .B(\us21\/_0072_ ), .Y(\us21\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1306_ ( .A1(\us21\/_0082_ ), .A2(\us21\/_0070_ ), .B1(\us21\/_0043_ ), .B2(\us21\/_0193_ ), .Y(\us21\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1307_ ( .A(\us21\/_0311_ ), .B(\us21\/_0520_ ), .C(\us21\/_0332_ ), .D(\us21\/_0522_ ), .X(\us21\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1308_ ( .A(\us21\/_0129_ ), .B(\us21\/_0218_ ), .X(\us21\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_1309_ ( .A(\us21\/_0235_ ), .B(\us21\/_0524_ ), .Y(\us21\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us21/_1310_ ( .A(\us21\/_0081_ ), .B(\us21\/_0085_ ), .Y(\us21\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1311_ ( .A1(\us21\/_0051_ ), .A2(\us21\/_0045_ ), .B1(\us21\/_0130_ ), .B2(\us21\/_0094_ ), .Y(\us21\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1312_ ( .A(\us21\/_0523_ ), .B(\us21\/_0525_ ), .C(\us21\/_0526_ ), .D(\us21\/_0527_ ), .X(\us21\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us21/_1313_ ( .A_N(\us21\/_0250_ ), .B(\us21\/_0521_ ), .Y(\us21\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1314_ ( .A(\us21\/_0128_ ), .B(\us21\/_0020_ ), .X(\us21\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1315_ ( .A(\us21\/_0530_ ), .Y(\us21\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1316_ ( .A(\us21\/_0099_ ), .B(\us21\/_0058_ ), .X(\us21\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1317_ ( .A(\us21\/_0533_ ), .Y(\us21\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us21/_1318_ ( .A_N(\us21\/_0529_ ), .B(\us21\/_0531_ ), .C(\us21\/_0534_ ), .D(\us21\/_0192_ ), .X(\us21\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1319_ ( .A(\us21\/_0434_ ), .B(\us21\/_0078_ ), .X(\us21\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us21/_1320_ ( .A1(\us21\/_0750_ ), .A2(\us21\/_0079_ ), .B1(\us21\/_0129_ ), .B2(\us21\/_0705_ ), .X(\us21\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1321_ ( .A1(\us21\/_0161_ ), .A2(\us21\/_0032_ ), .B1(\us21\/_0536_ ), .C1(\us21\/_0537_ ), .Y(\us21\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us21/_1322_ ( .A1(\us21\/_0747_ ), .A2(\us21\/_0162_ ), .B1(\us21\/_0079_ ), .B2(\us21\/_0043_ ), .X(\us21\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1323_ ( .A1(\us21\/_0093_ ), .A2(\us21\/_0247_ ), .B1(\us21\/_0240_ ), .C1(\us21\/_0539_ ), .Y(\us21\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1324_ ( .A(\us21\/_0434_ ), .B(\us21\/_0043_ ), .X(\us21\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us21/_1325_ ( .A1(\us21\/_0142_ ), .A2(\us21\/_0150_ ), .B1(\us21\/_0022_ ), .B2(\us21\/_0137_ ), .X(\us21\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1326_ ( .A1(\us21\/_0279_ ), .A2(\us21\/_0051_ ), .B1(\us21\/_0541_ ), .C1(\us21\/_0542_ ), .Y(\us21\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1327_ ( .A(\us21\/_0159_ ), .B(\us21\/_0035_ ), .X(\us21\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us21/_1328_ ( .A1(\us21\/_0271_ ), .A2(\us21\/_0434_ ), .B1(\us21\/_0027_ ), .X(\us21\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1329_ ( .A1(\us21\/_0091_ ), .A2(\us21\/_0128_ ), .B1(\us21\/_0545_ ), .C1(\us21\/_0546_ ), .Y(\us21\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1330_ ( .A(\us21\/_0538_ ), .B(\us21\/_0540_ ), .C(\us21\/_0544_ ), .D(\us21\/_0547_ ), .X(\us21\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1331_ ( .A(\us21\/_0099_ ), .B(\us21\/_0193_ ), .X(\us21\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us21/_1332_ ( .A(\us21\/_0549_ ), .B(\us21\/_0186_ ), .C(\us21\/_0187_ ), .Y(\us21\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1333_ ( .A(\us21\/_0062_ ), .B(\us21\/_0347_ ), .C(\us21\/_0749_ ), .D(\us21\/_0694_ ), .X(\us21\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1334_ ( .A1(\us21\/_0130_ ), .A2(\us21\/_0218_ ), .B1(\us21\/_0551_ ), .C1(\us21\/_0101_ ), .Y(\us21\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1335_ ( .A(\us21\/_0139_ ), .B(\us21\/_0640_ ), .Y(\us21\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1336_ ( .A1(\us21\/_0752_ ), .A2(\us21\/_0662_ ), .B1(\us21\/_0084_ ), .B2(\us21\/_0099_ ), .Y(\us21\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1337_ ( .A(\us21\/_0550_ ), .B(\us21\/_0552_ ), .C(\us21\/_0553_ ), .D(\us21\/_0555_ ), .X(\us21\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1338_ ( .A(\us21\/_0528_ ), .B(\us21\/_0535_ ), .C(\us21\/_0548_ ), .D(\us21\/_0556_ ), .X(\us21\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us21/_1339_ ( .A(\us21\/_0504_ ), .B(\us21\/_0519_ ), .C(\us21\/_0557_ ), .Y(\us21\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1340_ ( .A(\us21\/_0054_ ), .B(\us21\/_0507_ ), .X(\us21\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us21/_1341_ ( .A_N(\us21\/_0558_ ), .B(\us21\/_0408_ ), .C(\us21\/_0451_ ), .D(\us21\/_0452_ ), .X(\us21\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1342_ ( .A(\us21\/_0549_ ), .Y(\us21\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1343_ ( .A(\us21\/_0559_ ), .B(\us21\/_0403_ ), .C(\us21\/_0560_ ), .D(\us21\/_0371_ ), .X(\us21\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1344_ ( .A(\us21\/_0181_ ), .B(\us21\/_0178_ ), .X(\us21\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1345_ ( .A(\us21\/_0562_ ), .B(\us21\/_0552_ ), .C(\us21\/_0553_ ), .D(\us21\/_0555_ ), .X(\us21\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1346_ ( .A(\us21\/_0247_ ), .B(\us21\/_0020_ ), .Y(\us21\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1347_ ( .A(\us21\/_0051_ ), .B(\us21\/_0130_ ), .X(\us21\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1348_ ( .A(\us21\/_0566_ ), .Y(\us21\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1349_ ( .A(\us21\/_0159_ ), .B(\us21\/_0412_ ), .X(\us21\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1350_ ( .A1(\us21\/_0752_ ), .A2(\us21\/_0640_ ), .B1(\us21\/_0568_ ), .B2(\us21\/_0175_ ), .Y(\us21\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1351_ ( .A(\us21\/_0076_ ), .B(\us21\/_0565_ ), .C(\us21\/_0567_ ), .D(\us21\/_0569_ ), .X(\us21\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us21/_1352_ ( .A1(\us21\/_0035_ ), .A2(\us21\/_0142_ ), .B1(\us21\/_0161_ ), .X(\us21\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1353_ ( .A(\us21\/_0099_ ), .B(\us21\/_0662_ ), .Y(\us21\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us21/_1354_ ( .A(\us21\/_0420_ ), .B(\us21\/_0571_ ), .C_N(\us21\/_0572_ ), .Y(\us21\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1355_ ( .A(\us21\/_0051_ ), .B(\us21\/_0747_ ), .Y(\us21\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1356_ ( .A(\us21\/_0574_ ), .B(\us21\/_0319_ ), .C(\us21\/_0320_ ), .D(\us21\/_0411_ ), .X(\us21\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1357_ ( .A(\us21\/_0736_ ), .B(\us21\/_0035_ ), .Y(\us21\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1358_ ( .A(\us21\/_0736_ ), .B(\us21\/_0030_ ), .Y(\us21\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1359_ ( .A(\us21\/_0298_ ), .B(\us21\/_0208_ ), .C(\us21\/_0577_ ), .D(\us21\/_0578_ ), .X(\us21\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1360_ ( .A1(\us21\/_0020_ ), .A2(\us21\/_0137_ ), .B1(\us21\/_0261_ ), .B2(\us21\/_0128_ ), .Y(\us21\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1361_ ( .A(\us21\/_0573_ ), .B(\us21\/_0576_ ), .C(\us21\/_0579_ ), .D(\us21\/_0580_ ), .X(\us21\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1362_ ( .A(\us21\/_0561_ ), .B(\us21\/_0563_ ), .C(\us21\/_0570_ ), .D(\us21\/_0581_ ), .X(\us21\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1363_ ( .A(\us21\/_0128_ ), .B(\us21\/_0193_ ), .X(\us21\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1364_ ( .A(\us21\/_0082_ ), .B(\us21\/_0162_ ), .X(\us21\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us21/_1365_ ( .A(\us21\/_0583_ ), .B(\us21\/_0584_ ), .C_N(\us21\/_0437_ ), .Y(\us21\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us21/_1366_ ( .A(\us21\/_0150_ ), .B(\us21\/_0118_ ), .C(\us21\/_0380_ ), .Y(\us21\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us21/_1367_ ( .A_N(\us21\/_0182_ ), .B(\us21\/_0587_ ), .C(\us21\/_0323_ ), .X(\us21\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1368_ ( .A1(\us21\/_0575_ ), .A2(\us21\/_0153_ ), .B1(\us21\/_0727_ ), .B2(\us21\/_0058_ ), .Y(\us21\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1369_ ( .A1(\us21\/_0218_ ), .A2(\us21\/_0064_ ), .B1(\us21\/_0134_ ), .B2(\us21\/_0255_ ), .Y(\us21\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1370_ ( .A(\us21\/_0585_ ), .B(\us21\/_0588_ ), .C(\us21\/_0589_ ), .D(\us21\/_0590_ ), .X(\us21\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us21/_1371_ ( .A1(\us21\/_0091_ ), .A2(\us21\/_0139_ ), .B1(\us21\/_0250_ ), .Y(\us21\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1372_ ( .A1(\us21\/_0092_ ), .A2(\us21\/_0739_ ), .B1(\us21\/_0324_ ), .B2(\us21\/_0247_ ), .Y(\us21\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1373_ ( .A1(\us21\/_0144_ ), .A2(\us21\/_0153_ ), .B1(\us21\/_0683_ ), .B2(\us21\/_0056_ ), .Y(\us21\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1374_ ( .A1(\us21\/_0091_ ), .A2(\us21\/_0218_ ), .B1(\us21\/_0330_ ), .B2(\us21\/_0056_ ), .Y(\us21\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1375_ ( .A(\us21\/_0592_ ), .B(\us21\/_0593_ ), .C(\us21\/_0594_ ), .D(\us21\/_0595_ ), .X(\us21\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1376_ ( .A(\us21\/_0218_ ), .B(\us21\/_0144_ ), .Y(\us21\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1377_ ( .A(\us21\/_0312_ ), .B(\us21\/_0598_ ), .Y(\us21\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1378_ ( .A(\us21\/_0575_ ), .B(\us21\/_0147_ ), .Y(\us21\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1379_ ( .A1(\us21\/_0293_ ), .A2(\us21\/_0137_ ), .B1(\us21\/_0093_ ), .B2(\us21\/_0739_ ), .Y(\us21\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1380_ ( .A1(\us21\/_0734_ ), .A2(\us21\/_0531_ ), .B1(\us21\/_0600_ ), .C1(\us21\/_0601_ ), .Y(\us21\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1381_ ( .A1(\us21\/_0153_ ), .A2(\us21\/_0261_ ), .B1(\us21\/_0599_ ), .C1(\us21\/_0602_ ), .Y(\us21\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1382_ ( .A(\us21\/_0591_ ), .B(\us21\/_0596_ ), .C(\us21\/_0174_ ), .D(\us21\/_0603_ ), .X(\us21\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1383_ ( .A(\us21\/_0247_ ), .B(\us21\/_0144_ ), .Y(\us21\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1384_ ( .A(\us21\/_0113_ ), .B(\us21\/_0017_ ), .Y(\us21\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1385_ ( .A(\us21\/_0381_ ), .B(\us21\/_0605_ ), .C(\us21\/_0361_ ), .D(\us21\/_0606_ ), .X(\us21\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1386_ ( .A1(\us21\/_0016_ ), .A2(\us21\/_0727_ ), .B1(\us21\/_0733_ ), .Y(\us21\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1387_ ( .A1(\us21\/_0586_ ), .A2(\us21\/_0159_ ), .B1(\us21\/_0082_ ), .B2(\us21\/_0750_ ), .Y(\us21\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1388_ ( .A1(\us21\/_0142_ ), .A2(\us21\/_0162_ ), .B1(\us21\/_0079_ ), .B2(\us21\/_0054_ ), .Y(\us21\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1389_ ( .A(\us21\/_0610_ ), .B(\us21\/_0611_ ), .C(\us21\/_0105_ ), .D(\us21\/_0106_ ), .X(\us21\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1390_ ( .A1(\us21\/_0094_ ), .A2(\us21\/_0302_ ), .B1(\us21\/_0324_ ), .B2(\us21\/_0089_ ), .Y(\us21\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1391_ ( .A(\us21\/_0607_ ), .B(\us21\/_0609_ ), .C(\us21\/_0612_ ), .D(\us21\/_0613_ ), .X(\us21\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1392_ ( .A(\us21\/_0041_ ), .B(\us21\/_0170_ ), .X(\us21\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1393_ ( .A(\us21\/_0554_ ), .B(\us21\/_0027_ ), .X(\us21\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1394_ ( .A(\us21\/_0027_ ), .B(\us21\/_0261_ ), .Y(\us21\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us21/_1395_ ( .A_N(\us21\/_0616_ ), .B(\us21\/_0617_ ), .Y(\us21\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1396_ ( .A1(\us21\/_0147_ ), .A2(\us21\/_0302_ ), .B1(\us21\/_0342_ ), .C1(\us21\/_0618_ ), .Y(\us21\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1397_ ( .A(\us21\/_0614_ ), .B(\us21\/_0272_ ), .C(\us21\/_0615_ ), .D(\us21\/_0620_ ), .X(\us21\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us21/_1398_ ( .A(\us21\/_0582_ ), .B(\us21\/_0604_ ), .C(\us21\/_0621_ ), .Y(\us21\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1399_ ( .A1(\us21\/_0084_ ), .A2(\us21\/_0134_ ), .B1(\us21\/_0089_ ), .Y(\us21\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1400_ ( .A1(\us21\/_0144_ ), .A2(\us21\/_0608_ ), .A3(\us21\/_0330_ ), .B1(\us21\/_0089_ ), .Y(\us21\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1401_ ( .A1(\us21\/_0197_ ), .A2(\us21\/_0130_ ), .A3(\us21\/_0110_ ), .B1(\us21\/_0094_ ), .Y(\us21\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1402_ ( .A(\us21\/_0432_ ), .B(\us21\/_0622_ ), .C(\us21\/_0623_ ), .D(\us21\/_0624_ ), .X(\us21\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us21/_1403_ ( .A1(\us21\/_0554_ ), .A2(\us21\/_0017_ ), .A3(\us21\/_0022_ ), .B1(\us21\/_0161_ ), .X(\us21\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us21/_1404_ ( .A_N(\us21\/_0269_ ), .B(\us21\/_0170_ ), .X(\us21\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1405_ ( .A1(\us21\/_0109_ ), .A2(\us21\/_0064_ ), .A3(\us21\/_0733_ ), .B1(\us21\/_0355_ ), .Y(\us21\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us21/_1406_ ( .A_N(\us21\/_0626_ ), .B(\us21\/_0627_ ), .C(\us21\/_0353_ ), .D(\us21\/_0628_ ), .X(\us21\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1407_ ( .A1(\us21\/_0091_ ), .A2(\us21\/_0110_ ), .A3(\us21\/_0176_ ), .B1(\us21\/_0139_ ), .Y(\us21\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1408_ ( .A1(\us21\/_0020_ ), .A2(\us21\/_0261_ ), .B1(\us21\/_0147_ ), .Y(\us21\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1409_ ( .A(\us21\/_0631_ ), .B(\us21\/_0344_ ), .C(\us21\/_0421_ ), .D(\us21\/_0632_ ), .X(\us21\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us21/_1410_ ( .A1(\us21\/_0325_ ), .A2(\us21\/_0734_ ), .B1(\us21\/_0038_ ), .C1(\us21\/_0113_ ), .X(\us21\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1411_ ( .A1(\us21\/_0134_ ), .A2(\us21\/_0114_ ), .B1(\us21\/_0221_ ), .C1(\us21\/_0634_ ), .Y(\us21\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us21/_1412_ ( .A(\us21\/_0119_ ), .B_N(\us21\/_0111_ ), .Y(\us21\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1413_ ( .A1(\us21\/_0032_ ), .A2(\us21\/_0113_ ), .B1(\us21\/_0636_ ), .C1(\us21\/_0400_ ), .Y(\us21\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1414_ ( .A1(\us21\/_0731_ ), .A2(\us21\/_0293_ ), .A3(\us21\/_0251_ ), .B1(\us21\/_0099_ ), .Y(\us21\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1415_ ( .A(\us21\/_0189_ ), .B(\us21\/_0635_ ), .C(\us21\/_0637_ ), .D(\us21\/_0638_ ), .X(\us21\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1416_ ( .A(\us21\/_0625_ ), .B(\us21\/_0630_ ), .C(\us21\/_0633_ ), .D(\us21\/_0639_ ), .X(\us21\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1417_ ( .A(\us21\/_0747_ ), .B(\us21\/_0738_ ), .X(\us21\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1418_ ( .A(\us21\/_0736_ ), .B(\us21\/_0731_ ), .X(\us21\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us21/_1419_ ( .A_N(\us21\/_0643_ ), .B(\us21\/_0577_ ), .Y(\us21\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1420_ ( .A1(\us21\/_0084_ ), .A2(\us21\/_0739_ ), .B1(\us21\/_0642_ ), .C1(\us21\/_0644_ ), .Y(\us21\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1421_ ( .A1(\us21\/_0050_ ), .A2(\us21\/_0249_ ), .B1(\us21\/_0194_ ), .C1(\us21\/_0738_ ), .Y(\us21\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1422_ ( .A(\us21\/_0646_ ), .B(\us21\/_0232_ ), .C(\us21\/_0417_ ), .D(\us21\/_0578_ ), .X(\us21\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1423_ ( .A1(\us21\/_0064_ ), .A2(\us21\/_0733_ ), .B1(\us21\/_0727_ ), .Y(\us21\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1424_ ( .A1(\us21\/_0193_ ), .A2(\us21\/_0276_ ), .B1(\us21\/_0727_ ), .Y(\us21\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1425_ ( .A(\us21\/_0645_ ), .B(\us21\/_0647_ ), .C(\us21\/_0648_ ), .D(\us21\/_0649_ ), .X(\us21\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1426_ ( .A1(\us21\/_0325_ ), .A2(\us21\/_0734_ ), .B1(\us21\/_0038_ ), .C1(\us21\/_0247_ ), .Y(\us21\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1427_ ( .A1(\us21\/_0249_ ), .A2(\us21\/_0205_ ), .B1(\us21\/_0412_ ), .C1(\us21\/_0247_ ), .Y(\us21\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1428_ ( .A(\us21\/_0652_ ), .B(\us21\/_0653_ ), .X(\us21\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1429_ ( .A1(\us21\/_0733_ ), .A2(\us21\/_0748_ ), .A3(\us21\/_0324_ ), .B1(\us21\/_0016_ ), .Y(\us21\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1430_ ( .A1(\us21\/_0640_ ), .A2(\us21\/_0193_ ), .A3(\us21\/_0091_ ), .B1(\us21\/_0016_ ), .Y(\us21\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1431_ ( .A1(\us21\/_0102_ ), .A2(\us21\/_0301_ ), .B1(\sa21\[3\] ), .C1(\us21\/_0247_ ), .Y(\us21\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1432_ ( .A(\us21\/_0654_ ), .B(\us21\/_0655_ ), .C(\us21\/_0656_ ), .D(\us21\/_0657_ ), .X(\us21\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1433_ ( .A1(\us21\/_0118_ ), .A2(\us21\/_0050_ ), .B1(\us21\/_0038_ ), .C1(\us21\/_0478_ ), .Y(\us21\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us21/_1434_ ( .A_N(\us21\/_0250_ ), .B(\us21\/_0465_ ), .C(\us21\/_0659_ ), .X(\us21\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1435_ ( .A1(\us21\/_0683_ ), .A2(\us21\/_0324_ ), .B1(\us21\/_0255_ ), .Y(\us21\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1436_ ( .A1(\us21\/_0032_ ), .A2(\us21\/_0193_ ), .A3(\us21\/_0047_ ), .B1(\us21\/_0255_ ), .Y(\us21\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1437_ ( .A1(\us21\/_0144_ ), .A2(\us21\/_0586_ ), .A3(\us21\/_0047_ ), .B1(\us21\/_0218_ ), .Y(\us21\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1438_ ( .A(\us21\/_0660_ ), .B(\us21\/_0661_ ), .C(\us21\/_0663_ ), .D(\us21\/_0664_ ), .X(\us21\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1439_ ( .A1(\us21\/_0091_ ), .A2(\us21\/_0276_ ), .B1(\us21\/_0060_ ), .Y(\us21\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1440_ ( .A1(\us21\/_0144_ ), .A2(\us21\/_0608_ ), .B1(\us21\/_0056_ ), .Y(\us21\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1441_ ( .A1(\us21\/_0412_ ), .A2(\us21\/_0038_ ), .B1(\us21\/_0102_ ), .C1(\us21\/_0060_ ), .Y(\us21\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1442_ ( .A1(\sa21\[1\] ), .A2(\us21\/_0734_ ), .B1(\us21\/_0109_ ), .C1(\us21\/_0056_ ), .Y(\us21\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1443_ ( .A(\us21\/_0666_ ), .B(\us21\/_0667_ ), .C(\us21\/_0668_ ), .D(\us21\/_0669_ ), .X(\us21\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1444_ ( .A(\us21\/_0650_ ), .B(\us21\/_0658_ ), .C(\us21\/_0665_ ), .D(\us21\/_0670_ ), .X(\us21\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us21/_1445_ ( .A(\us21\/_0641_ ), .B(\us21\/_0174_ ), .C(\us21\/_0671_ ), .Y(\us21\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us21/_1446_ ( .A(\us21\/_0049_ ), .B(\us21\/_0618_ ), .C_N(\us21\/_0052_ ), .Y(\us21\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us21/_1447_ ( .A(\us21\/_0239_ ), .Y(\us21\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1448_ ( .A(\us21\/_0705_ ), .B(\us21\/_0032_ ), .Y(\us21\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1449_ ( .A1(\us21\/_0054_ ), .A2(\us21\/_0731_ ), .B1(\us21\/_0035_ ), .B2(\us21\/_0705_ ), .Y(\us21\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1450_ ( .A1(\us21\/_0304_ ), .A2(\us21\/_0731_ ), .B1(\us21\/_0047_ ), .B2(\us21\/_0750_ ), .Y(\us21\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1451_ ( .A(\us21\/_0674_ ), .B(\us21\/_0675_ ), .C(\us21\/_0676_ ), .D(\us21\/_0677_ ), .X(\us21\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us21/_1452_ ( .A_N(\us21\/_0584_ ), .B(\us21\/_0283_ ), .X(\us21\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1453_ ( .A(\us21\/_0673_ ), .B(\us21\/_0678_ ), .C(\us21\/_0679_ ), .D(\us21\/_0508_ ), .X(\us21\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1454_ ( .A1(\us21\/_0016_ ), .A2(\us21\/_0733_ ), .B1(\us21\/_0355_ ), .B2(\us21\/_0092_ ), .Y(\us21\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1455_ ( .A(\us21\/_0681_ ), .B(\us21\/_0034_ ), .X(\us21\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us21/_1456_ ( .A1(\us21\/_0330_ ), .A2(\us21\/_0139_ ), .B1(\us21\/_0324_ ), .B2(\us21\/_0089_ ), .X(\us21\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1457_ ( .A1(\us21\/_0146_ ), .A2(\us21\/_0147_ ), .B1(\us21\/_0133_ ), .C1(\us21\/_0684_ ), .Y(\us21\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1458_ ( .A(\us21\/_0113_ ), .B(\us21\/_0251_ ), .Y(\us21\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us21/_1459_ ( .A_N(\us21\/_0463_ ), .B(\us21\/_0686_ ), .C(\us21\/_0383_ ), .D(\us21\/_0464_ ), .X(\us21\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1460_ ( .A1(\us21\/_0051_ ), .A2(\us21\/_0293_ ), .B1(\us21\/_0084_ ), .B2(\us21\/_0705_ ), .Y(\us21\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1461_ ( .A1(\us21\/_0017_ ), .A2(\us21\/_0072_ ), .B1(\us21\/_0134_ ), .B2(\us21\/_0078_ ), .Y(\us21\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1462_ ( .A(\us21\/_0687_ ), .B(\us21\/_0236_ ), .C(\us21\/_0688_ ), .D(\us21\/_0689_ ), .X(\us21\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1463_ ( .A(\us21\/_0680_ ), .B(\us21\/_0682_ ), .C(\us21\/_0685_ ), .D(\us21\/_0690_ ), .X(\us21\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us21/_1464_ ( .A1(\us21\/_0532_ ), .A2(\us21\/_0380_ ), .B1(\us21\/_0102_ ), .C1(\us21\/_0355_ ), .X(\us21\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us21/_1465_ ( .A(\us21\/_0692_ ), .B(\us21\/_0338_ ), .C(\us21\/_0644_ ), .Y(\us21\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1466_ ( .A(\us21\/_0016_ ), .B(\us21\/_0020_ ), .Y(\us21\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1467_ ( .A1(\us21\/_0032_ ), .A2(\us21\/_0137_ ), .B1(\us21\/_0279_ ), .B2(\us21\/_0094_ ), .Y(\us21\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1468_ ( .A1(\us21\/_0575_ ), .A2(\us21\/_0153_ ), .B1(\us21\/_0161_ ), .B2(\us21\/_0293_ ), .Y(\us21\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1469_ ( .A(\us21\/_0259_ ), .B(\us21\/_0695_ ), .C(\us21\/_0696_ ), .D(\us21\/_0697_ ), .X(\us21\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us21/_1470_ ( .A1(\us21\/_0255_ ), .A2(\us21\/_0640_ ), .B1(\us21\/_0016_ ), .B2(\us21\/_0193_ ), .X(\us21\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1471_ ( .A1(\us21\/_0060_ ), .A2(\us21\/_0176_ ), .B1(\us21\/_0699_ ), .C1(\us21\/_0177_ ), .Y(\us21\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1472_ ( .A1(\us21\/_0091_ ), .A2(\us21\/_0218_ ), .B1(\us21\/_0092_ ), .B2(\us21\/_0705_ ), .Y(\us21\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us21/_1473_ ( .A1(\us21\/_0705_ ), .A2(\us21\/_0683_ ), .B1(\us21\/_0093_ ), .B2(\us21\/_0114_ ), .Y(\us21\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us21/_1474_ ( .A1(\us21\/_0683_ ), .A2(\us21\/_0084_ ), .B1(\us21\/_0094_ ), .Y(\us21\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us21/_1475_ ( .A1(\us21\/_0249_ ), .A2(\us21\/_0205_ ), .B1(\us21\/_0038_ ), .C1(\us21\/_0056_ ), .Y(\us21\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1476_ ( .A(\us21\/_0701_ ), .B(\us21\/_0702_ ), .C(\us21\/_0703_ ), .D(\us21\/_0704_ ), .X(\us21\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1477_ ( .A(\us21\/_0693_ ), .B(\us21\/_0698_ ), .C(\us21\/_0700_ ), .D(\us21\/_0706_ ), .X(\us21\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us21/_1478_ ( .A1(\us21\/_0113_ ), .A2(\us21\/_0640_ ), .B1(\us21\/_0099_ ), .B2(\us21\/_0058_ ), .X(\us21\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us21/_1479_ ( .A(\us21\/_0407_ ), .B(\us21\/_0708_ ), .C(\us21\/_0529_ ), .Y(\us21\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1480_ ( .A(\us21\/_0568_ ), .B(\us21\/_0175_ ), .Y(\us21\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us21/_1481_ ( .A1(\us21\/_0247_ ), .A2(\us21\/_0114_ ), .A3(\us21\/_0051_ ), .B1(\us21\/_0130_ ), .Y(\us21\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1482_ ( .A(\us21\/_0709_ ), .B(\us21\/_0550_ ), .C(\us21\/_0710_ ), .D(\us21\/_0711_ ), .X(\us21\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us21/_1483_ ( .A1(\us21\/_0114_ ), .A2(\us21\/_0064_ ), .B1(\us21\/_0261_ ), .B2(\us21\/_0089_ ), .X(\us21\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1484_ ( .A1(\us21\/_0355_ ), .A2(\us21\/_0261_ ), .B1(\us21\/_0198_ ), .C1(\us21\/_0713_ ), .Y(\us21\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1485_ ( .A(\us21\/_0586_ ), .B(\us21\/_0478_ ), .Y(\us21\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us21/_1486_ ( .A_N(\us21\/_0541_ ), .B(\us21\/_0267_ ), .C(\us21\/_0715_ ), .D(\us21\/_0320_ ), .X(\us21\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1487_ ( .A(\us21\/_0586_ ), .B(\us21\/_0070_ ), .Y(\us21\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us21/_1488_ ( .A_N(\us21\/_0211_ ), .B(\us21\/_0155_ ), .C(\us21\/_0202_ ), .D(\us21\/_0718_ ), .X(\us21\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us21/_1489_ ( .A(\us21\/_0150_ ), .B(\us21\/_0205_ ), .C(\us21\/_0380_ ), .Y(\us21\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us21/_1490_ ( .A(\us21\/_0411_ ), .B(\us21\/_0720_ ), .X(\us21\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us21/_1491_ ( .A1(\us21\/_0017_ ), .A2(\us21\/_0022_ ), .B1(\us21\/_0078_ ), .X(\us21\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us21/_1492_ ( .A1(\us21\/_0134_ ), .A2(\us21\/_0738_ ), .B1(\us21\/_0101_ ), .C1(\us21\/_0722_ ), .Y(\us21\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1493_ ( .A(\us21\/_0717_ ), .B(\us21\/_0719_ ), .C(\us21\/_0721_ ), .D(\us21\/_0723_ ), .X(\us21\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us21/_1494_ ( .A(\us21\/_0739_ ), .B(\us21\/_0193_ ), .Y(\us21\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1495_ ( .A(\us21\/_0344_ ), .B(\us21\/_0184_ ), .C(\us21\/_0449_ ), .D(\us21\/_0725_ ), .X(\us21\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us21/_1496_ ( .A(\us21\/_0712_ ), .B(\us21\/_0714_ ), .C(\us21\/_0724_ ), .D(\us21\/_0726_ ), .X(\us21\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \us21/_1497_ ( .A(\us21\/_0691_ ), .B(\us21\/_0707_ ), .C(\us21\/_0728_ ), .Y(\us21\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \us22/_0753_ ( .A(\sa22\[2\] ), .B_N(\sa22\[3\] ), .Y(\us22\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \us22/_0755_ ( .A(\sa22\[1\] ), .B(\sa22\[0\] ), .X(\us22\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us22/_0756_ ( .A(\us22\/_0096_ ), .B(\us22\/_0118_ ), .X(\us22\/_0129_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0757_ ( .A(\sa22\[7\] ), .B(\sa22\[6\] ), .X(\us22\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_0758_ ( .A(\sa22\[4\] ), .B(\sa22\[5\] ), .Y(\us22\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0759_ ( .A(\us22\/_0140_ ), .B(\us22\/_0151_ ), .X(\us22\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0761_ ( .A(\us22\/_0129_ ), .B(\us22\/_0162_ ), .X(\us22\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0762_ ( .A(\us22\/_0096_ ), .X(\us22\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \us22/_0763_ ( .A(\sa22\[1\] ), .B_N(\sa22\[0\] ), .Y(\us22\/_0205_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0764_ ( .A(\us22\/_0205_ ), .X(\us22\/_0216_ ) );
sky130_fd_sc_hd__and3_1 \us22/_0765_ ( .A(\us22\/_0162_ ), .B(\us22\/_0194_ ), .C(\us22\/_0216_ ), .X(\us22\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us22/_0766_ ( .A(\us22\/_0183_ ), .SLEEP(\us22\/_0227_ ), .X(\us22\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \us22/_0767_ ( .A(\sa22\[0\] ), .B_N(\sa22\[1\] ), .Y(\us22\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_0768_ ( .A(\sa22\[2\] ), .B(\sa22\[3\] ), .Y(\us22\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0769_ ( .A(\us22\/_0249_ ), .B(\us22\/_0260_ ), .X(\us22\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0771_ ( .A(\us22\/_0271_ ), .X(\us22\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0772_ ( .A(\us22\/_0162_ ), .X(\us22\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_0773_ ( .A(\us22\/_0293_ ), .B(\us22\/_0304_ ), .Y(\us22\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us22/_0774_ ( .A(\sa22\[1\] ), .Y(\us22\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us22/_0776_ ( .A(\sa22\[0\] ), .Y(\us22\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0777_ ( .A(\sa22\[2\] ), .B(\sa22\[3\] ), .X(\us22\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0779_ ( .A(\us22\/_0358_ ), .X(\us22\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_0780_ ( .A1(\us22\/_0325_ ), .A2(\us22\/_0347_ ), .B1(\us22\/_0380_ ), .C1(\us22\/_0304_ ), .Y(\us22\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us22/_0781_ ( .A_N(\us22\/_0238_ ), .B(\us22\/_0314_ ), .C(\us22\/_0391_ ), .X(\us22\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us22/_0782_ ( .A(\sa22\[3\] ), .B_N(\sa22\[2\] ), .Y(\us22\/_0412_ ) );
sky130_fd_sc_hd__buf_2 \us22/_0783_ ( .A(\us22\/_0412_ ), .X(\us22\/_0423_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0784_ ( .A(\us22\/_0423_ ), .B(\us22\/_0205_ ), .X(\us22\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \us22/_0787_ ( .A(\sa22\[5\] ), .B_N(\sa22\[4\] ), .Y(\us22\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0788_ ( .A(\us22\/_0467_ ), .B(\us22\/_0140_ ), .X(\us22\/_0478_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_0791_ ( .A(\us22\/_0134_ ), .B(\us22\/_0218_ ), .Y(\us22\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_0792_ ( .A(\us22\/_0478_ ), .B(\us22\/_0271_ ), .Y(\us22\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0793_ ( .A(\us22\/_0194_ ), .X(\us22\/_0532_ ) );
sky130_fd_sc_hd__buf_2 \us22/_0794_ ( .A(\us22\/_0249_ ), .X(\us22\/_0543_ ) );
sky130_fd_sc_hd__and2_1 \us22/_0795_ ( .A(\us22\/_0543_ ), .B(\us22\/_0358_ ), .X(\us22\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0797_ ( .A(\us22\/_0554_ ), .X(\us22\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us22/_0798_ ( .A(\us22\/_0216_ ), .B(\us22\/_0358_ ), .X(\us22\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0800_ ( .A(\us22\/_0586_ ), .X(\us22\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_0801_ ( .A1(\us22\/_0532_ ), .A2(\us22\/_0575_ ), .A3(\us22\/_0608_ ), .B1(\us22\/_0218_ ), .Y(\us22\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us22/_0802_ ( .A(\us22\/_0401_ ), .B(\us22\/_0510_ ), .C(\us22\/_0521_ ), .D(\us22\/_0619_ ), .X(\us22\/_0629_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0803_ ( .A(\us22\/_0358_ ), .B(\sa22\[1\] ), .X(\us22\/_0640_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0804_ ( .A(\us22\/_0640_ ), .X(\us22\/_0651_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0805_ ( .A(\us22\/_0205_ ), .B(\us22\/_0260_ ), .X(\us22\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0806_ ( .A(\us22\/_0662_ ), .X(\us22\/_0672_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0807_ ( .A(\us22\/_0672_ ), .X(\us22\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us22/_0808_ ( .A(\sa22\[6\] ), .B_N(\sa22\[7\] ), .Y(\us22\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \us22/_0809_ ( .A(\us22\/_0467_ ), .B(\us22\/_0694_ ), .X(\us22\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0811_ ( .A(\us22\/_0705_ ), .X(\us22\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_0812_ ( .A1(\us22\/_0651_ ), .A2(\us22\/_0293_ ), .A3(\us22\/_0683_ ), .B1(\us22\/_0727_ ), .Y(\us22\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_0813_ ( .A(\sa22\[1\] ), .B(\sa22\[0\] ), .Y(\us22\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0814_ ( .A(\us22\/_0730_ ), .B(\us22\/_0260_ ), .X(\us22\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0815_ ( .A(\us22\/_0731_ ), .X(\us22\/_0732_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0816_ ( .A(\us22\/_0732_ ), .X(\us22\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0817_ ( .A(\sa22\[0\] ), .X(\us22\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us22/_0818_ ( .A1(\us22\/_0325_ ), .A2(\us22\/_0734_ ), .B1(\us22\/_0423_ ), .X(\us22\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0819_ ( .A(\us22\/_0694_ ), .B(\us22\/_0151_ ), .X(\us22\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0821_ ( .A(\us22\/_0736_ ), .X(\us22\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0822_ ( .A(\us22\/_0738_ ), .X(\us22\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_0823_ ( .A1(\us22\/_0733_ ), .A2(\us22\/_0735_ ), .A3(\us22\/_0293_ ), .B1(\us22\/_0739_ ), .Y(\us22\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us22/_0824_ ( .A(\us22\/_0730_ ), .B_N(\us22\/_0358_ ), .Y(\us22\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_0825_ ( .A(\us22\/_0741_ ), .B(\us22\/_0739_ ), .Y(\us22\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_0827_ ( .A1(\us22\/_0118_ ), .A2(\us22\/_0216_ ), .B1(\us22\/_0532_ ), .C1(\us22\/_0739_ ), .Y(\us22\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us22/_0828_ ( .A(\us22\/_0729_ ), .B(\us22\/_0740_ ), .C(\us22\/_0742_ ), .D(\us22\/_0744_ ), .X(\us22\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0829_ ( .A(\us22\/_0423_ ), .B(\us22\/_0730_ ), .X(\us22\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0830_ ( .A(\us22\/_0746_ ), .X(\us22\/_0747_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0831_ ( .A(\us22\/_0747_ ), .X(\us22\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us22/_0832_ ( .A(\sa22\[4\] ), .B_N(\sa22\[5\] ), .Y(\us22\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0833_ ( .A(\us22\/_0749_ ), .B(\us22\/_0694_ ), .X(\us22\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0835_ ( .A(\us22\/_0750_ ), .X(\us22\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0836_ ( .A(\us22\/_0752_ ), .X(\us22\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0837_ ( .A(\us22\/_0118_ ), .B(\us22\/_0358_ ), .X(\us22\/_0017_ ) );
sky130_fd_sc_hd__buf_2 \us22/_0838_ ( .A(\us22\/_0017_ ), .X(\us22\/_0018_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0839_ ( .A(\us22\/_0752_ ), .B(\us22\/_0018_ ), .X(\us22\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0840_ ( .A(\us22\/_0358_ ), .B(\us22\/_0325_ ), .X(\us22\/_0020_ ) );
sky130_fd_sc_hd__buf_2 \us22/_0841_ ( .A(\us22\/_0020_ ), .X(\us22\/_0021_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0842_ ( .A(\us22\/_0096_ ), .B(\us22\/_0205_ ), .X(\us22\/_0022_ ) );
sky130_fd_sc_hd__buf_2 \us22/_0843_ ( .A(\us22\/_0022_ ), .X(\us22\/_0023_ ) );
sky130_fd_sc_hd__o21a_1 \us22/_0844_ ( .A1(\us22\/_0021_ ), .A2(\us22\/_0023_ ), .B1(\us22\/_0752_ ), .X(\us22\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_0845_ ( .A1(\us22\/_0748_ ), .A2(\us22\/_0016_ ), .B1(\us22\/_0019_ ), .C1(\us22\/_0024_ ), .Y(\us22\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \us22/_0846_ ( .A(\sa22\[4\] ), .B(\sa22\[5\] ), .X(\us22\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0847_ ( .A(\us22\/_0694_ ), .B(\us22\/_0026_ ), .X(\us22\/_0027_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0850_ ( .A(\us22\/_0358_ ), .B(\us22\/_0730_ ), .X(\us22\/_0030_ ) );
sky130_fd_sc_hd__buf_2 \us22/_0852_ ( .A(\us22\/_0030_ ), .X(\us22\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_0853_ ( .A(\us22\/_0247_ ), .B(\us22\/_0032_ ), .Y(\us22\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_0854_ ( .A(\us22\/_0247_ ), .B(\us22\/_0735_ ), .Y(\us22\/_0034_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0855_ ( .A(\us22\/_0118_ ), .B(\us22\/_0260_ ), .X(\us22\/_0035_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0856_ ( .A(\us22\/_0035_ ), .X(\us22\/_0036_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0857_ ( .A(\us22\/_0027_ ), .B(\us22\/_0036_ ), .X(\us22\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0858_ ( .A(\us22\/_0260_ ), .X(\us22\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_0859_ ( .A(\us22\/_0038_ ), .B(\us22\/_0347_ ), .Y(\us22\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us22/_0860_ ( .A_N(\us22\/_0039_ ), .B(\us22\/_0027_ ), .X(\us22\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_0861_ ( .A(\us22\/_0037_ ), .B(\us22\/_0040_ ), .Y(\us22\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us22/_0862_ ( .A(\us22\/_0025_ ), .B(\us22\/_0033_ ), .C(\us22\/_0034_ ), .D(\us22\/_0041_ ), .X(\us22\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0863_ ( .A(\us22\/_0749_ ), .B(\us22\/_0140_ ), .X(\us22\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us22/_0865_ ( .A(\sa22\[0\] ), .B(\sa22\[2\] ), .C(\sa22\[3\] ), .X(\us22\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0866_ ( .A(\us22\/_0043_ ), .B(\us22\/_0045_ ), .X(\us22\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0867_ ( .A(\us22\/_0096_ ), .B(\us22\/_0543_ ), .X(\us22\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0869_ ( .A(\us22\/_0047_ ), .B(\us22\/_0043_ ), .X(\us22\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0870_ ( .A(\us22\/_0730_ ), .X(\us22\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0871_ ( .A(\us22\/_0043_ ), .X(\us22\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_0872_ ( .A1(\us22\/_0118_ ), .A2(\us22\/_0050_ ), .B1(\us22\/_0194_ ), .C1(\us22\/_0051_ ), .Y(\us22\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us22/_0873_ ( .A(\us22\/_0046_ ), .B(\us22\/_0049_ ), .C_N(\us22\/_0052_ ), .Y(\us22\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0874_ ( .A(\us22\/_0026_ ), .B(\us22\/_0140_ ), .X(\us22\/_0054_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0876_ ( .A(\us22\/_0054_ ), .X(\us22\/_0056_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_0877_ ( .A1(\us22\/_0532_ ), .A2(\us22\/_0575_ ), .B1(\us22\/_0056_ ), .Y(\us22\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0878_ ( .A(\us22\/_0423_ ), .B(\us22\/_0325_ ), .X(\us22\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0880_ ( .A(\us22\/_0051_ ), .X(\us22\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_0881_ ( .A1(\us22\/_0732_ ), .A2(\us22\/_0036_ ), .A3(\us22\/_0058_ ), .B1(\us22\/_0060_ ), .Y(\us22\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0882_ ( .A(\us22\/_0260_ ), .B(\sa22\[1\] ), .X(\us22\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0884_ ( .A(\us22\/_0062_ ), .X(\us22\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_0885_ ( .A1(\us22\/_0064_ ), .A2(\us22\/_0748_ ), .A3(\us22\/_0683_ ), .B1(\us22\/_0056_ ), .Y(\us22\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us22/_0886_ ( .A(\us22\/_0053_ ), .B(\us22\/_0057_ ), .C(\us22\/_0061_ ), .D(\us22\/_0065_ ), .X(\us22\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us22/_0887_ ( .A(\us22\/_0629_ ), .B(\us22\/_0745_ ), .C(\us22\/_0042_ ), .D(\us22\/_0066_ ), .X(\us22\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us22/_0889_ ( .A(\sa22\[7\] ), .B_N(\sa22\[6\] ), .Y(\us22\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0890_ ( .A(\us22\/_0069_ ), .B(\us22\/_0151_ ), .X(\us22\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0892_ ( .A(\us22\/_0070_ ), .X(\us22\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_0893_ ( .A1(\us22\/_0129_ ), .A2(\us22\/_0586_ ), .B1(\us22\/_0072_ ), .Y(\us22\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_0894_ ( .A1(\us22\/_0380_ ), .A2(\us22\/_0347_ ), .B1(\us22\/_0194_ ), .B2(\us22\/_0216_ ), .Y(\us22\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us22/_0895_ ( .A(\us22\/_0074_ ), .B_N(\us22\/_0070_ ), .Y(\us22\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us22/_0896_ ( .A(\us22\/_0073_ ), .SLEEP(\us22\/_0075_ ), .X(\us22\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us22/_0897_ ( .A(\us22\/_0467_ ), .B(\us22\/_0069_ ), .X(\us22\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0898_ ( .A(\us22\/_0077_ ), .X(\us22\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0899_ ( .A(\us22\/_0412_ ), .B(\us22\/_0118_ ), .X(\us22\/_0079_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0900_ ( .A(\us22\/_0079_ ), .X(\us22\/_0080_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0901_ ( .A(\us22\/_0078_ ), .B(\us22\/_0080_ ), .X(\us22\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0902_ ( .A(\us22\/_0412_ ), .B(\us22\/_0249_ ), .X(\us22\/_0082_ ) );
sky130_fd_sc_hd__buf_2 \us22/_0904_ ( .A(\us22\/_0082_ ), .X(\us22\/_0084_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0905_ ( .A(\us22\/_0084_ ), .B(\us22\/_0078_ ), .X(\us22\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us22/_0906_ ( .A1(\sa22\[0\] ), .A2(\us22\/_0325_ ), .B1(\us22\/_0260_ ), .Y(\us22\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us22/_0907_ ( .A_N(\us22\/_0086_ ), .B(\us22\/_0078_ ), .X(\us22\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us22/_0908_ ( .A(\us22\/_0081_ ), .B(\us22\/_0085_ ), .C(\us22\/_0087_ ), .Y(\us22\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0909_ ( .A(\us22\/_0072_ ), .X(\us22\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_0910_ ( .A1(\us22\/_0733_ ), .A2(\us22\/_0748_ ), .A3(\us22\/_0683_ ), .B1(\us22\/_0089_ ), .Y(\us22\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0911_ ( .A(\us22\/_0129_ ), .X(\us22\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0912_ ( .A(\us22\/_0018_ ), .X(\us22\/_0092_ ) );
sky130_fd_sc_hd__buf_2 \us22/_0913_ ( .A(\us22\/_0023_ ), .X(\us22\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0914_ ( .A(\us22\/_0078_ ), .X(\us22\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_0915_ ( .A1(\us22\/_0091_ ), .A2(\us22\/_0092_ ), .A3(\us22\/_0093_ ), .B1(\us22\/_0094_ ), .Y(\us22\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us22/_0916_ ( .A(\us22\/_0076_ ), .B(\us22\/_0088_ ), .C(\us22\/_0090_ ), .D(\us22\/_0095_ ), .X(\us22\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us22/_0917_ ( .A(\us22\/_0069_ ), .B(\us22\/_0026_ ), .X(\us22\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \us22/_0918_ ( .A(\us22\/_0098_ ), .X(\us22\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0919_ ( .A(\us22\/_0434_ ), .B(\us22\/_0099_ ), .X(\us22\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0920_ ( .A(\us22\/_0080_ ), .B(\us22\/_0098_ ), .X(\us22\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0921_ ( .A(\us22\/_0325_ ), .X(\us22\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_0922_ ( .A1(\us22\/_0102_ ), .A2(\us22\/_0734_ ), .B1(\us22\/_0038_ ), .C1(\us22\/_0099_ ), .Y(\us22\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us22/_0923_ ( .A(\us22\/_0100_ ), .B(\us22\/_0101_ ), .C_N(\us22\/_0103_ ), .Y(\us22\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_0924_ ( .A1(\us22\/_0554_ ), .A2(\us22\/_0586_ ), .B1(\us22\/_0099_ ), .Y(\us22\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_0925_ ( .A(\us22\/_0129_ ), .B(\us22\/_0099_ ), .Y(\us22\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0926_ ( .A(\us22\/_0105_ ), .B(\us22\/_0106_ ), .X(\us22\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0927_ ( .A(\us22\/_0423_ ), .X(\us22\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us22/_0928_ ( .A(\us22\/_0260_ ), .B(\sa22\[0\] ), .X(\us22\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0929_ ( .A(\us22\/_0069_ ), .B(\us22\/_0749_ ), .X(\us22\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0931_ ( .A(\us22\/_0111_ ), .X(\us22\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0932_ ( .A(\us22\/_0113_ ), .X(\us22\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_0933_ ( .A1(\us22\/_0109_ ), .A2(\us22\/_0110_ ), .B1(\us22\/_0114_ ), .Y(\us22\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us22/_0934_ ( .A(\us22\/_0023_ ), .Y(\us22\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us22/_0935_ ( .A(\us22\/_0554_ ), .Y(\us22\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us22/_0936_ ( .A1(\us22\/_0050_ ), .A2(\us22\/_0118_ ), .B1(\us22\/_0194_ ), .Y(\us22\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us22/_0937_ ( .A(\us22\/_0113_ ), .Y(\us22\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us22/_0938_ ( .A1(\us22\/_0116_ ), .A2(\us22\/_0117_ ), .A3(\us22\/_0119_ ), .B1(\us22\/_0120_ ), .X(\us22\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us22/_0939_ ( .A(\us22\/_0104_ ), .B(\us22\/_0108_ ), .C(\us22\/_0115_ ), .D(\us22\/_0121_ ), .X(\us22\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_0940_ ( .A(\sa22\[7\] ), .B(\sa22\[6\] ), .Y(\us22\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0941_ ( .A(\us22\/_0749_ ), .B(\us22\/_0123_ ), .X(\us22\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0943_ ( .A(\us22\/_0082_ ), .B(\us22\/_0124_ ), .X(\us22\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_0944_ ( .A(\us22\/_0271_ ), .B(\us22\/_0124_ ), .Y(\us22\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0945_ ( .A(\us22\/_0124_ ), .X(\us22\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0946_ ( .A(\us22\/_0260_ ), .B(\us22\/_0325_ ), .X(\us22\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_0948_ ( .A(\us22\/_0128_ ), .B(\us22\/_0130_ ), .Y(\us22\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_0949_ ( .A(\us22\/_0127_ ), .B(\us22\/_0132_ ), .Y(\us22\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us22/_0950_ ( .A(\us22\/_0434_ ), .X(\us22\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_0951_ ( .A(\us22\/_0134_ ), .B(\us22\/_0128_ ), .Y(\us22\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us22/_0952_ ( .A(\us22\/_0126_ ), .B(\us22\/_0133_ ), .C_N(\us22\/_0135_ ), .Y(\us22\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us22/_0953_ ( .A(\us22\/_0026_ ), .B(\us22\/_0123_ ), .X(\us22\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0955_ ( .A(\us22\/_0137_ ), .X(\us22\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_0956_ ( .A1(\us22\/_0110_ ), .A2(\us22\/_0293_ ), .A3(\us22\/_0084_ ), .B1(\us22\/_0139_ ), .Y(\us22\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0957_ ( .A(\us22\/_0096_ ), .B(\us22\/_0730_ ), .X(\us22\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0959_ ( .A(\us22\/_0142_ ), .X(\us22\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_0960_ ( .A1(\us22\/_0021_ ), .A2(\us22\/_0144_ ), .A3(\us22\/_0018_ ), .B1(\us22\/_0139_ ), .Y(\us22\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \us22/_0961_ ( .A(\sa22\[2\] ), .B(\us22\/_0050_ ), .C_N(\sa22\[3\] ), .Y(\us22\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0962_ ( .A(\us22\/_0128_ ), .X(\us22\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_0963_ ( .A1(\us22\/_0146_ ), .A2(\us22\/_0032_ ), .A3(\us22\/_0651_ ), .B1(\us22\/_0147_ ), .Y(\us22\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us22/_0964_ ( .A(\us22\/_0136_ ), .B(\us22\/_0141_ ), .C(\us22\/_0145_ ), .D(\us22\/_0148_ ), .X(\us22\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0965_ ( .A(\us22\/_0123_ ), .B(\us22\/_0151_ ), .X(\us22\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0967_ ( .A(\us22\/_0150_ ), .X(\us22\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \us22/_0968_ ( .A(\us22\/_0150_ ), .B(\us22\/_0062_ ), .X(\us22\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_0969_ ( .A(\us22\/_0080_ ), .B(\us22\/_0150_ ), .Y(\us22\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us22/_0970_ ( .A(\us22\/_0150_ ), .B(\us22\/_0423_ ), .C(\us22\/_0543_ ), .Y(\us22\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_0971_ ( .A(\us22\/_0155_ ), .B(\us22\/_0156_ ), .Y(\us22\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_0972_ ( .A1(\us22\/_0153_ ), .A2(\us22\/_0134_ ), .B1(\us22\/_0154_ ), .C1(\us22\/_0157_ ), .Y(\us22\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0973_ ( .A(\us22\/_0467_ ), .B(\us22\/_0123_ ), .X(\us22\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_0975_ ( .A(\us22\/_0159_ ), .X(\us22\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us22/_0976_ ( .A_N(\us22\/_0119_ ), .B(\us22\/_0161_ ), .X(\us22\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us22/_0977_ ( .A(\us22\/_0163_ ), .Y(\us22\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_0978_ ( .A1(\us22\/_0146_ ), .A2(\us22\/_0575_ ), .A3(\us22\/_0608_ ), .B1(\us22\/_0153_ ), .Y(\us22\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_0979_ ( .A1(\us22\/_0062_ ), .A2(\us22\/_0084_ ), .A3(\us22\/_0134_ ), .B1(\us22\/_0161_ ), .Y(\us22\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us22/_0980_ ( .A(\us22\/_0158_ ), .B(\us22\/_0164_ ), .C(\us22\/_0165_ ), .D(\us22\/_0166_ ), .X(\us22\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us22/_0981_ ( .A(\us22\/_0097_ ), .B(\us22\/_0122_ ), .C(\us22\/_0149_ ), .D(\us22\/_0167_ ), .X(\us22\/_0168_ ) );
sky130_fd_sc_hd__and2_1 \us22/_0982_ ( .A(\us22\/_0672_ ), .B(\us22\/_0150_ ), .X(\us22\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_0983_ ( .A(\us22\/_0154_ ), .B(\us22\/_0169_ ), .Y(\us22\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us22/_0984_ ( .A(\us22\/_0123_ ), .B(\us22\/_0151_ ), .C(\us22\/_0038_ ), .X(\us22\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0985_ ( .A(\us22\/_0170_ ), .B(\us22\/_0171_ ), .X(\us22\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \us22/_0986_ ( .A(\us22\/_0172_ ), .Y(\us22\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \us22/_0987_ ( .A(\us22\/_0067_ ), .B(\us22\/_0168_ ), .C(\us22\/_0174_ ), .Y(\us22\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us22/_0988_ ( .A(\sa22\[1\] ), .B(\sa22\[0\] ), .Y(\us22\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us22/_0989_ ( .A(\us22\/_0175_ ), .B(\us22\/_0358_ ), .X(\us22\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0990_ ( .A(\us22\/_0176_ ), .B(\us22\/_0478_ ), .X(\us22\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_0991_ ( .A(\us22\/_0084_ ), .B(\us22\/_0113_ ), .Y(\us22\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0992_ ( .A(\us22\/_0111_ ), .B(\us22\/_0062_ ), .X(\us22\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0993_ ( .A(\us22\/_0111_ ), .B(\us22\/_0672_ ), .X(\us22\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_0994_ ( .A(\us22\/_0179_ ), .B(\us22\/_0180_ ), .Y(\us22\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0995_ ( .A(\us22\/_0054_ ), .B(\us22\/_0058_ ), .X(\us22\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us22/_0996_ ( .A(\us22\/_0182_ ), .Y(\us22\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us22/_0997_ ( .A_N(\us22\/_0177_ ), .B(\us22\/_0178_ ), .C(\us22\/_0181_ ), .D(\us22\/_0184_ ), .X(\us22\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0998_ ( .A(\us22\/_0098_ ), .B(\us22\/_0741_ ), .X(\us22\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us22/_0999_ ( .A(\us22\/_0047_ ), .B(\us22\/_0098_ ), .X(\us22\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us22/_1000_ ( .A(\us22\/_0186_ ), .B(\us22\/_0187_ ), .X(\us22\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1001_ ( .A(\us22\/_0188_ ), .Y(\us22\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1002_ ( .A(\us22\/_0738_ ), .B(\us22\/_0735_ ), .X(\us22\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1003_ ( .A(\us22\/_0271_ ), .B(\us22\/_0736_ ), .X(\us22\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_1004_ ( .A(\us22\/_0190_ ), .B(\us22\/_0191_ ), .Y(\us22\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us22/_1005_ ( .A(\us22\/_0096_ ), .B(\us22\/_0325_ ), .X(\us22\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1006_ ( .A1(\us22\/_0193_ ), .A2(\us22\/_0176_ ), .B1(\us22\/_0043_ ), .Y(\us22\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1007_ ( .A(\us22\/_0185_ ), .B(\us22\/_0189_ ), .C(\us22\/_0192_ ), .D(\us22\/_0195_ ), .X(\us22\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us22/_1008_ ( .A_N(\sa22\[3\] ), .B(\us22\/_0734_ ), .C(\sa22\[2\] ), .X(\us22\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1009_ ( .A(\us22\/_0137_ ), .B(\us22\/_0197_ ), .X(\us22\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_1010_ ( .A(\us22\/_0198_ ), .B(\us22\/_0040_ ), .Y(\us22\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1011_ ( .A(\us22\/_0293_ ), .B(\us22\/_0137_ ), .X(\us22\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1012_ ( .A(\us22\/_0200_ ), .Y(\us22\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1013_ ( .A(\us22\/_0137_ ), .B(\us22\/_0110_ ), .Y(\us22\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1014_ ( .A(\us22\/_0139_ ), .B(\us22\/_0021_ ), .Y(\us22\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1015_ ( .A(\us22\/_0199_ ), .B(\us22\/_0201_ ), .C(\us22\/_0202_ ), .D(\us22\/_0203_ ), .X(\us22\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us22/_1016_ ( .A1(\us22\/_0532_ ), .A2(\us22\/_0109_ ), .B1(\us22\/_0102_ ), .C1(\us22\/_0727_ ), .X(\us22\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1017_ ( .A(\us22\/_0023_ ), .B(\us22\/_0078_ ), .Y(\us22\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1018_ ( .A(\us22\/_0078_ ), .B(\us22\/_0142_ ), .Y(\us22\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1019_ ( .A(\us22\/_0207_ ), .B(\us22\/_0208_ ), .Y(\us22\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1020_ ( .A1(\us22\/_0094_ ), .A2(\us22\/_0176_ ), .B1(\us22\/_0206_ ), .C1(\us22\/_0209_ ), .Y(\us22\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1021_ ( .A(\us22\/_0662_ ), .B(\us22\/_0070_ ), .X(\us22\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us22/_1022_ ( .A(\us22\/_0732_ ), .B(\us22\/_0123_ ), .C(\us22\/_0749_ ), .Y(\us22\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us22/_1023_ ( .A(\us22\/_0732_ ), .B(\us22\/_0467_ ), .C(\us22\/_0069_ ), .Y(\us22\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us22/_1024_ ( .A_N(\us22\/_0211_ ), .B(\us22\/_0127_ ), .C(\us22\/_0212_ ), .D(\us22\/_0213_ ), .X(\us22\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1025_ ( .A(\us22\/_0137_ ), .Y(\us22\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1026_ ( .A(\us22\/_0128_ ), .B(\us22\/_0036_ ), .Y(\us22\/_0217_ ) );
sky130_fd_sc_hd__buf_2 \us22/_1027_ ( .A(\us22\/_0478_ ), .X(\us22\/_0218_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1028_ ( .A1(\us22\/_0159_ ), .A2(\us22\/_0747_ ), .B1(\us22\/_0434_ ), .B2(\us22\/_0218_ ), .Y(\us22\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us22/_1029_ ( .A1(\us22\/_0116_ ), .A2(\us22\/_0215_ ), .B1(\us22\/_0217_ ), .C1(\us22\/_0219_ ), .X(\us22\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1030_ ( .A(\us22\/_0113_ ), .B(\us22\/_0746_ ), .X(\us22\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us22/_1031_ ( .A1(\us22\/_0098_ ), .A2(\us22\/_0746_ ), .B1(\us22\/_0434_ ), .B2(\us22\/_0750_ ), .X(\us22\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1032_ ( .A1(\us22\/_0047_ ), .A2(\us22\/_0113_ ), .B1(\us22\/_0221_ ), .C1(\us22\/_0222_ ), .Y(\us22\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us22/_1033_ ( .A1(\us22\/_0129_ ), .A2(\us22\/_0162_ ), .B1(\us22\/_0271_ ), .B2(\us22\/_0705_ ), .X(\us22\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1034_ ( .A1(\us22\/_0093_ ), .A2(\us22\/_0738_ ), .B1(\us22\/_0081_ ), .C1(\us22\/_0224_ ), .Y(\us22\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1035_ ( .A(\us22\/_0214_ ), .B(\us22\/_0220_ ), .C(\us22\/_0223_ ), .D(\us22\/_0225_ ), .X(\us22\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1036_ ( .A(\us22\/_0196_ ), .B(\us22\/_0204_ ), .C(\us22\/_0210_ ), .D(\us22\/_0226_ ), .X(\us22\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1037_ ( .A(\us22\/_0111_ ), .B(\us22\/_0554_ ), .X(\us22\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1038_ ( .A(\us22\/_0229_ ), .Y(\us22\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1039_ ( .A(\us22\/_0111_ ), .B(\us22\/_0129_ ), .Y(\us22\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1040_ ( .A(\us22\/_0018_ ), .B(\us22\/_0738_ ), .Y(\us22\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1041_ ( .A(\us22\/_0030_ ), .B(\us22\/_0304_ ), .Y(\us22\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1042_ ( .A(\us22\/_0230_ ), .B(\us22\/_0231_ ), .C(\us22\/_0232_ ), .D(\us22\/_0233_ ), .X(\us22\/_0234_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1043_ ( .A(\us22\/_0047_ ), .B(\us22\/_0478_ ), .X(\us22\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1044_ ( .A1(\us22\/_0129_ ), .A2(\us22\/_0554_ ), .B1(\us22\/_0137_ ), .Y(\us22\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us22/_1045_ ( .A(\us22\/_0235_ ), .B(\us22\/_0049_ ), .C_N(\us22\/_0236_ ), .Y(\us22\/_0237_ ) );
sky130_fd_sc_hd__and2_1 \us22/_1046_ ( .A(\us22\/_0047_ ), .B(\us22\/_0077_ ), .X(\us22\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1047_ ( .A(\us22\/_0070_ ), .B(\us22\/_0036_ ), .X(\us22\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us22/_1048_ ( .A1(\us22\/_0047_ ), .A2(\us22\/_0736_ ), .B1(\us22\/_0023_ ), .B2(\us22\/_0099_ ), .X(\us22\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us22/_1049_ ( .A(\us22\/_0239_ ), .B(\us22\/_0240_ ), .C(\us22\/_0241_ ), .Y(\us22\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1050_ ( .A(\us22\/_0554_ ), .B(\us22\/_0072_ ), .X(\us22\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us22/_1051_ ( .A1(\us22\/_0142_ ), .A2(\us22\/_0137_ ), .B1(\us22\/_0159_ ), .B2(\us22\/_0082_ ), .X(\us22\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1052_ ( .A1(\us22\/_0608_ ), .A2(\us22\/_0072_ ), .B1(\us22\/_0243_ ), .C1(\us22\/_0244_ ), .Y(\us22\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1053_ ( .A(\us22\/_0234_ ), .B(\us22\/_0237_ ), .C(\us22\/_0242_ ), .D(\us22\/_0245_ ), .X(\us22\/_0246_ ) );
sky130_fd_sc_hd__buf_2 \us22/_1054_ ( .A(\us22\/_0027_ ), .X(\us22\/_0247_ ) );
sky130_fd_sc_hd__o21a_1 \us22/_1055_ ( .A1(\us22\/_0554_ ), .A2(\us22\/_0586_ ), .B1(\us22\/_0247_ ), .X(\us22\/_0248_ ) );
sky130_fd_sc_hd__and2_1 \us22/_1056_ ( .A(\us22\/_0082_ ), .B(\us22\/_0478_ ), .X(\us22\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_1057_ ( .A(\us22\/_0080_ ), .X(\us22\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1058_ ( .A(\us22\/_0251_ ), .B(\us22\/_0478_ ), .X(\us22\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_1059_ ( .A(\us22\/_0250_ ), .B(\us22\/_0252_ ), .Y(\us22\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1060_ ( .A(\us22\/_0016_ ), .B(\us22\/_0064_ ), .Y(\us22\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_1061_ ( .A(\us22\/_0304_ ), .X(\us22\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1062_ ( .A(\us22\/_0255_ ), .B(\us22\/_0651_ ), .Y(\us22\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us22/_1063_ ( .A_N(\us22\/_0248_ ), .B(\us22\/_0253_ ), .C(\us22\/_0254_ ), .D(\us22\/_0256_ ), .X(\us22\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1064_ ( .A(\us22\/_0099_ ), .B(\us22\/_0110_ ), .X(\us22\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us22/_1065_ ( .A1(\us22\/_0161_ ), .A2(\us22\/_0130_ ), .B1(\us22\/_0258_ ), .Y(\us22\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1066_ ( .A(\us22\/_0194_ ), .B(\sa22\[1\] ), .X(\us22\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1068_ ( .A(\us22\/_0261_ ), .B(\us22\/_0153_ ), .Y(\us22\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us22/_1069_ ( .A_N(\us22\/_0154_ ), .B(\us22\/_0259_ ), .C(\us22\/_0263_ ), .X(\us22\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1070_ ( .A(\us22\/_0246_ ), .B(\us22\/_0174_ ), .C(\us22\/_0257_ ), .D(\us22\/_0264_ ), .X(\us22\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us22/_1071_ ( .A1(\us22\/_0261_ ), .A2(\us22\/_0554_ ), .B1(\us22\/_0159_ ), .X(\us22\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1072_ ( .A(\us22\/_0747_ ), .B(\us22\/_0150_ ), .Y(\us22\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1073_ ( .A(\us22\/_0175_ ), .Y(\us22\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us22/_1074_ ( .A(\us22\/_0423_ ), .B(\us22\/_0123_ ), .C(\us22\/_0151_ ), .X(\us22\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1075_ ( .A(\us22\/_0268_ ), .B(\us22\/_0269_ ), .Y(\us22\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us22/_1076_ ( .A_N(\us22\/_0266_ ), .B(\us22\/_0267_ ), .C(\us22\/_0270_ ), .X(\us22\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1077_ ( .A(\us22\/_0554_ ), .B(\us22\/_0150_ ), .X(\us22\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1078_ ( .A(\us22\/_0273_ ), .Y(\us22\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1079_ ( .A1(\us22\/_0734_ ), .A2(\us22\/_0325_ ), .B1(\us22\/_0380_ ), .Y(\us22\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1080_ ( .A(\us22\/_0275_ ), .Y(\us22\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1081_ ( .A(\us22\/_0276_ ), .B(\us22\/_0153_ ), .Y(\us22\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us22/_1082_ ( .A(\us22\/_0272_ ), .B(\us22\/_0274_ ), .C(\us22\/_0277_ ), .X(\us22\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_1083_ ( .A(\us22\/_0036_ ), .X(\us22\/_0279_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1085_ ( .A1(\us22\/_0218_ ), .A2(\us22\/_0279_ ), .B1(\us22\/_0084_ ), .B2(\us22\/_0060_ ), .Y(\us22\/_0281_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1086_ ( .A1(\us22\/_0251_ ), .A2(\us22\/_0434_ ), .B1(\us22\/_0304_ ), .Y(\us22\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1087_ ( .A(\us22\/_0091_ ), .B(\us22\/_0056_ ), .Y(\us22\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1088_ ( .A1(\us22\/_0118_ ), .A2(\us22\/_0050_ ), .B1(\us22\/_0038_ ), .C1(\us22\/_0255_ ), .Y(\us22\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1089_ ( .A(\us22\/_0281_ ), .B(\us22\/_0283_ ), .C(\us22\/_0284_ ), .D(\us22\/_0285_ ), .X(\us22\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1090_ ( .A(\us22\/_0082_ ), .B(\us22\/_0027_ ), .X(\us22\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1091_ ( .A(\us22\/_0129_ ), .B(\us22\/_0027_ ), .X(\us22\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_1092_ ( .A(\us22\/_0287_ ), .B(\us22\/_0288_ ), .Y(\us22\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1093_ ( .A1(\us22\/_0752_ ), .A2(\us22\/_0683_ ), .B1(\us22\/_0093_ ), .B2(\us22\/_0247_ ), .Y(\us22\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1094_ ( .A1(\us22\/_0092_ ), .A2(\us22\/_0575_ ), .B1(\us22\/_0056_ ), .Y(\us22\/_0291_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1096_ ( .A1(\us22\/_0218_ ), .A2(\us22\/_0672_ ), .B1(\us22\/_0084_ ), .B2(\us22\/_0056_ ), .Y(\us22\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1097_ ( .A(\us22\/_0289_ ), .B(\us22\/_0290_ ), .C(\us22\/_0291_ ), .D(\us22\/_0294_ ), .X(\us22\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1098_ ( .A(\us22\/_0750_ ), .B(\us22\/_0193_ ), .X(\us22\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1099_ ( .A(\us22\/_0705_ ), .B(\us22\/_0380_ ), .X(\us22\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1100_ ( .A(\us22\/_0752_ ), .B(\us22\/_0129_ ), .Y(\us22\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us22/_1101_ ( .A(\us22\/_0296_ ), .B(\us22\/_0297_ ), .C_N(\us22\/_0298_ ), .Y(\us22\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1102_ ( .A(\us22\/_0089_ ), .B(\us22\/_0532_ ), .Y(\us22\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1103_ ( .A(\sa22\[2\] ), .Y(\us22\/_0301_ ) );
sky130_fd_sc_hd__nor3_2 \us22/_1104_ ( .A(\us22\/_0301_ ), .B(\sa22\[3\] ), .C(\us22\/_0118_ ), .Y(\us22\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1105_ ( .A(\us22\/_0072_ ), .B(\us22\/_0302_ ), .X(\us22\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1106_ ( .A(\us22\/_0303_ ), .Y(\us22\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1107_ ( .A(\us22\/_0147_ ), .B(\us22\/_0302_ ), .Y(\us22\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1108_ ( .A(\us22\/_0299_ ), .B(\us22\/_0300_ ), .C(\us22\/_0305_ ), .D(\us22\/_0306_ ), .X(\us22\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1109_ ( .A(\us22\/_0278_ ), .B(\us22\/_0286_ ), .C(\us22\/_0295_ ), .D(\us22\/_0307_ ), .X(\us22\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us22/_1110_ ( .A(\us22\/_0228_ ), .B(\us22\/_0265_ ), .C(\us22\/_0308_ ), .Y(\us22\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1111_ ( .A(\us22\/_0235_ ), .Y(\us22\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1112_ ( .A(\us22\/_0478_ ), .B(\us22\/_0640_ ), .X(\us22\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1113_ ( .A(\us22\/_0310_ ), .Y(\us22\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1114_ ( .A(\us22\/_0023_ ), .B(\us22\/_0218_ ), .Y(\us22\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1115_ ( .A(\us22\/_0218_ ), .B(\us22\/_0032_ ), .Y(\us22\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1116_ ( .A(\us22\/_0309_ ), .B(\us22\/_0311_ ), .C(\us22\/_0312_ ), .D(\us22\/_0313_ ), .X(\us22\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1117_ ( .A(\us22\/_0218_ ), .B(\us22\/_0064_ ), .Y(\us22\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1118_ ( .A(\us22\/_0218_ ), .B(\us22\/_0683_ ), .Y(\us22\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1119_ ( .A(\us22\/_0315_ ), .B(\us22\/_0316_ ), .C(\us22\/_0317_ ), .D(\us22\/_0253_ ), .X(\us22\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1120_ ( .A(\us22\/_0047_ ), .B(\us22\/_0304_ ), .Y(\us22\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1121_ ( .A(\us22\/_0586_ ), .B(\us22\/_0162_ ), .Y(\us22\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1122_ ( .A(\us22\/_0319_ ), .B(\us22\/_0320_ ), .Y(\us22\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_1123_ ( .A(\us22\/_0321_ ), .B(\us22\/_0238_ ), .Y(\us22\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1124_ ( .A(\us22\/_0304_ ), .B(\us22\/_0062_ ), .Y(\us22\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_1125_ ( .A(\us22\/_0251_ ), .X(\us22\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1126_ ( .A1(\us22\/_0324_ ), .A2(\us22\/_0084_ ), .B1(\us22\/_0255_ ), .Y(\us22\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1127_ ( .A1(\us22\/_0050_ ), .A2(\us22\/_0216_ ), .B1(\us22\/_0109_ ), .C1(\us22\/_0255_ ), .Y(\us22\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1128_ ( .A(\us22\/_0322_ ), .B(\us22\/_0323_ ), .C(\us22\/_0326_ ), .D(\us22\/_0327_ ), .X(\us22\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1129_ ( .A1(\us22\/_0733_ ), .A2(\us22\/_0279_ ), .A3(\us22\/_0058_ ), .B1(\us22\/_0056_ ), .Y(\us22\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_1130_ ( .A(\us22\/_0047_ ), .X(\us22\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1131_ ( .A(\us22\/_0330_ ), .B(\us22\/_0056_ ), .Y(\us22\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1132_ ( .A(\us22\/_0054_ ), .B(\us22\/_0045_ ), .Y(\us22\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1133_ ( .A(\us22\/_0329_ ), .B(\us22\/_0331_ ), .C(\us22\/_0284_ ), .D(\us22\/_0332_ ), .X(\us22\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us22/_1134_ ( .A1(\us22\/_0543_ ), .A2(\us22\/_0216_ ), .B1(\us22\/_0532_ ), .C1(\us22\/_0060_ ), .X(\us22\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1135_ ( .A(\us22\/_0084_ ), .B(\us22\/_0060_ ), .Y(\us22\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1136_ ( .A(\us22\/_0324_ ), .B(\us22\/_0060_ ), .Y(\us22\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1137_ ( .A(\us22\/_0335_ ), .B(\us22\/_0337_ ), .Y(\us22\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1138_ ( .A1(\us22\/_0276_ ), .A2(\us22\/_0060_ ), .B1(\us22\/_0334_ ), .C1(\us22\/_0338_ ), .Y(\us22\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1139_ ( .A(\us22\/_0318_ ), .B(\us22\/_0328_ ), .C(\us22\/_0333_ ), .D(\us22\/_0339_ ), .X(\us22\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us22/_1140_ ( .A1(\us22\/_0747_ ), .A2(\us22\/_0134_ ), .B1(\us22\/_0128_ ), .X(\us22\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us22/_1141_ ( .A_N(\us22\/_0086_ ), .B(\us22\/_0128_ ), .X(\us22\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1142_ ( .A(\us22\/_0080_ ), .B(\us22\/_0124_ ), .X(\us22\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_1143_ ( .A(\us22\/_0126_ ), .B(\us22\/_0343_ ), .Y(\us22\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us22/_1144_ ( .A(\us22\/_0341_ ), .B(\us22\/_0342_ ), .C_N(\us22\/_0344_ ), .Y(\us22\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1146_ ( .A1(\us22\/_0193_ ), .A2(\us22\/_0092_ ), .A3(\us22\/_0330_ ), .B1(\us22\/_0147_ ), .Y(\us22\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1147_ ( .A1(\us22\/_0130_ ), .A2(\us22\/_0084_ ), .A3(\us22\/_0134_ ), .B1(\us22\/_0139_ ), .Y(\us22\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1148_ ( .A1(\us22\/_0144_ ), .A2(\us22\/_0608_ ), .A3(\us22\/_0092_ ), .B1(\us22\/_0139_ ), .Y(\us22\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1149_ ( .A(\us22\/_0345_ ), .B(\us22\/_0348_ ), .C(\us22\/_0349_ ), .D(\us22\/_0350_ ), .X(\us22\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us22/_1150_ ( .A(\us22\/_0150_ ), .B(\us22\/_0194_ ), .C(\us22\/_0543_ ), .X(\us22\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us22/_1151_ ( .A(\us22\/_0277_ ), .SLEEP(\us22\/_0352_ ), .X(\us22\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us22/_1152_ ( .A1(\us22\/_0268_ ), .A2(\us22\/_0171_ ), .B1(\us22\/_0157_ ), .Y(\us22\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us22/_1153_ ( .A(\us22\/_0161_ ), .X(\us22\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1154_ ( .A1(\us22\/_0279_ ), .A2(\us22\/_0084_ ), .B1(\us22\/_0355_ ), .Y(\us22\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1155_ ( .A1(\us22\/_0021_ ), .A2(\us22\/_0193_ ), .A3(\us22\/_0091_ ), .B1(\us22\/_0355_ ), .Y(\us22\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1156_ ( .A(\us22\/_0353_ ), .B(\us22\/_0354_ ), .C(\us22\/_0356_ ), .D(\us22\/_0357_ ), .X(\us22\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1157_ ( .A(\us22\/_0111_ ), .B(\us22\/_0586_ ), .X(\us22\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1158_ ( .A(\us22\/_0360_ ), .Y(\us22\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us22/_1159_ ( .A1(\us22\/_0119_ ), .A2(\us22\/_0120_ ), .B1(\us22\/_0230_ ), .C1(\us22\/_0361_ ), .X(\us22\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1160_ ( .A1(\us22\/_0672_ ), .A2(\us22\/_0251_ ), .A3(\us22\/_0134_ ), .B1(\us22\/_0114_ ), .Y(\us22\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1162_ ( .A1(\us22\/_0036_ ), .A2(\us22\/_0251_ ), .A3(\us22\/_0134_ ), .B1(\us22\/_0099_ ), .Y(\us22\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1163_ ( .A1(\us22\/_0193_ ), .A2(\us22\/_0608_ ), .B1(\us22\/_0099_ ), .Y(\us22\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1164_ ( .A(\us22\/_0362_ ), .B(\us22\/_0363_ ), .C(\us22\/_0365_ ), .D(\us22\/_0366_ ), .X(\us22\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1165_ ( .A1(\us22\/_0575_ ), .A2(\us22\/_0092_ ), .A3(\us22\/_0330_ ), .B1(\us22\/_0089_ ), .Y(\us22\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1166_ ( .A1(\us22\/_0586_ ), .A2(\us22\/_0018_ ), .A3(\us22\/_0330_ ), .B1(\us22\/_0094_ ), .Y(\us22\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \us22/_1167_ ( .A1(\us22\/_0293_ ), .A2(\us22\/_0134_ ), .B1(\us22\/_0089_ ), .Y(\us22\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1168_ ( .A1(\us22\/_0279_ ), .A2(\us22\/_0134_ ), .B1(\us22\/_0094_ ), .Y(\us22\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1169_ ( .A(\us22\/_0368_ ), .B(\us22\/_0370_ ), .C(\us22\/_0371_ ), .D(\us22\/_0372_ ), .X(\us22\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1170_ ( .A(\us22\/_0351_ ), .B(\us22\/_0359_ ), .C(\us22\/_0367_ ), .D(\us22\/_0373_ ), .X(\us22\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1171_ ( .A1(\us22\/_0102_ ), .A2(\us22\/_0347_ ), .B1(\us22\/_0109_ ), .C1(\us22\/_0247_ ), .Y(\us22\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1172_ ( .A1(\us22\/_0102_ ), .A2(\us22\/_0347_ ), .B1(\us22\/_0532_ ), .C1(\us22\/_0247_ ), .Y(\us22\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1173_ ( .A1(\us22\/_0050_ ), .A2(\us22\/_0543_ ), .B1(\us22\/_0380_ ), .C1(\us22\/_0247_ ), .Y(\us22\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1174_ ( .A(\us22\/_0041_ ), .B(\us22\/_0375_ ), .C(\us22\/_0376_ ), .D(\us22\/_0377_ ), .X(\us22\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1175_ ( .A(\us22\/_0047_ ), .B(\us22\/_0750_ ), .X(\us22\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1176_ ( .A(\us22\/_0379_ ), .Y(\us22\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1177_ ( .A(\us22\/_0016_ ), .B(\us22\/_0608_ ), .Y(\us22\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1178_ ( .A(\us22\/_0752_ ), .B(\us22\/_0554_ ), .Y(\us22\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1179_ ( .A1(\sa22\[1\] ), .A2(\us22\/_0734_ ), .B1(\us22\/_0109_ ), .C1(\us22\/_0016_ ), .Y(\us22\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1180_ ( .A(\us22\/_0381_ ), .B(\us22\/_0382_ ), .C(\us22\/_0383_ ), .D(\us22\/_0384_ ), .X(\us22\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us22/_1181_ ( .A(\us22\/_0086_ ), .B_N(\us22\/_0736_ ), .X(\us22\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1182_ ( .A1(\us22\/_0748_ ), .A2(\us22\/_0134_ ), .B1(\us22\/_0739_ ), .Y(\us22\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1183_ ( .A1(\us22\/_0118_ ), .A2(\us22\/_0543_ ), .B1(\us22\/_0109_ ), .C1(\us22\/_0739_ ), .Y(\us22\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1184_ ( .A1(\us22\/_0102_ ), .A2(\us22\/_0301_ ), .B1(\sa22\[3\] ), .C1(\us22\/_0739_ ), .Y(\us22\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1185_ ( .A(\us22\/_0386_ ), .B(\us22\/_0387_ ), .C(\us22\/_0388_ ), .D(\us22\/_0389_ ), .X(\us22\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1186_ ( .A(\us22\/_0021_ ), .Y(\us22\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1187_ ( .A(\us22\/_0727_ ), .Y(\us22\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1188_ ( .A(\us22\/_0727_ ), .B(\us22\/_0064_ ), .Y(\us22\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1189_ ( .A1(\us22\/_0102_ ), .A2(\us22\/_0734_ ), .B1(\us22\/_0532_ ), .C1(\us22\/_0727_ ), .Y(\us22\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us22/_1190_ ( .A1(\us22\/_0392_ ), .A2(\us22\/_0393_ ), .B1(\us22\/_0394_ ), .C1(\us22\/_0395_ ), .X(\us22\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1191_ ( .A(\us22\/_0378_ ), .B(\us22\/_0385_ ), .C(\us22\/_0390_ ), .D(\us22\/_0396_ ), .X(\us22\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us22/_1192_ ( .A(\us22\/_0340_ ), .B(\us22\/_0374_ ), .C(\us22\/_0397_ ), .Y(\us22\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1193_ ( .A(\us22\/_0077_ ), .B(\us22\/_0129_ ), .X(\us22\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_1194_ ( .A(\us22\/_0398_ ), .B(\us22\/_0239_ ), .Y(\us22\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1195_ ( .A(\us22\/_0023_ ), .B(\us22\/_0111_ ), .X(\us22\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us22/_1196_ ( .A_N(\us22\/_0400_ ), .B(\us22\/_0231_ ), .Y(\us22\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us22/_1197_ ( .A(\us22\/_0399_ ), .SLEEP(\us22\/_0402_ ), .X(\us22\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_1198_ ( .A(\us22\/_0747_ ), .B(\us22\/_0251_ ), .Y(\us22\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us22/_1199_ ( .A_N(\us22\/_0404_ ), .B(\us22\/_0752_ ), .Y(\us22\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us22/_1200_ ( .A(\us22\/_0467_ ), .B(\us22\/_0194_ ), .C(\us22\/_0694_ ), .X(\us22\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us22/_1201_ ( .A_N(\us22\/_0175_ ), .B(\us22\/_0406_ ), .X(\us22\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1202_ ( .A(\us22\/_0407_ ), .Y(\us22\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1203_ ( .A1(\us22\/_0094_ ), .A2(\us22\/_0197_ ), .B1(\us22\/_0114_ ), .B2(\us22\/_0651_ ), .Y(\us22\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1204_ ( .A(\us22\/_0403_ ), .B(\us22\/_0405_ ), .C(\us22\/_0408_ ), .D(\us22\/_0409_ ), .X(\us22\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1205_ ( .A(\us22\/_0030_ ), .B(\us22\/_0150_ ), .Y(\us22\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us22/_1206_ ( .A_N(\us22\/_0169_ ), .B(\us22\/_0289_ ), .C(\us22\/_0411_ ), .X(\us22\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us22/_1207_ ( .A1(\us22\/_0467_ ), .A2(\us22\/_0151_ ), .B1(\us22\/_0140_ ), .C1(\us22\/_0129_ ), .X(\us22\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1208_ ( .A1(\us22\/_0608_ ), .A2(\us22\/_0099_ ), .B1(\us22\/_0037_ ), .C1(\us22\/_0414_ ), .Y(\us22\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1209_ ( .A(\us22\/_0738_ ), .Y(\us22\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1210_ ( .A(\us22\/_0586_ ), .B(\us22\/_0736_ ), .Y(\us22\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1211_ ( .A1(\us22\/_0194_ ), .A2(\us22\/_0038_ ), .B1(\us22\/_0118_ ), .C1(\us22\/_0153_ ), .Y(\us22\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us22/_1212_ ( .A1(\us22\/_0416_ ), .A2(\us22\/_0117_ ), .B1(\us22\/_0417_ ), .C1(\us22\/_0418_ ), .X(\us22\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1213_ ( .A(\us22\/_0077_ ), .B(\us22\/_0035_ ), .X(\us22\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1214_ ( .A(\us22\/_0672_ ), .B(\us22\/_0124_ ), .Y(\us22\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1215_ ( .A(\us22\/_0030_ ), .B(\us22\/_0137_ ), .Y(\us22\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1216_ ( .A(\us22\/_0072_ ), .B(\us22\/_0732_ ), .Y(\us22\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us22/_1217_ ( .A_N(\us22\/_0420_ ), .B(\us22\/_0421_ ), .C(\us22\/_0422_ ), .D(\us22\/_0424_ ), .X(\us22\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1218_ ( .A(\us22\/_0413_ ), .B(\us22\/_0415_ ), .C(\us22\/_0419_ ), .D(\us22\/_0425_ ), .X(\us22\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us22/_1219_ ( .A(\us22\/_0355_ ), .B(\us22\/_0102_ ), .C(\us22\/_0109_ ), .Y(\us22\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1220_ ( .A(\us22\/_0077_ ), .B(\us22\/_0018_ ), .X(\us22\/_0428_ ) );
sky130_fd_sc_hd__and2_1 \us22/_1221_ ( .A(\us22\/_0077_ ), .B(\us22\/_0554_ ), .X(\us22\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us22/_1222_ ( .A1(\us22\/_0050_ ), .A2(\us22\/_0216_ ), .B1(\us22\/_0380_ ), .C1(\us22\/_0078_ ), .X(\us22\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us22/_1223_ ( .A(\us22\/_0428_ ), .B(\us22\/_0429_ ), .C(\us22\/_0430_ ), .Y(\us22\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us22/_1224_ ( .A_N(\us22\/_0209_ ), .B(\us22\/_0431_ ), .X(\us22\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us22/_1225_ ( .A1(\us22\/_0215_ ), .A2(\us22\/_0404_ ), .B1(\us22\/_0427_ ), .C1(\us22\/_0432_ ), .X(\us22\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1226_ ( .A(\us22\/_0043_ ), .B(\us22\/_0058_ ), .Y(\us22\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1227_ ( .A(\us22\/_0195_ ), .B(\us22\/_0233_ ), .C(\us22\/_0320_ ), .D(\us22\/_0435_ ), .X(\us22\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1228_ ( .A(\us22\/_0261_ ), .B(\us22\/_0738_ ), .Y(\us22\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1229_ ( .A1(\us22\/_0218_ ), .A2(\us22\/_0651_ ), .B1(\us22\/_0261_ ), .B2(\us22\/_0056_ ), .Y(\us22\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1230_ ( .A(\us22\/_0436_ ), .B(\us22\/_0394_ ), .C(\us22\/_0437_ ), .D(\us22\/_0438_ ), .X(\us22\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1231_ ( .A(\us22\/_0410_ ), .B(\us22\/_0426_ ), .C(\us22\/_0433_ ), .D(\us22\/_0439_ ), .X(\us22\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us22/_1232_ ( .A(\us22\/_0135_ ), .SLEEP(\us22\/_0273_ ), .X(\us22\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1233_ ( .A1(\us22\/_0279_ ), .A2(\us22\/_0134_ ), .B1(\us22\/_0099_ ), .Y(\us22\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1234_ ( .A(\us22\/_0441_ ), .B(\us22\/_0164_ ), .C(\us22\/_0270_ ), .D(\us22\/_0442_ ), .X(\us22\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1235_ ( .A(\us22\/_0051_ ), .B(\us22\/_0672_ ), .Y(\us22\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1236_ ( .A(\us22\/_0051_ ), .B(\us22\/_0271_ ), .Y(\us22\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1237_ ( .A(\us22\/_0444_ ), .B(\us22\/_0446_ ), .X(\us22\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1238_ ( .A(\us22\/_0193_ ), .B(\us22\/_0304_ ), .X(\us22\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1239_ ( .A(\us22\/_0448_ ), .Y(\us22\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1240_ ( .A(\us22\/_0162_ ), .B(\us22\/_0130_ ), .X(\us22\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1241_ ( .A(\us22\/_0450_ ), .Y(\us22\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1242_ ( .A1(\us22\/_0129_ ), .A2(\us22\/_0554_ ), .B1(\us22\/_0043_ ), .Y(\us22\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1243_ ( .A(\us22\/_0447_ ), .B(\us22\/_0449_ ), .C(\us22\/_0451_ ), .D(\us22\/_0452_ ), .X(\us22\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1244_ ( .A(\us22\/_0056_ ), .B(\us22\/_0064_ ), .Y(\us22\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us22/_1245_ ( .A_N(\us22\/_0248_ ), .B(\us22\/_0454_ ), .C(\us22\/_0254_ ), .D(\us22\/_0256_ ), .X(\us22\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1246_ ( .A1(\us22\/_0330_ ), .A2(\us22\/_0099_ ), .B1(\us22\/_0134_ ), .B2(\us22\/_0705_ ), .Y(\us22\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1247_ ( .A1(\us22\/_0748_ ), .A2(\us22\/_0738_ ), .B1(\us22\/_0092_ ), .B2(\us22\/_0752_ ), .Y(\us22\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1248_ ( .A1(\us22\/_0072_ ), .A2(\us22\/_0036_ ), .B1(\us22\/_0748_ ), .B2(\us22\/_0056_ ), .Y(\us22\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1249_ ( .A1(\us22\/_0748_ ), .A2(\us22\/_0251_ ), .B1(\us22\/_0247_ ), .Y(\us22\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1250_ ( .A(\us22\/_0457_ ), .B(\us22\/_0458_ ), .C(\us22\/_0459_ ), .D(\us22\/_0460_ ), .X(\us22\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1251_ ( .A(\us22\/_0443_ ), .B(\us22\/_0453_ ), .C(\us22\/_0455_ ), .D(\us22\/_0461_ ), .X(\us22\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1252_ ( .A(\us22\/_0705_ ), .B(\us22\/_0080_ ), .X(\us22\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1253_ ( .A(\us22\/_0586_ ), .B(\us22\/_0124_ ), .Y(\us22\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1254_ ( .A(\us22\/_0218_ ), .B(\us22\/_0747_ ), .Y(\us22\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us22/_1255_ ( .A_N(\us22\/_0463_ ), .B(\us22\/_0464_ ), .C(\us22\/_0465_ ), .X(\us22\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us22/_1256_ ( .A1(\us22\/_0271_ ), .A2(\us22\/_0072_ ), .B1(\us22\/_0142_ ), .B2(\us22\/_0027_ ), .X(\us22\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1257_ ( .A1(\us22\/_0144_ ), .A2(\us22\/_0099_ ), .B1(\us22\/_0360_ ), .C1(\us22\/_0468_ ), .Y(\us22\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us22/_1258_ ( .A1(\us22\/_0672_ ), .A2(\us22\/_0251_ ), .B1(\us22\/_0218_ ), .X(\us22\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1259_ ( .A1(\us22\/_0575_ ), .A2(\us22\/_0056_ ), .B1(\us22\/_0379_ ), .C1(\us22\/_0470_ ), .Y(\us22\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1260_ ( .A(\us22\/_0466_ ), .B(\us22\/_0469_ ), .C(\us22\/_0471_ ), .D(\us22\/_0305_ ), .X(\us22\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us22/_1261_ ( .A1(\us22\/_0247_ ), .A2(\us22\/_0683_ ), .B1(\us22\/_0324_ ), .B2(\us22\/_0056_ ), .X(\us22\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1262_ ( .A(\us22\/_0084_ ), .B(\us22\/_0099_ ), .X(\us22\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us22/_1263_ ( .A1(\us22\/_0092_ ), .A2(\us22\/_0247_ ), .B1(\us22\/_0474_ ), .X(\us22\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us22/_1264_ ( .A(\us22\/_0075_ ), .B(\us22\/_0473_ ), .C(\us22\/_0475_ ), .Y(\us22\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1265_ ( .A1(\us22\/_0279_ ), .A2(\us22\/_0255_ ), .B1(\us22\/_0084_ ), .B2(\us22\/_0060_ ), .Y(\us22\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1266_ ( .A1(\us22\/_0093_ ), .A2(\us22\/_0056_ ), .B1(\us22\/_0134_ ), .B2(\us22\/_0114_ ), .Y(\us22\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1267_ ( .A1(\us22\/_0161_ ), .A2(\us22\/_0032_ ), .B1(\us22\/_0324_ ), .B2(\us22\/_0147_ ), .Y(\us22\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1268_ ( .A1(\us22\/_0054_ ), .A2(\us22\/_0732_ ), .B1(\us22\/_0748_ ), .B2(\us22\/_0304_ ), .Y(\us22\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1269_ ( .A(\us22\/_0477_ ), .B(\us22\/_0479_ ), .C(\us22\/_0480_ ), .D(\us22\/_0481_ ), .X(\us22\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1270_ ( .A(\us22\/_0161_ ), .B(\us22\/_0064_ ), .Y(\us22\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us22/_1271_ ( .A(\us22\/_0732_ ), .B(\us22\/_0123_ ), .C(\us22\/_0467_ ), .Y(\us22\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1272_ ( .A(\us22\/_0483_ ), .B(\us22\/_0484_ ), .Y(\us22\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1273_ ( .A(\us22\/_0297_ ), .Y(\us22\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us22/_1274_ ( .A_N(\us22\/_0485_ ), .B(\us22\/_0181_ ), .C(\us22\/_0486_ ), .D(\us22\/_0386_ ), .X(\us22\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1275_ ( .A(\us22\/_0472_ ), .B(\us22\/_0476_ ), .C(\us22\/_0482_ ), .D(\us22\/_0487_ ), .X(\us22\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \us22/_1276_ ( .A(\us22\/_0440_ ), .B(\us22\/_0462_ ), .C(\us22\/_0488_ ), .Y(\us22\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1277_ ( .A(\us22\/_0403_ ), .B(\us22\/_0230_ ), .C(\us22\/_0451_ ), .D(\us22\/_0361_ ), .X(\us22\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1278_ ( .A1(\us22\/_0118_ ), .A2(\us22\/_0050_ ), .B1(\us22\/_0109_ ), .C1(\us22\/_0139_ ), .Y(\us22\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1279_ ( .A(\us22\/_0447_ ), .B(\us22\/_0437_ ), .C(\us22\/_0491_ ), .D(\us22\/_0427_ ), .X(\us22\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1280_ ( .A1(\us22\/_0084_ ), .A2(\us22\/_0255_ ), .B1(\us22\/_0608_ ), .B2(\us22\/_0247_ ), .Y(\us22\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1281_ ( .A1(\us22\/_0144_ ), .A2(\us22\/_0147_ ), .B1(\us22\/_0355_ ), .B2(\us22\/_0093_ ), .Y(\us22\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1282_ ( .A1(\us22\/_0705_ ), .A2(\us22\/_0279_ ), .B1(\us22\/_0330_ ), .B2(\us22\/_0247_ ), .Y(\us22\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1283_ ( .A1(\us22\/_0279_ ), .A2(\us22\/_0084_ ), .B1(\us22\/_0114_ ), .Y(\us22\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1284_ ( .A(\us22\/_0493_ ), .B(\us22\/_0494_ ), .C(\us22\/_0495_ ), .D(\us22\/_0496_ ), .X(\us22\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1285_ ( .A1(\us22\/_0134_ ), .A2(\us22\/_0137_ ), .B1(\us22\/_0355_ ), .B2(\us22\/_0575_ ), .Y(\us22\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1286_ ( .A1(\us22\/_0099_ ), .A2(\us22\/_0733_ ), .B1(\us22\/_0093_ ), .B2(\us22\/_0218_ ), .Y(\us22\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1287_ ( .A(\us22\/_0147_ ), .B(\us22\/_0651_ ), .Y(\us22\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1288_ ( .A1(\us22\/_0153_ ), .A2(\us22\/_0056_ ), .B1(\us22\/_0748_ ), .Y(\us22\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1289_ ( .A(\us22\/_0498_ ), .B(\us22\/_0500_ ), .C(\us22\/_0501_ ), .D(\us22\/_0502_ ), .X(\us22\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1290_ ( .A(\us22\/_0490_ ), .B(\us22\/_0492_ ), .C(\us22\/_0497_ ), .D(\us22\/_0503_ ), .X(\us22\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us22/_1291_ ( .A_N(\us22\/_0275_ ), .B(\us22\/_0705_ ), .X(\us22\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1292_ ( .A(\us22\/_0505_ ), .Y(\us22\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1293_ ( .A(\us22\/_0380_ ), .B(\us22\/_0347_ ), .X(\us22\/_0507_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1294_ ( .A1(\us22\/_0507_ ), .A2(\us22\/_0093_ ), .B1(\us22\/_0056_ ), .Y(\us22\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1295_ ( .A(\us22\/_0322_ ), .B(\us22\/_0277_ ), .C(\us22\/_0506_ ), .D(\us22\/_0508_ ), .X(\us22\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1296_ ( .A(\us22\/_0084_ ), .B(\us22\/_0705_ ), .X(\us22\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1297_ ( .A1(\us22\/_0733_ ), .A2(\us22\/_0114_ ), .B1(\us22\/_0429_ ), .C1(\us22\/_0511_ ), .Y(\us22\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_1298_ ( .A(\us22\/_0019_ ), .B(\us22\/_0024_ ), .Y(\us22\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1299_ ( .A(\us22\/_0512_ ), .B(\us22\/_0513_ ), .C(\us22\/_0742_ ), .D(\us22\/_0306_ ), .X(\us22\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1300_ ( .A1(\us22\/_0532_ ), .A2(\us22\/_0089_ ), .B1(\us22\/_0154_ ), .C1(\us22\/_0169_ ), .Y(\us22\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us22/_1301_ ( .A1(\us22\/_0749_ ), .A2(\us22\/_0026_ ), .B1(\us22\/_0069_ ), .C1(\us22\/_0032_ ), .X(\us22\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us22/_1302_ ( .A1(\us22\/_0324_ ), .A2(\us22\/_0355_ ), .B1(\us22\/_0330_ ), .B2(\us22\/_0727_ ), .X(\us22\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us22/_1303_ ( .A(\us22\/_0133_ ), .B(\us22\/_0516_ ), .C(\us22\/_0517_ ), .Y(\us22\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1304_ ( .A(\us22\/_0509_ ), .B(\us22\/_0514_ ), .C(\us22\/_0515_ ), .D(\us22\/_0518_ ), .X(\us22\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1305_ ( .A(\us22\/_0747_ ), .B(\us22\/_0072_ ), .Y(\us22\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1306_ ( .A1(\us22\/_0082_ ), .A2(\us22\/_0070_ ), .B1(\us22\/_0043_ ), .B2(\us22\/_0193_ ), .Y(\us22\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1307_ ( .A(\us22\/_0311_ ), .B(\us22\/_0520_ ), .C(\us22\/_0332_ ), .D(\us22\/_0522_ ), .X(\us22\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1308_ ( .A(\us22\/_0129_ ), .B(\us22\/_0218_ ), .X(\us22\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_1309_ ( .A(\us22\/_0235_ ), .B(\us22\/_0524_ ), .Y(\us22\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us22/_1310_ ( .A(\us22\/_0081_ ), .B(\us22\/_0085_ ), .Y(\us22\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1311_ ( .A1(\us22\/_0051_ ), .A2(\us22\/_0045_ ), .B1(\us22\/_0130_ ), .B2(\us22\/_0094_ ), .Y(\us22\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1312_ ( .A(\us22\/_0523_ ), .B(\us22\/_0525_ ), .C(\us22\/_0526_ ), .D(\us22\/_0527_ ), .X(\us22\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us22/_1313_ ( .A_N(\us22\/_0250_ ), .B(\us22\/_0521_ ), .Y(\us22\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1314_ ( .A(\us22\/_0128_ ), .B(\us22\/_0021_ ), .X(\us22\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1315_ ( .A(\us22\/_0530_ ), .Y(\us22\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1316_ ( .A(\us22\/_0099_ ), .B(\us22\/_0058_ ), .X(\us22\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1317_ ( .A(\us22\/_0533_ ), .Y(\us22\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us22/_1318_ ( .A_N(\us22\/_0529_ ), .B(\us22\/_0531_ ), .C(\us22\/_0534_ ), .D(\us22\/_0192_ ), .X(\us22\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1319_ ( .A(\us22\/_0434_ ), .B(\us22\/_0078_ ), .X(\us22\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us22/_1320_ ( .A1(\us22\/_0750_ ), .A2(\us22\/_0080_ ), .B1(\us22\/_0129_ ), .B2(\us22\/_0705_ ), .X(\us22\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1321_ ( .A1(\us22\/_0161_ ), .A2(\us22\/_0032_ ), .B1(\us22\/_0536_ ), .C1(\us22\/_0537_ ), .Y(\us22\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us22/_1322_ ( .A1(\us22\/_0747_ ), .A2(\us22\/_0162_ ), .B1(\us22\/_0080_ ), .B2(\us22\/_0043_ ), .X(\us22\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1323_ ( .A1(\us22\/_0093_ ), .A2(\us22\/_0247_ ), .B1(\us22\/_0240_ ), .C1(\us22\/_0539_ ), .Y(\us22\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1324_ ( .A(\us22\/_0434_ ), .B(\us22\/_0043_ ), .X(\us22\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us22/_1325_ ( .A1(\us22\/_0142_ ), .A2(\us22\/_0150_ ), .B1(\us22\/_0023_ ), .B2(\us22\/_0137_ ), .X(\us22\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1326_ ( .A1(\us22\/_0279_ ), .A2(\us22\/_0051_ ), .B1(\us22\/_0541_ ), .C1(\us22\/_0542_ ), .Y(\us22\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1327_ ( .A(\us22\/_0159_ ), .B(\us22\/_0036_ ), .X(\us22\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us22/_1328_ ( .A1(\us22\/_0271_ ), .A2(\us22\/_0434_ ), .B1(\us22\/_0027_ ), .X(\us22\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1329_ ( .A1(\us22\/_0091_ ), .A2(\us22\/_0128_ ), .B1(\us22\/_0545_ ), .C1(\us22\/_0546_ ), .Y(\us22\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1330_ ( .A(\us22\/_0538_ ), .B(\us22\/_0540_ ), .C(\us22\/_0544_ ), .D(\us22\/_0547_ ), .X(\us22\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1331_ ( .A(\us22\/_0099_ ), .B(\us22\/_0193_ ), .X(\us22\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us22/_1332_ ( .A(\us22\/_0549_ ), .B(\us22\/_0186_ ), .C(\us22\/_0187_ ), .Y(\us22\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1333_ ( .A(\us22\/_0062_ ), .B(\us22\/_0347_ ), .C(\us22\/_0749_ ), .D(\us22\/_0694_ ), .X(\us22\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1334_ ( .A1(\us22\/_0130_ ), .A2(\us22\/_0218_ ), .B1(\us22\/_0551_ ), .C1(\us22\/_0101_ ), .Y(\us22\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1335_ ( .A(\us22\/_0139_ ), .B(\us22\/_0651_ ), .Y(\us22\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1336_ ( .A1(\us22\/_0752_ ), .A2(\us22\/_0672_ ), .B1(\us22\/_0084_ ), .B2(\us22\/_0099_ ), .Y(\us22\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1337_ ( .A(\us22\/_0550_ ), .B(\us22\/_0552_ ), .C(\us22\/_0553_ ), .D(\us22\/_0555_ ), .X(\us22\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1338_ ( .A(\us22\/_0528_ ), .B(\us22\/_0535_ ), .C(\us22\/_0548_ ), .D(\us22\/_0556_ ), .X(\us22\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us22/_1339_ ( .A(\us22\/_0504_ ), .B(\us22\/_0519_ ), .C(\us22\/_0557_ ), .Y(\us22\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1340_ ( .A(\us22\/_0054_ ), .B(\us22\/_0507_ ), .X(\us22\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us22/_1341_ ( .A_N(\us22\/_0558_ ), .B(\us22\/_0408_ ), .C(\us22\/_0451_ ), .D(\us22\/_0452_ ), .X(\us22\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1342_ ( .A(\us22\/_0549_ ), .Y(\us22\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1343_ ( .A(\us22\/_0559_ ), .B(\us22\/_0403_ ), .C(\us22\/_0560_ ), .D(\us22\/_0371_ ), .X(\us22\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1344_ ( .A(\us22\/_0181_ ), .B(\us22\/_0178_ ), .X(\us22\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1345_ ( .A(\us22\/_0562_ ), .B(\us22\/_0552_ ), .C(\us22\/_0553_ ), .D(\us22\/_0555_ ), .X(\us22\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1346_ ( .A(\us22\/_0247_ ), .B(\us22\/_0021_ ), .Y(\us22\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1347_ ( .A(\us22\/_0051_ ), .B(\us22\/_0130_ ), .X(\us22\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1348_ ( .A(\us22\/_0566_ ), .Y(\us22\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1349_ ( .A(\us22\/_0159_ ), .B(\us22\/_0423_ ), .X(\us22\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1350_ ( .A1(\us22\/_0752_ ), .A2(\us22\/_0651_ ), .B1(\us22\/_0568_ ), .B2(\us22\/_0175_ ), .Y(\us22\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1351_ ( .A(\us22\/_0076_ ), .B(\us22\/_0565_ ), .C(\us22\/_0567_ ), .D(\us22\/_0569_ ), .X(\us22\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us22/_1352_ ( .A1(\us22\/_0036_ ), .A2(\us22\/_0142_ ), .B1(\us22\/_0161_ ), .X(\us22\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1353_ ( .A(\us22\/_0099_ ), .B(\us22\/_0672_ ), .Y(\us22\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us22/_1354_ ( .A(\us22\/_0420_ ), .B(\us22\/_0571_ ), .C_N(\us22\/_0572_ ), .Y(\us22\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1355_ ( .A(\us22\/_0051_ ), .B(\us22\/_0747_ ), .Y(\us22\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1356_ ( .A(\us22\/_0574_ ), .B(\us22\/_0319_ ), .C(\us22\/_0320_ ), .D(\us22\/_0411_ ), .X(\us22\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1357_ ( .A(\us22\/_0736_ ), .B(\us22\/_0035_ ), .Y(\us22\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1358_ ( .A(\us22\/_0736_ ), .B(\us22\/_0030_ ), .Y(\us22\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1359_ ( .A(\us22\/_0298_ ), .B(\us22\/_0208_ ), .C(\us22\/_0577_ ), .D(\us22\/_0578_ ), .X(\us22\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1360_ ( .A1(\us22\/_0021_ ), .A2(\us22\/_0137_ ), .B1(\us22\/_0261_ ), .B2(\us22\/_0128_ ), .Y(\us22\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1361_ ( .A(\us22\/_0573_ ), .B(\us22\/_0576_ ), .C(\us22\/_0579_ ), .D(\us22\/_0580_ ), .X(\us22\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1362_ ( .A(\us22\/_0561_ ), .B(\us22\/_0563_ ), .C(\us22\/_0570_ ), .D(\us22\/_0581_ ), .X(\us22\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1363_ ( .A(\us22\/_0128_ ), .B(\us22\/_0193_ ), .X(\us22\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1364_ ( .A(\us22\/_0082_ ), .B(\us22\/_0162_ ), .X(\us22\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us22/_1365_ ( .A(\us22\/_0583_ ), .B(\us22\/_0584_ ), .C_N(\us22\/_0437_ ), .Y(\us22\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us22/_1366_ ( .A(\us22\/_0150_ ), .B(\us22\/_0118_ ), .C(\us22\/_0380_ ), .Y(\us22\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us22/_1367_ ( .A_N(\us22\/_0182_ ), .B(\us22\/_0587_ ), .C(\us22\/_0323_ ), .X(\us22\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1368_ ( .A1(\us22\/_0575_ ), .A2(\us22\/_0153_ ), .B1(\us22\/_0727_ ), .B2(\us22\/_0058_ ), .Y(\us22\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1369_ ( .A1(\us22\/_0218_ ), .A2(\us22\/_0064_ ), .B1(\us22\/_0134_ ), .B2(\us22\/_0255_ ), .Y(\us22\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1370_ ( .A(\us22\/_0585_ ), .B(\us22\/_0588_ ), .C(\us22\/_0589_ ), .D(\us22\/_0590_ ), .X(\us22\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us22/_1371_ ( .A1(\us22\/_0091_ ), .A2(\us22\/_0139_ ), .B1(\us22\/_0250_ ), .Y(\us22\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1372_ ( .A1(\us22\/_0092_ ), .A2(\us22\/_0739_ ), .B1(\us22\/_0324_ ), .B2(\us22\/_0247_ ), .Y(\us22\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1373_ ( .A1(\us22\/_0144_ ), .A2(\us22\/_0153_ ), .B1(\us22\/_0683_ ), .B2(\us22\/_0056_ ), .Y(\us22\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1374_ ( .A1(\us22\/_0091_ ), .A2(\us22\/_0218_ ), .B1(\us22\/_0330_ ), .B2(\us22\/_0056_ ), .Y(\us22\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1375_ ( .A(\us22\/_0592_ ), .B(\us22\/_0593_ ), .C(\us22\/_0594_ ), .D(\us22\/_0595_ ), .X(\us22\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1376_ ( .A(\us22\/_0218_ ), .B(\us22\/_0144_ ), .Y(\us22\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1377_ ( .A(\us22\/_0312_ ), .B(\us22\/_0598_ ), .Y(\us22\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1378_ ( .A(\us22\/_0575_ ), .B(\us22\/_0147_ ), .Y(\us22\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1379_ ( .A1(\us22\/_0293_ ), .A2(\us22\/_0137_ ), .B1(\us22\/_0093_ ), .B2(\us22\/_0739_ ), .Y(\us22\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1380_ ( .A1(\us22\/_0734_ ), .A2(\us22\/_0531_ ), .B1(\us22\/_0600_ ), .C1(\us22\/_0601_ ), .Y(\us22\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1381_ ( .A1(\us22\/_0153_ ), .A2(\us22\/_0261_ ), .B1(\us22\/_0599_ ), .C1(\us22\/_0602_ ), .Y(\us22\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1382_ ( .A(\us22\/_0591_ ), .B(\us22\/_0596_ ), .C(\us22\/_0174_ ), .D(\us22\/_0603_ ), .X(\us22\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1383_ ( .A(\us22\/_0247_ ), .B(\us22\/_0144_ ), .Y(\us22\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1384_ ( .A(\us22\/_0113_ ), .B(\us22\/_0018_ ), .Y(\us22\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1385_ ( .A(\us22\/_0381_ ), .B(\us22\/_0605_ ), .C(\us22\/_0361_ ), .D(\us22\/_0606_ ), .X(\us22\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1386_ ( .A1(\us22\/_0016_ ), .A2(\us22\/_0727_ ), .B1(\us22\/_0733_ ), .Y(\us22\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1387_ ( .A1(\us22\/_0586_ ), .A2(\us22\/_0159_ ), .B1(\us22\/_0082_ ), .B2(\us22\/_0750_ ), .Y(\us22\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1388_ ( .A1(\us22\/_0142_ ), .A2(\us22\/_0162_ ), .B1(\us22\/_0080_ ), .B2(\us22\/_0054_ ), .Y(\us22\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1389_ ( .A(\us22\/_0610_ ), .B(\us22\/_0611_ ), .C(\us22\/_0105_ ), .D(\us22\/_0106_ ), .X(\us22\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1390_ ( .A1(\us22\/_0094_ ), .A2(\us22\/_0302_ ), .B1(\us22\/_0324_ ), .B2(\us22\/_0089_ ), .Y(\us22\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1391_ ( .A(\us22\/_0607_ ), .B(\us22\/_0609_ ), .C(\us22\/_0612_ ), .D(\us22\/_0613_ ), .X(\us22\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1392_ ( .A(\us22\/_0041_ ), .B(\us22\/_0170_ ), .X(\us22\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1393_ ( .A(\us22\/_0554_ ), .B(\us22\/_0027_ ), .X(\us22\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1394_ ( .A(\us22\/_0027_ ), .B(\us22\/_0261_ ), .Y(\us22\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us22/_1395_ ( .A_N(\us22\/_0616_ ), .B(\us22\/_0617_ ), .Y(\us22\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1396_ ( .A1(\us22\/_0147_ ), .A2(\us22\/_0302_ ), .B1(\us22\/_0342_ ), .C1(\us22\/_0618_ ), .Y(\us22\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1397_ ( .A(\us22\/_0614_ ), .B(\us22\/_0272_ ), .C(\us22\/_0615_ ), .D(\us22\/_0620_ ), .X(\us22\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us22/_1398_ ( .A(\us22\/_0582_ ), .B(\us22\/_0604_ ), .C(\us22\/_0621_ ), .Y(\us22\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1399_ ( .A1(\us22\/_0084_ ), .A2(\us22\/_0134_ ), .B1(\us22\/_0089_ ), .Y(\us22\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1400_ ( .A1(\us22\/_0144_ ), .A2(\us22\/_0608_ ), .A3(\us22\/_0330_ ), .B1(\us22\/_0089_ ), .Y(\us22\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1401_ ( .A1(\us22\/_0197_ ), .A2(\us22\/_0130_ ), .A3(\us22\/_0110_ ), .B1(\us22\/_0094_ ), .Y(\us22\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1402_ ( .A(\us22\/_0432_ ), .B(\us22\/_0622_ ), .C(\us22\/_0623_ ), .D(\us22\/_0624_ ), .X(\us22\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us22/_1403_ ( .A1(\us22\/_0554_ ), .A2(\us22\/_0018_ ), .A3(\us22\/_0023_ ), .B1(\us22\/_0161_ ), .X(\us22\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us22/_1404_ ( .A_N(\us22\/_0269_ ), .B(\us22\/_0170_ ), .X(\us22\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1405_ ( .A1(\us22\/_0109_ ), .A2(\us22\/_0064_ ), .A3(\us22\/_0733_ ), .B1(\us22\/_0355_ ), .Y(\us22\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us22/_1406_ ( .A_N(\us22\/_0626_ ), .B(\us22\/_0627_ ), .C(\us22\/_0353_ ), .D(\us22\/_0628_ ), .X(\us22\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1407_ ( .A1(\us22\/_0091_ ), .A2(\us22\/_0110_ ), .A3(\us22\/_0176_ ), .B1(\us22\/_0139_ ), .Y(\us22\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1408_ ( .A1(\us22\/_0021_ ), .A2(\us22\/_0261_ ), .B1(\us22\/_0147_ ), .Y(\us22\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1409_ ( .A(\us22\/_0631_ ), .B(\us22\/_0344_ ), .C(\us22\/_0421_ ), .D(\us22\/_0632_ ), .X(\us22\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us22/_1410_ ( .A1(\us22\/_0325_ ), .A2(\us22\/_0734_ ), .B1(\us22\/_0038_ ), .C1(\us22\/_0113_ ), .X(\us22\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1411_ ( .A1(\us22\/_0134_ ), .A2(\us22\/_0114_ ), .B1(\us22\/_0221_ ), .C1(\us22\/_0634_ ), .Y(\us22\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us22/_1412_ ( .A(\us22\/_0119_ ), .B_N(\us22\/_0111_ ), .Y(\us22\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1413_ ( .A1(\us22\/_0032_ ), .A2(\us22\/_0113_ ), .B1(\us22\/_0636_ ), .C1(\us22\/_0400_ ), .Y(\us22\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1414_ ( .A1(\us22\/_0732_ ), .A2(\us22\/_0293_ ), .A3(\us22\/_0251_ ), .B1(\us22\/_0099_ ), .Y(\us22\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1415_ ( .A(\us22\/_0189_ ), .B(\us22\/_0635_ ), .C(\us22\/_0637_ ), .D(\us22\/_0638_ ), .X(\us22\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1416_ ( .A(\us22\/_0625_ ), .B(\us22\/_0630_ ), .C(\us22\/_0633_ ), .D(\us22\/_0639_ ), .X(\us22\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1417_ ( .A(\us22\/_0747_ ), .B(\us22\/_0738_ ), .X(\us22\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1418_ ( .A(\us22\/_0736_ ), .B(\us22\/_0731_ ), .X(\us22\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us22/_1419_ ( .A_N(\us22\/_0643_ ), .B(\us22\/_0577_ ), .Y(\us22\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1420_ ( .A1(\us22\/_0084_ ), .A2(\us22\/_0739_ ), .B1(\us22\/_0642_ ), .C1(\us22\/_0644_ ), .Y(\us22\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1421_ ( .A1(\us22\/_0050_ ), .A2(\us22\/_0543_ ), .B1(\us22\/_0194_ ), .C1(\us22\/_0738_ ), .Y(\us22\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1422_ ( .A(\us22\/_0646_ ), .B(\us22\/_0232_ ), .C(\us22\/_0417_ ), .D(\us22\/_0578_ ), .X(\us22\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1423_ ( .A1(\us22\/_0064_ ), .A2(\us22\/_0733_ ), .B1(\us22\/_0727_ ), .Y(\us22\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1424_ ( .A1(\us22\/_0193_ ), .A2(\us22\/_0276_ ), .B1(\us22\/_0727_ ), .Y(\us22\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1425_ ( .A(\us22\/_0645_ ), .B(\us22\/_0647_ ), .C(\us22\/_0648_ ), .D(\us22\/_0649_ ), .X(\us22\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1426_ ( .A1(\us22\/_0325_ ), .A2(\us22\/_0734_ ), .B1(\us22\/_0038_ ), .C1(\us22\/_0247_ ), .Y(\us22\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1427_ ( .A1(\us22\/_0543_ ), .A2(\us22\/_0216_ ), .B1(\us22\/_0423_ ), .C1(\us22\/_0247_ ), .Y(\us22\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1428_ ( .A(\us22\/_0652_ ), .B(\us22\/_0653_ ), .X(\us22\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1429_ ( .A1(\us22\/_0733_ ), .A2(\us22\/_0748_ ), .A3(\us22\/_0324_ ), .B1(\us22\/_0016_ ), .Y(\us22\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1430_ ( .A1(\us22\/_0651_ ), .A2(\us22\/_0193_ ), .A3(\us22\/_0091_ ), .B1(\us22\/_0016_ ), .Y(\us22\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1431_ ( .A1(\us22\/_0102_ ), .A2(\us22\/_0301_ ), .B1(\sa22\[3\] ), .C1(\us22\/_0247_ ), .Y(\us22\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1432_ ( .A(\us22\/_0654_ ), .B(\us22\/_0655_ ), .C(\us22\/_0656_ ), .D(\us22\/_0657_ ), .X(\us22\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1433_ ( .A1(\us22\/_0118_ ), .A2(\us22\/_0050_ ), .B1(\us22\/_0038_ ), .C1(\us22\/_0478_ ), .Y(\us22\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us22/_1434_ ( .A_N(\us22\/_0250_ ), .B(\us22\/_0465_ ), .C(\us22\/_0659_ ), .X(\us22\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1435_ ( .A1(\us22\/_0683_ ), .A2(\us22\/_0324_ ), .B1(\us22\/_0255_ ), .Y(\us22\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1436_ ( .A1(\us22\/_0032_ ), .A2(\us22\/_0193_ ), .A3(\us22\/_0047_ ), .B1(\us22\/_0255_ ), .Y(\us22\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1437_ ( .A1(\us22\/_0144_ ), .A2(\us22\/_0586_ ), .A3(\us22\/_0047_ ), .B1(\us22\/_0218_ ), .Y(\us22\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1438_ ( .A(\us22\/_0660_ ), .B(\us22\/_0661_ ), .C(\us22\/_0663_ ), .D(\us22\/_0664_ ), .X(\us22\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1439_ ( .A1(\us22\/_0091_ ), .A2(\us22\/_0276_ ), .B1(\us22\/_0060_ ), .Y(\us22\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1440_ ( .A1(\us22\/_0144_ ), .A2(\us22\/_0608_ ), .B1(\us22\/_0056_ ), .Y(\us22\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1441_ ( .A1(\us22\/_0423_ ), .A2(\us22\/_0038_ ), .B1(\us22\/_0102_ ), .C1(\us22\/_0060_ ), .Y(\us22\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1442_ ( .A1(\sa22\[1\] ), .A2(\us22\/_0734_ ), .B1(\us22\/_0109_ ), .C1(\us22\/_0056_ ), .Y(\us22\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1443_ ( .A(\us22\/_0666_ ), .B(\us22\/_0667_ ), .C(\us22\/_0668_ ), .D(\us22\/_0669_ ), .X(\us22\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1444_ ( .A(\us22\/_0650_ ), .B(\us22\/_0658_ ), .C(\us22\/_0665_ ), .D(\us22\/_0670_ ), .X(\us22\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us22/_1445_ ( .A(\us22\/_0641_ ), .B(\us22\/_0174_ ), .C(\us22\/_0671_ ), .Y(\us22\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us22/_1446_ ( .A(\us22\/_0049_ ), .B(\us22\/_0618_ ), .C_N(\us22\/_0052_ ), .Y(\us22\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us22/_1447_ ( .A(\us22\/_0239_ ), .Y(\us22\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1448_ ( .A(\us22\/_0705_ ), .B(\us22\/_0032_ ), .Y(\us22\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1449_ ( .A1(\us22\/_0054_ ), .A2(\us22\/_0732_ ), .B1(\us22\/_0036_ ), .B2(\us22\/_0705_ ), .Y(\us22\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1450_ ( .A1(\us22\/_0304_ ), .A2(\us22\/_0732_ ), .B1(\us22\/_0047_ ), .B2(\us22\/_0750_ ), .Y(\us22\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1451_ ( .A(\us22\/_0674_ ), .B(\us22\/_0675_ ), .C(\us22\/_0676_ ), .D(\us22\/_0677_ ), .X(\us22\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us22/_1452_ ( .A_N(\us22\/_0584_ ), .B(\us22\/_0283_ ), .X(\us22\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1453_ ( .A(\us22\/_0673_ ), .B(\us22\/_0678_ ), .C(\us22\/_0679_ ), .D(\us22\/_0508_ ), .X(\us22\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1454_ ( .A1(\us22\/_0016_ ), .A2(\us22\/_0733_ ), .B1(\us22\/_0355_ ), .B2(\us22\/_0092_ ), .Y(\us22\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1455_ ( .A(\us22\/_0681_ ), .B(\us22\/_0034_ ), .X(\us22\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us22/_1456_ ( .A1(\us22\/_0330_ ), .A2(\us22\/_0139_ ), .B1(\us22\/_0324_ ), .B2(\us22\/_0089_ ), .X(\us22\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1457_ ( .A1(\us22\/_0146_ ), .A2(\us22\/_0147_ ), .B1(\us22\/_0133_ ), .C1(\us22\/_0684_ ), .Y(\us22\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1458_ ( .A(\us22\/_0113_ ), .B(\us22\/_0251_ ), .Y(\us22\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us22/_1459_ ( .A_N(\us22\/_0463_ ), .B(\us22\/_0686_ ), .C(\us22\/_0383_ ), .D(\us22\/_0464_ ), .X(\us22\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1460_ ( .A1(\us22\/_0051_ ), .A2(\us22\/_0293_ ), .B1(\us22\/_0084_ ), .B2(\us22\/_0705_ ), .Y(\us22\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1461_ ( .A1(\us22\/_0018_ ), .A2(\us22\/_0072_ ), .B1(\us22\/_0134_ ), .B2(\us22\/_0078_ ), .Y(\us22\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1462_ ( .A(\us22\/_0687_ ), .B(\us22\/_0236_ ), .C(\us22\/_0688_ ), .D(\us22\/_0689_ ), .X(\us22\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1463_ ( .A(\us22\/_0680_ ), .B(\us22\/_0682_ ), .C(\us22\/_0685_ ), .D(\us22\/_0690_ ), .X(\us22\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us22/_1464_ ( .A1(\us22\/_0532_ ), .A2(\us22\/_0380_ ), .B1(\us22\/_0102_ ), .C1(\us22\/_0355_ ), .X(\us22\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us22/_1465_ ( .A(\us22\/_0692_ ), .B(\us22\/_0338_ ), .C(\us22\/_0644_ ), .Y(\us22\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1466_ ( .A(\us22\/_0016_ ), .B(\us22\/_0021_ ), .Y(\us22\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1467_ ( .A1(\us22\/_0032_ ), .A2(\us22\/_0137_ ), .B1(\us22\/_0279_ ), .B2(\us22\/_0094_ ), .Y(\us22\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1468_ ( .A1(\us22\/_0575_ ), .A2(\us22\/_0153_ ), .B1(\us22\/_0161_ ), .B2(\us22\/_0293_ ), .Y(\us22\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1469_ ( .A(\us22\/_0259_ ), .B(\us22\/_0695_ ), .C(\us22\/_0696_ ), .D(\us22\/_0697_ ), .X(\us22\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us22/_1470_ ( .A1(\us22\/_0255_ ), .A2(\us22\/_0651_ ), .B1(\us22\/_0016_ ), .B2(\us22\/_0193_ ), .X(\us22\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1471_ ( .A1(\us22\/_0060_ ), .A2(\us22\/_0176_ ), .B1(\us22\/_0699_ ), .C1(\us22\/_0177_ ), .Y(\us22\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1472_ ( .A1(\us22\/_0091_ ), .A2(\us22\/_0218_ ), .B1(\us22\/_0092_ ), .B2(\us22\/_0705_ ), .Y(\us22\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us22/_1473_ ( .A1(\us22\/_0705_ ), .A2(\us22\/_0683_ ), .B1(\us22\/_0093_ ), .B2(\us22\/_0114_ ), .Y(\us22\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us22/_1474_ ( .A1(\us22\/_0683_ ), .A2(\us22\/_0084_ ), .B1(\us22\/_0094_ ), .Y(\us22\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us22/_1475_ ( .A1(\us22\/_0543_ ), .A2(\us22\/_0216_ ), .B1(\us22\/_0038_ ), .C1(\us22\/_0056_ ), .Y(\us22\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1476_ ( .A(\us22\/_0701_ ), .B(\us22\/_0702_ ), .C(\us22\/_0703_ ), .D(\us22\/_0704_ ), .X(\us22\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1477_ ( .A(\us22\/_0693_ ), .B(\us22\/_0698_ ), .C(\us22\/_0700_ ), .D(\us22\/_0706_ ), .X(\us22\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us22/_1478_ ( .A1(\us22\/_0113_ ), .A2(\us22\/_0640_ ), .B1(\us22\/_0099_ ), .B2(\us22\/_0058_ ), .X(\us22\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us22/_1479_ ( .A(\us22\/_0407_ ), .B(\us22\/_0708_ ), .C(\us22\/_0529_ ), .Y(\us22\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1480_ ( .A(\us22\/_0568_ ), .B(\us22\/_0175_ ), .Y(\us22\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us22/_1481_ ( .A1(\us22\/_0247_ ), .A2(\us22\/_0114_ ), .A3(\us22\/_0051_ ), .B1(\us22\/_0130_ ), .Y(\us22\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1482_ ( .A(\us22\/_0709_ ), .B(\us22\/_0550_ ), .C(\us22\/_0710_ ), .D(\us22\/_0711_ ), .X(\us22\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us22/_1483_ ( .A1(\us22\/_0114_ ), .A2(\us22\/_0064_ ), .B1(\us22\/_0261_ ), .B2(\us22\/_0089_ ), .X(\us22\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1484_ ( .A1(\us22\/_0355_ ), .A2(\us22\/_0261_ ), .B1(\us22\/_0198_ ), .C1(\us22\/_0713_ ), .Y(\us22\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1485_ ( .A(\us22\/_0586_ ), .B(\us22\/_0478_ ), .Y(\us22\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us22/_1486_ ( .A_N(\us22\/_0541_ ), .B(\us22\/_0267_ ), .C(\us22\/_0715_ ), .D(\us22\/_0320_ ), .X(\us22\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1487_ ( .A(\us22\/_0586_ ), .B(\us22\/_0070_ ), .Y(\us22\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us22/_1488_ ( .A_N(\us22\/_0211_ ), .B(\us22\/_0155_ ), .C(\us22\/_0202_ ), .D(\us22\/_0718_ ), .X(\us22\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us22/_1489_ ( .A(\us22\/_0150_ ), .B(\us22\/_0216_ ), .C(\us22\/_0380_ ), .Y(\us22\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us22/_1490_ ( .A(\us22\/_0411_ ), .B(\us22\/_0720_ ), .X(\us22\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us22/_1491_ ( .A1(\us22\/_0018_ ), .A2(\us22\/_0023_ ), .B1(\us22\/_0078_ ), .X(\us22\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us22/_1492_ ( .A1(\us22\/_0134_ ), .A2(\us22\/_0738_ ), .B1(\us22\/_0101_ ), .C1(\us22\/_0722_ ), .Y(\us22\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1493_ ( .A(\us22\/_0717_ ), .B(\us22\/_0719_ ), .C(\us22\/_0721_ ), .D(\us22\/_0723_ ), .X(\us22\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us22/_1494_ ( .A(\us22\/_0739_ ), .B(\us22\/_0193_ ), .Y(\us22\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1495_ ( .A(\us22\/_0344_ ), .B(\us22\/_0184_ ), .C(\us22\/_0449_ ), .D(\us22\/_0725_ ), .X(\us22\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us22/_1496_ ( .A(\us22\/_0712_ ), .B(\us22\/_0714_ ), .C(\us22\/_0724_ ), .D(\us22\/_0726_ ), .X(\us22\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \us22/_1497_ ( .A(\us22\/_0691_ ), .B(\us22\/_0707_ ), .C(\us22\/_0728_ ), .Y(\us22\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \us23/_0753_ ( .A(\sa23\[2\] ), .B_N(\sa23\[3\] ), .Y(\us23\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \us23/_0755_ ( .A(\sa23\[1\] ), .B(\sa23\[0\] ), .X(\us23\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us23/_0756_ ( .A(\us23\/_0096_ ), .B(\us23\/_0118_ ), .X(\us23\/_0129_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0757_ ( .A(\sa23\[7\] ), .B(\sa23\[6\] ), .X(\us23\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_0758_ ( .A(\sa23\[4\] ), .B(\sa23\[5\] ), .Y(\us23\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0759_ ( .A(\us23\/_0140_ ), .B(\us23\/_0151_ ), .X(\us23\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0761_ ( .A(\us23\/_0129_ ), .B(\us23\/_0162_ ), .X(\us23\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0762_ ( .A(\us23\/_0096_ ), .X(\us23\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \us23/_0763_ ( .A(\sa23\[1\] ), .B_N(\sa23\[0\] ), .Y(\us23\/_0205_ ) );
sky130_fd_sc_hd__and3_1 \us23/_0765_ ( .A(\us23\/_0162_ ), .B(\us23\/_0194_ ), .C(\us23\/_0205_ ), .X(\us23\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us23/_0766_ ( .A(\us23\/_0183_ ), .SLEEP(\us23\/_0227_ ), .X(\us23\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \us23/_0767_ ( .A(\sa23\[0\] ), .B_N(\sa23\[1\] ), .Y(\us23\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_0768_ ( .A(\sa23\[2\] ), .B(\sa23\[3\] ), .Y(\us23\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0769_ ( .A(\us23\/_0249_ ), .B(\us23\/_0260_ ), .X(\us23\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0771_ ( .A(\us23\/_0271_ ), .X(\us23\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0772_ ( .A(\us23\/_0162_ ), .X(\us23\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_0773_ ( .A(\us23\/_0293_ ), .B(\us23\/_0304_ ), .Y(\us23\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us23/_0774_ ( .A(\sa23\[1\] ), .Y(\us23\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us23/_0776_ ( .A(\sa23\[0\] ), .Y(\us23\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0777_ ( .A(\sa23\[2\] ), .B(\sa23\[3\] ), .X(\us23\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0779_ ( .A(\us23\/_0358_ ), .X(\us23\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_0780_ ( .A1(\us23\/_0325_ ), .A2(\us23\/_0347_ ), .B1(\us23\/_0380_ ), .C1(\us23\/_0304_ ), .Y(\us23\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us23/_0781_ ( .A_N(\us23\/_0238_ ), .B(\us23\/_0314_ ), .C(\us23\/_0391_ ), .X(\us23\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us23/_0782_ ( .A(\sa23\[3\] ), .B_N(\sa23\[2\] ), .Y(\us23\/_0412_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0783_ ( .A(\us23\/_0412_ ), .X(\us23\/_0423_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0784_ ( .A(\us23\/_0423_ ), .B(\us23\/_0205_ ), .X(\us23\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \us23/_0787_ ( .A(\sa23\[5\] ), .B_N(\sa23\[4\] ), .Y(\us23\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0788_ ( .A(\us23\/_0467_ ), .B(\us23\/_0140_ ), .X(\us23\/_0478_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_0791_ ( .A(\us23\/_0134_ ), .B(\us23\/_0218_ ), .Y(\us23\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_0792_ ( .A(\us23\/_0478_ ), .B(\us23\/_0271_ ), .Y(\us23\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0793_ ( .A(\us23\/_0194_ ), .X(\us23\/_0532_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0794_ ( .A(\us23\/_0249_ ), .X(\us23\/_0543_ ) );
sky130_fd_sc_hd__and2_1 \us23/_0795_ ( .A(\us23\/_0543_ ), .B(\us23\/_0358_ ), .X(\us23\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0797_ ( .A(\us23\/_0554_ ), .X(\us23\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us23/_0798_ ( .A(\us23\/_0205_ ), .B(\us23\/_0358_ ), .X(\us23\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0800_ ( .A(\us23\/_0586_ ), .X(\us23\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_0801_ ( .A1(\us23\/_0532_ ), .A2(\us23\/_0575_ ), .A3(\us23\/_0608_ ), .B1(\us23\/_0218_ ), .Y(\us23\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us23/_0802_ ( .A(\us23\/_0401_ ), .B(\us23\/_0510_ ), .C(\us23\/_0521_ ), .D(\us23\/_0619_ ), .X(\us23\/_0629_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0803_ ( .A(\us23\/_0358_ ), .B(\sa23\[1\] ), .X(\us23\/_0640_ ) );
sky130_fd_sc_hd__and2_1 \us23/_0805_ ( .A(\us23\/_0205_ ), .B(\us23\/_0260_ ), .X(\us23\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0807_ ( .A(\us23\/_0662_ ), .X(\us23\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us23/_0808_ ( .A(\sa23\[6\] ), .B_N(\sa23\[7\] ), .Y(\us23\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \us23/_0809_ ( .A(\us23\/_0467_ ), .B(\us23\/_0694_ ), .X(\us23\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0811_ ( .A(\us23\/_0705_ ), .X(\us23\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_0812_ ( .A1(\us23\/_0640_ ), .A2(\us23\/_0293_ ), .A3(\us23\/_0683_ ), .B1(\us23\/_0727_ ), .Y(\us23\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_0813_ ( .A(\sa23\[1\] ), .B(\sa23\[0\] ), .Y(\us23\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0814_ ( .A(\us23\/_0730_ ), .B(\us23\/_0260_ ), .X(\us23\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0816_ ( .A(\us23\/_0731_ ), .X(\us23\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0817_ ( .A(\sa23\[0\] ), .X(\us23\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us23/_0818_ ( .A1(\us23\/_0325_ ), .A2(\us23\/_0734_ ), .B1(\us23\/_0423_ ), .X(\us23\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0819_ ( .A(\us23\/_0694_ ), .B(\us23\/_0151_ ), .X(\us23\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0821_ ( .A(\us23\/_0736_ ), .X(\us23\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0822_ ( .A(\us23\/_0738_ ), .X(\us23\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_0823_ ( .A1(\us23\/_0733_ ), .A2(\us23\/_0735_ ), .A3(\us23\/_0293_ ), .B1(\us23\/_0739_ ), .Y(\us23\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us23/_0824_ ( .A(\us23\/_0730_ ), .B_N(\us23\/_0358_ ), .Y(\us23\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_0825_ ( .A(\us23\/_0741_ ), .B(\us23\/_0739_ ), .Y(\us23\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_0827_ ( .A1(\us23\/_0118_ ), .A2(\us23\/_0205_ ), .B1(\us23\/_0532_ ), .C1(\us23\/_0739_ ), .Y(\us23\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us23/_0828_ ( .A(\us23\/_0729_ ), .B(\us23\/_0740_ ), .C(\us23\/_0742_ ), .D(\us23\/_0744_ ), .X(\us23\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0829_ ( .A(\us23\/_0423_ ), .B(\us23\/_0730_ ), .X(\us23\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0831_ ( .A(\us23\/_0746_ ), .X(\us23\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us23/_0832_ ( .A(\sa23\[4\] ), .B_N(\sa23\[5\] ), .Y(\us23\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0833_ ( .A(\us23\/_0749_ ), .B(\us23\/_0694_ ), .X(\us23\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0835_ ( .A(\us23\/_0750_ ), .X(\us23\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0836_ ( .A(\us23\/_0752_ ), .X(\us23\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0837_ ( .A(\us23\/_0118_ ), .B(\us23\/_0358_ ), .X(\us23\/_0017_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0839_ ( .A(\us23\/_0752_ ), .B(\us23\/_0017_ ), .X(\us23\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0840_ ( .A(\us23\/_0358_ ), .B(\us23\/_0325_ ), .X(\us23\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0842_ ( .A(\us23\/_0096_ ), .B(\us23\/_0205_ ), .X(\us23\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \us23/_0844_ ( .A1(\us23\/_0020_ ), .A2(\us23\/_0022_ ), .B1(\us23\/_0752_ ), .X(\us23\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_0845_ ( .A1(\us23\/_0748_ ), .A2(\us23\/_0016_ ), .B1(\us23\/_0019_ ), .C1(\us23\/_0024_ ), .Y(\us23\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \us23/_0846_ ( .A(\sa23\[4\] ), .B(\sa23\[5\] ), .X(\us23\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0847_ ( .A(\us23\/_0694_ ), .B(\us23\/_0026_ ), .X(\us23\/_0027_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0850_ ( .A(\us23\/_0358_ ), .B(\us23\/_0730_ ), .X(\us23\/_0030_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0852_ ( .A(\us23\/_0030_ ), .X(\us23\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_0853_ ( .A(\us23\/_0247_ ), .B(\us23\/_0032_ ), .Y(\us23\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_0854_ ( .A(\us23\/_0247_ ), .B(\us23\/_0735_ ), .Y(\us23\/_0034_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0855_ ( .A(\us23\/_0118_ ), .B(\us23\/_0260_ ), .X(\us23\/_0035_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0857_ ( .A(\us23\/_0027_ ), .B(\us23\/_0035_ ), .X(\us23\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0858_ ( .A(\us23\/_0260_ ), .X(\us23\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_0859_ ( .A(\us23\/_0038_ ), .B(\us23\/_0347_ ), .Y(\us23\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us23/_0860_ ( .A_N(\us23\/_0039_ ), .B(\us23\/_0027_ ), .X(\us23\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_0861_ ( .A(\us23\/_0037_ ), .B(\us23\/_0040_ ), .Y(\us23\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us23/_0862_ ( .A(\us23\/_0025_ ), .B(\us23\/_0033_ ), .C(\us23\/_0034_ ), .D(\us23\/_0041_ ), .X(\us23\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0863_ ( .A(\us23\/_0749_ ), .B(\us23\/_0140_ ), .X(\us23\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us23/_0865_ ( .A(\sa23\[0\] ), .B(\sa23\[2\] ), .C(\sa23\[3\] ), .X(\us23\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0866_ ( .A(\us23\/_0043_ ), .B(\us23\/_0045_ ), .X(\us23\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0867_ ( .A(\us23\/_0096_ ), .B(\us23\/_0543_ ), .X(\us23\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0869_ ( .A(\us23\/_0047_ ), .B(\us23\/_0043_ ), .X(\us23\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0870_ ( .A(\us23\/_0730_ ), .X(\us23\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0871_ ( .A(\us23\/_0043_ ), .X(\us23\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_0872_ ( .A1(\us23\/_0118_ ), .A2(\us23\/_0050_ ), .B1(\us23\/_0194_ ), .C1(\us23\/_0051_ ), .Y(\us23\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us23/_0873_ ( .A(\us23\/_0046_ ), .B(\us23\/_0049_ ), .C_N(\us23\/_0052_ ), .Y(\us23\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0874_ ( .A(\us23\/_0026_ ), .B(\us23\/_0140_ ), .X(\us23\/_0054_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0876_ ( .A(\us23\/_0054_ ), .X(\us23\/_0056_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_0877_ ( .A1(\us23\/_0532_ ), .A2(\us23\/_0575_ ), .B1(\us23\/_0056_ ), .Y(\us23\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0878_ ( .A(\us23\/_0423_ ), .B(\us23\/_0325_ ), .X(\us23\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0880_ ( .A(\us23\/_0051_ ), .X(\us23\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_0881_ ( .A1(\us23\/_0731_ ), .A2(\us23\/_0035_ ), .A3(\us23\/_0058_ ), .B1(\us23\/_0060_ ), .Y(\us23\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0882_ ( .A(\us23\/_0260_ ), .B(\sa23\[1\] ), .X(\us23\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0884_ ( .A(\us23\/_0062_ ), .X(\us23\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_0885_ ( .A1(\us23\/_0064_ ), .A2(\us23\/_0748_ ), .A3(\us23\/_0683_ ), .B1(\us23\/_0056_ ), .Y(\us23\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us23/_0886_ ( .A(\us23\/_0053_ ), .B(\us23\/_0057_ ), .C(\us23\/_0061_ ), .D(\us23\/_0065_ ), .X(\us23\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us23/_0887_ ( .A(\us23\/_0629_ ), .B(\us23\/_0745_ ), .C(\us23\/_0042_ ), .D(\us23\/_0066_ ), .X(\us23\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us23/_0889_ ( .A(\sa23\[7\] ), .B_N(\sa23\[6\] ), .Y(\us23\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0890_ ( .A(\us23\/_0069_ ), .B(\us23\/_0151_ ), .X(\us23\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0892_ ( .A(\us23\/_0070_ ), .X(\us23\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_0893_ ( .A1(\us23\/_0129_ ), .A2(\us23\/_0586_ ), .B1(\us23\/_0072_ ), .Y(\us23\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_0894_ ( .A1(\us23\/_0380_ ), .A2(\us23\/_0347_ ), .B1(\us23\/_0194_ ), .B2(\us23\/_0205_ ), .Y(\us23\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us23/_0895_ ( .A(\us23\/_0074_ ), .B_N(\us23\/_0070_ ), .Y(\us23\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us23/_0896_ ( .A(\us23\/_0073_ ), .SLEEP(\us23\/_0075_ ), .X(\us23\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us23/_0897_ ( .A(\us23\/_0467_ ), .B(\us23\/_0069_ ), .X(\us23\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0898_ ( .A(\us23\/_0077_ ), .X(\us23\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0899_ ( .A(\us23\/_0412_ ), .B(\us23\/_0118_ ), .X(\us23\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0901_ ( .A(\us23\/_0078_ ), .B(\us23\/_0079_ ), .X(\us23\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0902_ ( .A(\us23\/_0412_ ), .B(\us23\/_0249_ ), .X(\us23\/_0082_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0905_ ( .A(\us23\/_0280_ ), .B(\us23\/_0078_ ), .X(\us23\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us23/_0906_ ( .A1(\sa23\[0\] ), .A2(\us23\/_0325_ ), .B1(\us23\/_0260_ ), .Y(\us23\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us23/_0907_ ( .A_N(\us23\/_0086_ ), .B(\us23\/_0078_ ), .X(\us23\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us23/_0908_ ( .A(\us23\/_0081_ ), .B(\us23\/_0085_ ), .C(\us23\/_0087_ ), .Y(\us23\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0909_ ( .A(\us23\/_0072_ ), .X(\us23\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_0910_ ( .A1(\us23\/_0733_ ), .A2(\us23\/_0748_ ), .A3(\us23\/_0683_ ), .B1(\us23\/_0089_ ), .Y(\us23\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0911_ ( .A(\us23\/_0129_ ), .X(\us23\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0912_ ( .A(\us23\/_0017_ ), .X(\us23\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0913_ ( .A(\us23\/_0022_ ), .X(\us23\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0914_ ( .A(\us23\/_0078_ ), .X(\us23\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_0915_ ( .A1(\us23\/_0091_ ), .A2(\us23\/_0092_ ), .A3(\us23\/_0093_ ), .B1(\us23\/_0094_ ), .Y(\us23\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us23/_0916_ ( .A(\us23\/_0076_ ), .B(\us23\/_0088_ ), .C(\us23\/_0090_ ), .D(\us23\/_0095_ ), .X(\us23\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us23/_0917_ ( .A(\us23\/_0069_ ), .B(\us23\/_0026_ ), .X(\us23\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \us23/_0918_ ( .A(\us23\/_0098_ ), .X(\us23\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0919_ ( .A(\us23\/_0434_ ), .B(\us23\/_0099_ ), .X(\us23\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0920_ ( .A(\us23\/_0079_ ), .B(\us23\/_0098_ ), .X(\us23\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0921_ ( .A(\us23\/_0325_ ), .X(\us23\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_0922_ ( .A1(\us23\/_0102_ ), .A2(\us23\/_0734_ ), .B1(\us23\/_0038_ ), .C1(\us23\/_0099_ ), .Y(\us23\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us23/_0923_ ( .A(\us23\/_0100_ ), .B(\us23\/_0101_ ), .C_N(\us23\/_0103_ ), .Y(\us23\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_0924_ ( .A1(\us23\/_0554_ ), .A2(\us23\/_0586_ ), .B1(\us23\/_0099_ ), .Y(\us23\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_0925_ ( .A(\us23\/_0129_ ), .B(\us23\/_0099_ ), .Y(\us23\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0926_ ( .A(\us23\/_0105_ ), .B(\us23\/_0106_ ), .X(\us23\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0927_ ( .A(\us23\/_0423_ ), .X(\us23\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us23/_0928_ ( .A(\us23\/_0260_ ), .B(\sa23\[0\] ), .X(\us23\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0929_ ( .A(\us23\/_0069_ ), .B(\us23\/_0749_ ), .X(\us23\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0931_ ( .A(\us23\/_0111_ ), .X(\us23\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0932_ ( .A(\us23\/_0113_ ), .X(\us23\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_0933_ ( .A1(\us23\/_0109_ ), .A2(\us23\/_0110_ ), .B1(\us23\/_0114_ ), .Y(\us23\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us23/_0934_ ( .A(\us23\/_0022_ ), .Y(\us23\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us23/_0935_ ( .A(\us23\/_0554_ ), .Y(\us23\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us23/_0936_ ( .A1(\us23\/_0050_ ), .A2(\us23\/_0118_ ), .B1(\us23\/_0194_ ), .Y(\us23\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us23/_0937_ ( .A(\us23\/_0113_ ), .Y(\us23\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us23/_0938_ ( .A1(\us23\/_0116_ ), .A2(\us23\/_0117_ ), .A3(\us23\/_0119_ ), .B1(\us23\/_0120_ ), .X(\us23\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us23/_0939_ ( .A(\us23\/_0104_ ), .B(\us23\/_0108_ ), .C(\us23\/_0115_ ), .D(\us23\/_0121_ ), .X(\us23\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_0940_ ( .A(\sa23\[7\] ), .B(\sa23\[6\] ), .Y(\us23\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0941_ ( .A(\us23\/_0749_ ), .B(\us23\/_0123_ ), .X(\us23\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0943_ ( .A(\us23\/_0082_ ), .B(\us23\/_0124_ ), .X(\us23\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_0944_ ( .A(\us23\/_0271_ ), .B(\us23\/_0124_ ), .Y(\us23\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0945_ ( .A(\us23\/_0124_ ), .X(\us23\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0946_ ( .A(\us23\/_0260_ ), .B(\us23\/_0325_ ), .X(\us23\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_0948_ ( .A(\us23\/_0128_ ), .B(\us23\/_0130_ ), .Y(\us23\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_0949_ ( .A(\us23\/_0127_ ), .B(\us23\/_0132_ ), .Y(\us23\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us23/_0950_ ( .A(\us23\/_0434_ ), .X(\us23\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_0951_ ( .A(\us23\/_0134_ ), .B(\us23\/_0128_ ), .Y(\us23\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us23/_0952_ ( .A(\us23\/_0126_ ), .B(\us23\/_0133_ ), .C_N(\us23\/_0135_ ), .Y(\us23\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us23/_0953_ ( .A(\us23\/_0026_ ), .B(\us23\/_0123_ ), .X(\us23\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0955_ ( .A(\us23\/_0137_ ), .X(\us23\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_0956_ ( .A1(\us23\/_0110_ ), .A2(\us23\/_0293_ ), .A3(\us23\/_0280_ ), .B1(\us23\/_0139_ ), .Y(\us23\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0957_ ( .A(\us23\/_0096_ ), .B(\us23\/_0730_ ), .X(\us23\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0959_ ( .A(\us23\/_0142_ ), .X(\us23\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_0960_ ( .A1(\us23\/_0020_ ), .A2(\us23\/_0144_ ), .A3(\us23\/_0017_ ), .B1(\us23\/_0139_ ), .Y(\us23\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \us23/_0961_ ( .A(\sa23\[2\] ), .B(\us23\/_0050_ ), .C_N(\sa23\[3\] ), .Y(\us23\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0962_ ( .A(\us23\/_0128_ ), .X(\us23\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_0963_ ( .A1(\us23\/_0146_ ), .A2(\us23\/_0032_ ), .A3(\us23\/_0640_ ), .B1(\us23\/_0147_ ), .Y(\us23\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us23/_0964_ ( .A(\us23\/_0136_ ), .B(\us23\/_0141_ ), .C(\us23\/_0145_ ), .D(\us23\/_0148_ ), .X(\us23\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0965_ ( .A(\us23\/_0123_ ), .B(\us23\/_0151_ ), .X(\us23\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0967_ ( .A(\us23\/_0150_ ), .X(\us23\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \us23/_0968_ ( .A(\us23\/_0150_ ), .B(\us23\/_0062_ ), .X(\us23\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_0969_ ( .A(\us23\/_0079_ ), .B(\us23\/_0150_ ), .Y(\us23\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us23/_0970_ ( .A(\us23\/_0150_ ), .B(\us23\/_0423_ ), .C(\us23\/_0543_ ), .Y(\us23\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_0971_ ( .A(\us23\/_0155_ ), .B(\us23\/_0156_ ), .Y(\us23\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_0972_ ( .A1(\us23\/_0153_ ), .A2(\us23\/_0134_ ), .B1(\us23\/_0154_ ), .C1(\us23\/_0157_ ), .Y(\us23\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0973_ ( .A(\us23\/_0467_ ), .B(\us23\/_0123_ ), .X(\us23\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_0975_ ( .A(\us23\/_0159_ ), .X(\us23\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us23/_0976_ ( .A_N(\us23\/_0119_ ), .B(\us23\/_0161_ ), .X(\us23\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us23/_0977_ ( .A(\us23\/_0163_ ), .Y(\us23\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_0978_ ( .A1(\us23\/_0146_ ), .A2(\us23\/_0575_ ), .A3(\us23\/_0608_ ), .B1(\us23\/_0153_ ), .Y(\us23\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_0979_ ( .A1(\us23\/_0062_ ), .A2(\us23\/_0280_ ), .A3(\us23\/_0134_ ), .B1(\us23\/_0161_ ), .Y(\us23\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us23/_0980_ ( .A(\us23\/_0158_ ), .B(\us23\/_0164_ ), .C(\us23\/_0165_ ), .D(\us23\/_0166_ ), .X(\us23\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us23/_0981_ ( .A(\us23\/_0097_ ), .B(\us23\/_0122_ ), .C(\us23\/_0149_ ), .D(\us23\/_0167_ ), .X(\us23\/_0168_ ) );
sky130_fd_sc_hd__and2_1 \us23/_0982_ ( .A(\us23\/_0662_ ), .B(\us23\/_0150_ ), .X(\us23\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_0983_ ( .A(\us23\/_0154_ ), .B(\us23\/_0169_ ), .Y(\us23\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us23/_0984_ ( .A(\us23\/_0123_ ), .B(\us23\/_0151_ ), .C(\us23\/_0038_ ), .X(\us23\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0985_ ( .A(\us23\/_0170_ ), .B(\us23\/_0171_ ), .X(\us23\/_0172_ ) );
sky130_fd_sc_hd__inv_2 \us23/_0986_ ( .A(\us23\/_0172_ ), .Y(\us23\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \us23/_0987_ ( .A(\us23\/_0067_ ), .B(\us23\/_0168_ ), .C(\us23\/_0174_ ), .Y(\us23\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us23/_0988_ ( .A(\sa23\[1\] ), .B(\sa23\[0\] ), .Y(\us23\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us23/_0989_ ( .A(\us23\/_0175_ ), .B(\us23\/_0358_ ), .X(\us23\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0990_ ( .A(\us23\/_0176_ ), .B(\us23\/_0478_ ), .X(\us23\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_0991_ ( .A(\us23\/_0280_ ), .B(\us23\/_0113_ ), .Y(\us23\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0992_ ( .A(\us23\/_0111_ ), .B(\us23\/_0062_ ), .X(\us23\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0993_ ( .A(\us23\/_0111_ ), .B(\us23\/_0662_ ), .X(\us23\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_0994_ ( .A(\us23\/_0179_ ), .B(\us23\/_0180_ ), .Y(\us23\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0995_ ( .A(\us23\/_0054_ ), .B(\us23\/_0058_ ), .X(\us23\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us23/_0996_ ( .A(\us23\/_0182_ ), .Y(\us23\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us23/_0997_ ( .A_N(\us23\/_0177_ ), .B(\us23\/_0178_ ), .C(\us23\/_0181_ ), .D(\us23\/_0184_ ), .X(\us23\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0998_ ( .A(\us23\/_0098_ ), .B(\us23\/_0741_ ), .X(\us23\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us23/_0999_ ( .A(\us23\/_0047_ ), .B(\us23\/_0098_ ), .X(\us23\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us23/_1000_ ( .A(\us23\/_0186_ ), .B(\us23\/_0187_ ), .X(\us23\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1001_ ( .A(\us23\/_0188_ ), .Y(\us23\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1002_ ( .A(\us23\/_0738_ ), .B(\us23\/_0735_ ), .X(\us23\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1003_ ( .A(\us23\/_0271_ ), .B(\us23\/_0736_ ), .X(\us23\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_1004_ ( .A(\us23\/_0190_ ), .B(\us23\/_0191_ ), .Y(\us23\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us23/_1005_ ( .A(\us23\/_0096_ ), .B(\us23\/_0325_ ), .X(\us23\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1006_ ( .A1(\us23\/_0193_ ), .A2(\us23\/_0176_ ), .B1(\us23\/_0043_ ), .Y(\us23\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1007_ ( .A(\us23\/_0185_ ), .B(\us23\/_0189_ ), .C(\us23\/_0192_ ), .D(\us23\/_0195_ ), .X(\us23\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us23/_1008_ ( .A_N(\sa23\[3\] ), .B(\us23\/_0734_ ), .C(\sa23\[2\] ), .X(\us23\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1009_ ( .A(\us23\/_0137_ ), .B(\us23\/_0197_ ), .X(\us23\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_1010_ ( .A(\us23\/_0198_ ), .B(\us23\/_0040_ ), .Y(\us23\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1011_ ( .A(\us23\/_0293_ ), .B(\us23\/_0137_ ), .X(\us23\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1012_ ( .A(\us23\/_0200_ ), .Y(\us23\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1013_ ( .A(\us23\/_0137_ ), .B(\us23\/_0110_ ), .Y(\us23\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1014_ ( .A(\us23\/_0139_ ), .B(\us23\/_0020_ ), .Y(\us23\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1015_ ( .A(\us23\/_0199_ ), .B(\us23\/_0201_ ), .C(\us23\/_0202_ ), .D(\us23\/_0203_ ), .X(\us23\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us23/_1016_ ( .A1(\us23\/_0532_ ), .A2(\us23\/_0109_ ), .B1(\us23\/_0102_ ), .C1(\us23\/_0727_ ), .X(\us23\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1017_ ( .A(\us23\/_0022_ ), .B(\us23\/_0078_ ), .Y(\us23\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1018_ ( .A(\us23\/_0078_ ), .B(\us23\/_0142_ ), .Y(\us23\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1019_ ( .A(\us23\/_0207_ ), .B(\us23\/_0208_ ), .Y(\us23\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1020_ ( .A1(\us23\/_0094_ ), .A2(\us23\/_0176_ ), .B1(\us23\/_0206_ ), .C1(\us23\/_0209_ ), .Y(\us23\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1021_ ( .A(\us23\/_0662_ ), .B(\us23\/_0070_ ), .X(\us23\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us23/_1022_ ( .A(\us23\/_0731_ ), .B(\us23\/_0123_ ), .C(\us23\/_0749_ ), .Y(\us23\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us23/_1023_ ( .A(\us23\/_0731_ ), .B(\us23\/_0467_ ), .C(\us23\/_0069_ ), .Y(\us23\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us23/_1024_ ( .A_N(\us23\/_0211_ ), .B(\us23\/_0127_ ), .C(\us23\/_0212_ ), .D(\us23\/_0213_ ), .X(\us23\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1025_ ( .A(\us23\/_0137_ ), .Y(\us23\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1026_ ( .A(\us23\/_0128_ ), .B(\us23\/_0035_ ), .Y(\us23\/_0217_ ) );
sky130_fd_sc_hd__buf_2 \us23/_1027_ ( .A(\us23\/_0478_ ), .X(\us23\/_0218_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1028_ ( .A1(\us23\/_0159_ ), .A2(\us23\/_0746_ ), .B1(\us23\/_0434_ ), .B2(\us23\/_0218_ ), .Y(\us23\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us23/_1029_ ( .A1(\us23\/_0116_ ), .A2(\us23\/_0215_ ), .B1(\us23\/_0217_ ), .C1(\us23\/_0219_ ), .X(\us23\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1030_ ( .A(\us23\/_0113_ ), .B(\us23\/_0746_ ), .X(\us23\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us23/_1031_ ( .A1(\us23\/_0098_ ), .A2(\us23\/_0746_ ), .B1(\us23\/_0434_ ), .B2(\us23\/_0750_ ), .X(\us23\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1032_ ( .A1(\us23\/_0047_ ), .A2(\us23\/_0113_ ), .B1(\us23\/_0221_ ), .C1(\us23\/_0222_ ), .Y(\us23\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us23/_1033_ ( .A1(\us23\/_0129_ ), .A2(\us23\/_0162_ ), .B1(\us23\/_0271_ ), .B2(\us23\/_0705_ ), .X(\us23\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1034_ ( .A1(\us23\/_0093_ ), .A2(\us23\/_0738_ ), .B1(\us23\/_0081_ ), .C1(\us23\/_0224_ ), .Y(\us23\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1035_ ( .A(\us23\/_0214_ ), .B(\us23\/_0220_ ), .C(\us23\/_0223_ ), .D(\us23\/_0225_ ), .X(\us23\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1036_ ( .A(\us23\/_0196_ ), .B(\us23\/_0204_ ), .C(\us23\/_0210_ ), .D(\us23\/_0226_ ), .X(\us23\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1037_ ( .A(\us23\/_0111_ ), .B(\us23\/_0554_ ), .X(\us23\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1038_ ( .A(\us23\/_0229_ ), .Y(\us23\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1039_ ( .A(\us23\/_0111_ ), .B(\us23\/_0129_ ), .Y(\us23\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1040_ ( .A(\us23\/_0017_ ), .B(\us23\/_0738_ ), .Y(\us23\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1041_ ( .A(\us23\/_0030_ ), .B(\us23\/_0304_ ), .Y(\us23\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1042_ ( .A(\us23\/_0230_ ), .B(\us23\/_0231_ ), .C(\us23\/_0232_ ), .D(\us23\/_0233_ ), .X(\us23\/_0234_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1043_ ( .A(\us23\/_0047_ ), .B(\us23\/_0478_ ), .X(\us23\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1044_ ( .A1(\us23\/_0129_ ), .A2(\us23\/_0554_ ), .B1(\us23\/_0137_ ), .Y(\us23\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us23/_1045_ ( .A(\us23\/_0235_ ), .B(\us23\/_0049_ ), .C_N(\us23\/_0236_ ), .Y(\us23\/_0237_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1046_ ( .A(\us23\/_0047_ ), .B(\us23\/_0077_ ), .X(\us23\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1047_ ( .A(\us23\/_0070_ ), .B(\us23\/_0035_ ), .X(\us23\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us23/_1048_ ( .A1(\us23\/_0047_ ), .A2(\us23\/_0736_ ), .B1(\us23\/_0022_ ), .B2(\us23\/_0099_ ), .X(\us23\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us23/_1049_ ( .A(\us23\/_0239_ ), .B(\us23\/_0240_ ), .C(\us23\/_0241_ ), .Y(\us23\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1050_ ( .A(\us23\/_0554_ ), .B(\us23\/_0072_ ), .X(\us23\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us23/_1051_ ( .A1(\us23\/_0142_ ), .A2(\us23\/_0137_ ), .B1(\us23\/_0159_ ), .B2(\us23\/_0082_ ), .X(\us23\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1052_ ( .A1(\us23\/_0608_ ), .A2(\us23\/_0072_ ), .B1(\us23\/_0243_ ), .C1(\us23\/_0244_ ), .Y(\us23\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1053_ ( .A(\us23\/_0234_ ), .B(\us23\/_0237_ ), .C(\us23\/_0242_ ), .D(\us23\/_0245_ ), .X(\us23\/_0246_ ) );
sky130_fd_sc_hd__buf_2 \us23/_1054_ ( .A(\us23\/_0027_ ), .X(\us23\/_0247_ ) );
sky130_fd_sc_hd__o21a_1 \us23/_1055_ ( .A1(\us23\/_0554_ ), .A2(\us23\/_0586_ ), .B1(\us23\/_0247_ ), .X(\us23\/_0248_ ) );
sky130_fd_sc_hd__and2_1 \us23/_1056_ ( .A(\us23\/_0082_ ), .B(\us23\/_0478_ ), .X(\us23\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_1057_ ( .A(\us23\/_0079_ ), .X(\us23\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1058_ ( .A(\us23\/_0251_ ), .B(\us23\/_0478_ ), .X(\us23\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_1059_ ( .A(\us23\/_0250_ ), .B(\us23\/_0252_ ), .Y(\us23\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1060_ ( .A(\us23\/_0016_ ), .B(\us23\/_0064_ ), .Y(\us23\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_1061_ ( .A(\us23\/_0304_ ), .X(\us23\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1062_ ( .A(\us23\/_0255_ ), .B(\us23\/_0640_ ), .Y(\us23\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us23/_1063_ ( .A_N(\us23\/_0248_ ), .B(\us23\/_0253_ ), .C(\us23\/_0254_ ), .D(\us23\/_0256_ ), .X(\us23\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1064_ ( .A(\us23\/_0099_ ), .B(\us23\/_0110_ ), .X(\us23\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us23/_1065_ ( .A1(\us23\/_0161_ ), .A2(\us23\/_0130_ ), .B1(\us23\/_0258_ ), .Y(\us23\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1066_ ( .A(\us23\/_0194_ ), .B(\sa23\[1\] ), .X(\us23\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1068_ ( .A(\us23\/_0261_ ), .B(\us23\/_0153_ ), .Y(\us23\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us23/_1069_ ( .A_N(\us23\/_0154_ ), .B(\us23\/_0259_ ), .C(\us23\/_0263_ ), .X(\us23\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1070_ ( .A(\us23\/_0246_ ), .B(\us23\/_0174_ ), .C(\us23\/_0257_ ), .D(\us23\/_0264_ ), .X(\us23\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us23/_1071_ ( .A1(\us23\/_0261_ ), .A2(\us23\/_0554_ ), .B1(\us23\/_0159_ ), .X(\us23\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1072_ ( .A(\us23\/_0746_ ), .B(\us23\/_0150_ ), .Y(\us23\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1073_ ( .A(\us23\/_0175_ ), .Y(\us23\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us23/_1074_ ( .A(\us23\/_0423_ ), .B(\us23\/_0123_ ), .C(\us23\/_0151_ ), .X(\us23\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1075_ ( .A(\us23\/_0268_ ), .B(\us23\/_0269_ ), .Y(\us23\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us23/_1076_ ( .A_N(\us23\/_0266_ ), .B(\us23\/_0267_ ), .C(\us23\/_0270_ ), .X(\us23\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1077_ ( .A(\us23\/_0554_ ), .B(\us23\/_0150_ ), .X(\us23\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1078_ ( .A(\us23\/_0273_ ), .Y(\us23\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1079_ ( .A1(\us23\/_0734_ ), .A2(\us23\/_0325_ ), .B1(\us23\/_0380_ ), .Y(\us23\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1080_ ( .A(\us23\/_0275_ ), .Y(\us23\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1081_ ( .A(\us23\/_0276_ ), .B(\us23\/_0153_ ), .Y(\us23\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us23/_1082_ ( .A(\us23\/_0272_ ), .B(\us23\/_0274_ ), .C(\us23\/_0277_ ), .X(\us23\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_1083_ ( .A(\us23\/_0035_ ), .X(\us23\/_0279_ ) );
sky130_fd_sc_hd__buf_2 \us23/_1084_ ( .A(\us23\/_0082_ ), .X(\us23\/_0280_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1085_ ( .A1(\us23\/_0218_ ), .A2(\us23\/_0279_ ), .B1(\us23\/_0280_ ), .B2(\us23\/_0060_ ), .Y(\us23\/_0281_ ) );
sky130_fd_sc_hd__o21ai_1 \us23/_1086_ ( .A1(\us23\/_0251_ ), .A2(\us23\/_0434_ ), .B1(\us23\/_0304_ ), .Y(\us23\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1087_ ( .A(\us23\/_0091_ ), .B(\us23\/_0056_ ), .Y(\us23\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1088_ ( .A1(\us23\/_0118_ ), .A2(\us23\/_0050_ ), .B1(\us23\/_0038_ ), .C1(\us23\/_0255_ ), .Y(\us23\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1089_ ( .A(\us23\/_0281_ ), .B(\us23\/_0283_ ), .C(\us23\/_0284_ ), .D(\us23\/_0285_ ), .X(\us23\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1090_ ( .A(\us23\/_0082_ ), .B(\us23\/_0027_ ), .X(\us23\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1091_ ( .A(\us23\/_0129_ ), .B(\us23\/_0027_ ), .X(\us23\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_1092_ ( .A(\us23\/_0287_ ), .B(\us23\/_0288_ ), .Y(\us23\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1093_ ( .A1(\us23\/_0752_ ), .A2(\us23\/_0683_ ), .B1(\us23\/_0093_ ), .B2(\us23\/_0247_ ), .Y(\us23\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1094_ ( .A1(\us23\/_0092_ ), .A2(\us23\/_0575_ ), .B1(\us23\/_0056_ ), .Y(\us23\/_0291_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1096_ ( .A1(\us23\/_0218_ ), .A2(\us23\/_0662_ ), .B1(\us23\/_0280_ ), .B2(\us23\/_0056_ ), .Y(\us23\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1097_ ( .A(\us23\/_0289_ ), .B(\us23\/_0290_ ), .C(\us23\/_0291_ ), .D(\us23\/_0294_ ), .X(\us23\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1098_ ( .A(\us23\/_0750_ ), .B(\us23\/_0193_ ), .X(\us23\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1099_ ( .A(\us23\/_0705_ ), .B(\us23\/_0380_ ), .X(\us23\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1100_ ( .A(\us23\/_0752_ ), .B(\us23\/_0129_ ), .Y(\us23\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us23/_1101_ ( .A(\us23\/_0296_ ), .B(\us23\/_0297_ ), .C_N(\us23\/_0298_ ), .Y(\us23\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1102_ ( .A(\us23\/_0089_ ), .B(\us23\/_0532_ ), .Y(\us23\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1103_ ( .A(\sa23\[2\] ), .Y(\us23\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \us23/_1104_ ( .A(\us23\/_0301_ ), .B(\sa23\[3\] ), .C(\us23\/_0118_ ), .Y(\us23\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1105_ ( .A(\us23\/_0072_ ), .B(\us23\/_0302_ ), .X(\us23\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1106_ ( .A(\us23\/_0303_ ), .Y(\us23\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1107_ ( .A(\us23\/_0147_ ), .B(\us23\/_0302_ ), .Y(\us23\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1108_ ( .A(\us23\/_0299_ ), .B(\us23\/_0300_ ), .C(\us23\/_0305_ ), .D(\us23\/_0306_ ), .X(\us23\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1109_ ( .A(\us23\/_0278_ ), .B(\us23\/_0286_ ), .C(\us23\/_0295_ ), .D(\us23\/_0307_ ), .X(\us23\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us23/_1110_ ( .A(\us23\/_0228_ ), .B(\us23\/_0265_ ), .C(\us23\/_0308_ ), .Y(\us23\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1111_ ( .A(\us23\/_0235_ ), .Y(\us23\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1112_ ( .A(\us23\/_0478_ ), .B(\us23\/_0640_ ), .X(\us23\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1113_ ( .A(\us23\/_0310_ ), .Y(\us23\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1114_ ( .A(\us23\/_0022_ ), .B(\us23\/_0218_ ), .Y(\us23\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1115_ ( .A(\us23\/_0218_ ), .B(\us23\/_0032_ ), .Y(\us23\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1116_ ( .A(\us23\/_0309_ ), .B(\us23\/_0311_ ), .C(\us23\/_0312_ ), .D(\us23\/_0313_ ), .X(\us23\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1117_ ( .A(\us23\/_0218_ ), .B(\us23\/_0064_ ), .Y(\us23\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1118_ ( .A(\us23\/_0218_ ), .B(\us23\/_0683_ ), .Y(\us23\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1119_ ( .A(\us23\/_0315_ ), .B(\us23\/_0316_ ), .C(\us23\/_0317_ ), .D(\us23\/_0253_ ), .X(\us23\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1120_ ( .A(\us23\/_0047_ ), .B(\us23\/_0304_ ), .Y(\us23\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1121_ ( .A(\us23\/_0586_ ), .B(\us23\/_0162_ ), .Y(\us23\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1122_ ( .A(\us23\/_0319_ ), .B(\us23\/_0320_ ), .Y(\us23\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_1123_ ( .A(\us23\/_0321_ ), .B(\us23\/_0238_ ), .Y(\us23\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1124_ ( .A(\us23\/_0304_ ), .B(\us23\/_0062_ ), .Y(\us23\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_1125_ ( .A(\us23\/_0251_ ), .X(\us23\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1126_ ( .A1(\us23\/_0324_ ), .A2(\us23\/_0280_ ), .B1(\us23\/_0255_ ), .Y(\us23\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1127_ ( .A1(\us23\/_0050_ ), .A2(\us23\/_0205_ ), .B1(\us23\/_0109_ ), .C1(\us23\/_0255_ ), .Y(\us23\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1128_ ( .A(\us23\/_0322_ ), .B(\us23\/_0323_ ), .C(\us23\/_0326_ ), .D(\us23\/_0327_ ), .X(\us23\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1129_ ( .A1(\us23\/_0733_ ), .A2(\us23\/_0279_ ), .A3(\us23\/_0058_ ), .B1(\us23\/_0056_ ), .Y(\us23\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_1130_ ( .A(\us23\/_0047_ ), .X(\us23\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1131_ ( .A(\us23\/_0330_ ), .B(\us23\/_0056_ ), .Y(\us23\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1132_ ( .A(\us23\/_0054_ ), .B(\us23\/_0045_ ), .Y(\us23\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1133_ ( .A(\us23\/_0329_ ), .B(\us23\/_0331_ ), .C(\us23\/_0284_ ), .D(\us23\/_0332_ ), .X(\us23\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us23/_1134_ ( .A1(\us23\/_0543_ ), .A2(\us23\/_0205_ ), .B1(\us23\/_0532_ ), .C1(\us23\/_0060_ ), .X(\us23\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1135_ ( .A(\us23\/_0280_ ), .B(\us23\/_0060_ ), .Y(\us23\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1136_ ( .A(\us23\/_0324_ ), .B(\us23\/_0060_ ), .Y(\us23\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1137_ ( .A(\us23\/_0335_ ), .B(\us23\/_0337_ ), .Y(\us23\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1138_ ( .A1(\us23\/_0276_ ), .A2(\us23\/_0060_ ), .B1(\us23\/_0334_ ), .C1(\us23\/_0338_ ), .Y(\us23\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1139_ ( .A(\us23\/_0318_ ), .B(\us23\/_0328_ ), .C(\us23\/_0333_ ), .D(\us23\/_0339_ ), .X(\us23\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us23/_1140_ ( .A1(\us23\/_0746_ ), .A2(\us23\/_0134_ ), .B1(\us23\/_0128_ ), .X(\us23\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us23/_1141_ ( .A_N(\us23\/_0086_ ), .B(\us23\/_0128_ ), .X(\us23\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1142_ ( .A(\us23\/_0079_ ), .B(\us23\/_0124_ ), .X(\us23\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_1143_ ( .A(\us23\/_0126_ ), .B(\us23\/_0343_ ), .Y(\us23\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us23/_1144_ ( .A(\us23\/_0341_ ), .B(\us23\/_0342_ ), .C_N(\us23\/_0344_ ), .Y(\us23\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1146_ ( .A1(\us23\/_0193_ ), .A2(\us23\/_0092_ ), .A3(\us23\/_0330_ ), .B1(\us23\/_0147_ ), .Y(\us23\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1147_ ( .A1(\us23\/_0130_ ), .A2(\us23\/_0280_ ), .A3(\us23\/_0134_ ), .B1(\us23\/_0139_ ), .Y(\us23\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1148_ ( .A1(\us23\/_0144_ ), .A2(\us23\/_0608_ ), .A3(\us23\/_0092_ ), .B1(\us23\/_0139_ ), .Y(\us23\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1149_ ( .A(\us23\/_0345_ ), .B(\us23\/_0348_ ), .C(\us23\/_0349_ ), .D(\us23\/_0350_ ), .X(\us23\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us23/_1150_ ( .A(\us23\/_0150_ ), .B(\us23\/_0194_ ), .C(\us23\/_0543_ ), .X(\us23\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us23/_1151_ ( .A(\us23\/_0277_ ), .SLEEP(\us23\/_0352_ ), .X(\us23\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us23/_1152_ ( .A1(\us23\/_0268_ ), .A2(\us23\/_0171_ ), .B1(\us23\/_0157_ ), .Y(\us23\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us23/_1153_ ( .A(\us23\/_0161_ ), .X(\us23\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1154_ ( .A1(\us23\/_0279_ ), .A2(\us23\/_0280_ ), .B1(\us23\/_0355_ ), .Y(\us23\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1155_ ( .A1(\us23\/_0020_ ), .A2(\us23\/_0193_ ), .A3(\us23\/_0091_ ), .B1(\us23\/_0355_ ), .Y(\us23\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1156_ ( .A(\us23\/_0353_ ), .B(\us23\/_0354_ ), .C(\us23\/_0356_ ), .D(\us23\/_0357_ ), .X(\us23\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1157_ ( .A(\us23\/_0111_ ), .B(\us23\/_0586_ ), .X(\us23\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1158_ ( .A(\us23\/_0360_ ), .Y(\us23\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us23/_1159_ ( .A1(\us23\/_0119_ ), .A2(\us23\/_0120_ ), .B1(\us23\/_0230_ ), .C1(\us23\/_0361_ ), .X(\us23\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1160_ ( .A1(\us23\/_0662_ ), .A2(\us23\/_0251_ ), .A3(\us23\/_0134_ ), .B1(\us23\/_0114_ ), .Y(\us23\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1162_ ( .A1(\us23\/_0035_ ), .A2(\us23\/_0251_ ), .A3(\us23\/_0134_ ), .B1(\us23\/_0099_ ), .Y(\us23\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1163_ ( .A1(\us23\/_0193_ ), .A2(\us23\/_0608_ ), .B1(\us23\/_0099_ ), .Y(\us23\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1164_ ( .A(\us23\/_0362_ ), .B(\us23\/_0363_ ), .C(\us23\/_0365_ ), .D(\us23\/_0366_ ), .X(\us23\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1165_ ( .A1(\us23\/_0575_ ), .A2(\us23\/_0092_ ), .A3(\us23\/_0330_ ), .B1(\us23\/_0089_ ), .Y(\us23\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1166_ ( .A1(\us23\/_0586_ ), .A2(\us23\/_0017_ ), .A3(\us23\/_0330_ ), .B1(\us23\/_0094_ ), .Y(\us23\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \us23/_1167_ ( .A1(\us23\/_0293_ ), .A2(\us23\/_0134_ ), .B1(\us23\/_0089_ ), .Y(\us23\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1168_ ( .A1(\us23\/_0279_ ), .A2(\us23\/_0134_ ), .B1(\us23\/_0094_ ), .Y(\us23\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1169_ ( .A(\us23\/_0368_ ), .B(\us23\/_0370_ ), .C(\us23\/_0371_ ), .D(\us23\/_0372_ ), .X(\us23\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1170_ ( .A(\us23\/_0351_ ), .B(\us23\/_0359_ ), .C(\us23\/_0367_ ), .D(\us23\/_0373_ ), .X(\us23\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1171_ ( .A1(\us23\/_0102_ ), .A2(\us23\/_0347_ ), .B1(\us23\/_0109_ ), .C1(\us23\/_0247_ ), .Y(\us23\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1172_ ( .A1(\us23\/_0102_ ), .A2(\us23\/_0347_ ), .B1(\us23\/_0532_ ), .C1(\us23\/_0247_ ), .Y(\us23\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1173_ ( .A1(\us23\/_0050_ ), .A2(\us23\/_0543_ ), .B1(\us23\/_0380_ ), .C1(\us23\/_0247_ ), .Y(\us23\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1174_ ( .A(\us23\/_0041_ ), .B(\us23\/_0375_ ), .C(\us23\/_0376_ ), .D(\us23\/_0377_ ), .X(\us23\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1175_ ( .A(\us23\/_0047_ ), .B(\us23\/_0750_ ), .X(\us23\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1176_ ( .A(\us23\/_0379_ ), .Y(\us23\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1177_ ( .A(\us23\/_0016_ ), .B(\us23\/_0608_ ), .Y(\us23\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1178_ ( .A(\us23\/_0752_ ), .B(\us23\/_0554_ ), .Y(\us23\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1179_ ( .A1(\sa23\[1\] ), .A2(\us23\/_0734_ ), .B1(\us23\/_0109_ ), .C1(\us23\/_0016_ ), .Y(\us23\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1180_ ( .A(\us23\/_0381_ ), .B(\us23\/_0382_ ), .C(\us23\/_0383_ ), .D(\us23\/_0384_ ), .X(\us23\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us23/_1181_ ( .A(\us23\/_0086_ ), .B_N(\us23\/_0736_ ), .X(\us23\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1182_ ( .A1(\us23\/_0748_ ), .A2(\us23\/_0134_ ), .B1(\us23\/_0739_ ), .Y(\us23\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1183_ ( .A1(\us23\/_0118_ ), .A2(\us23\/_0543_ ), .B1(\us23\/_0109_ ), .C1(\us23\/_0739_ ), .Y(\us23\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1184_ ( .A1(\us23\/_0102_ ), .A2(\us23\/_0301_ ), .B1(\sa23\[3\] ), .C1(\us23\/_0739_ ), .Y(\us23\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1185_ ( .A(\us23\/_0386_ ), .B(\us23\/_0387_ ), .C(\us23\/_0388_ ), .D(\us23\/_0389_ ), .X(\us23\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1186_ ( .A(\us23\/_0020_ ), .Y(\us23\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1187_ ( .A(\us23\/_0727_ ), .Y(\us23\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1188_ ( .A(\us23\/_0727_ ), .B(\us23\/_0064_ ), .Y(\us23\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1189_ ( .A1(\us23\/_0102_ ), .A2(\us23\/_0734_ ), .B1(\us23\/_0532_ ), .C1(\us23\/_0727_ ), .Y(\us23\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us23/_1190_ ( .A1(\us23\/_0392_ ), .A2(\us23\/_0393_ ), .B1(\us23\/_0394_ ), .C1(\us23\/_0395_ ), .X(\us23\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1191_ ( .A(\us23\/_0378_ ), .B(\us23\/_0385_ ), .C(\us23\/_0390_ ), .D(\us23\/_0396_ ), .X(\us23\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us23/_1192_ ( .A(\us23\/_0340_ ), .B(\us23\/_0374_ ), .C(\us23\/_0397_ ), .Y(\us23\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1193_ ( .A(\us23\/_0077_ ), .B(\us23\/_0129_ ), .X(\us23\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_1194_ ( .A(\us23\/_0398_ ), .B(\us23\/_0239_ ), .Y(\us23\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1195_ ( .A(\us23\/_0022_ ), .B(\us23\/_0111_ ), .X(\us23\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us23/_1196_ ( .A_N(\us23\/_0400_ ), .B(\us23\/_0231_ ), .Y(\us23\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us23/_1197_ ( .A(\us23\/_0399_ ), .SLEEP(\us23\/_0402_ ), .X(\us23\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_1198_ ( .A(\us23\/_0746_ ), .B(\us23\/_0251_ ), .Y(\us23\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us23/_1199_ ( .A_N(\us23\/_0404_ ), .B(\us23\/_0752_ ), .Y(\us23\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us23/_1200_ ( .A(\us23\/_0467_ ), .B(\us23\/_0194_ ), .C(\us23\/_0694_ ), .X(\us23\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us23/_1201_ ( .A_N(\us23\/_0175_ ), .B(\us23\/_0406_ ), .X(\us23\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1202_ ( .A(\us23\/_0407_ ), .Y(\us23\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1203_ ( .A1(\us23\/_0094_ ), .A2(\us23\/_0197_ ), .B1(\us23\/_0114_ ), .B2(\us23\/_0640_ ), .Y(\us23\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1204_ ( .A(\us23\/_0403_ ), .B(\us23\/_0405_ ), .C(\us23\/_0408_ ), .D(\us23\/_0409_ ), .X(\us23\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1205_ ( .A(\us23\/_0030_ ), .B(\us23\/_0150_ ), .Y(\us23\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us23/_1206_ ( .A_N(\us23\/_0169_ ), .B(\us23\/_0289_ ), .C(\us23\/_0411_ ), .X(\us23\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us23/_1207_ ( .A1(\us23\/_0467_ ), .A2(\us23\/_0151_ ), .B1(\us23\/_0140_ ), .C1(\us23\/_0129_ ), .X(\us23\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1208_ ( .A1(\us23\/_0608_ ), .A2(\us23\/_0099_ ), .B1(\us23\/_0037_ ), .C1(\us23\/_0414_ ), .Y(\us23\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1209_ ( .A(\us23\/_0738_ ), .Y(\us23\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1210_ ( .A(\us23\/_0586_ ), .B(\us23\/_0736_ ), .Y(\us23\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1211_ ( .A1(\us23\/_0194_ ), .A2(\us23\/_0038_ ), .B1(\us23\/_0118_ ), .C1(\us23\/_0153_ ), .Y(\us23\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us23/_1212_ ( .A1(\us23\/_0416_ ), .A2(\us23\/_0117_ ), .B1(\us23\/_0417_ ), .C1(\us23\/_0418_ ), .X(\us23\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1213_ ( .A(\us23\/_0077_ ), .B(\us23\/_0035_ ), .X(\us23\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1214_ ( .A(\us23\/_0662_ ), .B(\us23\/_0124_ ), .Y(\us23\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1215_ ( .A(\us23\/_0030_ ), .B(\us23\/_0137_ ), .Y(\us23\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1216_ ( .A(\us23\/_0072_ ), .B(\us23\/_0731_ ), .Y(\us23\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us23/_1217_ ( .A_N(\us23\/_0420_ ), .B(\us23\/_0421_ ), .C(\us23\/_0422_ ), .D(\us23\/_0424_ ), .X(\us23\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1218_ ( .A(\us23\/_0413_ ), .B(\us23\/_0415_ ), .C(\us23\/_0419_ ), .D(\us23\/_0425_ ), .X(\us23\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us23/_1219_ ( .A(\us23\/_0355_ ), .B(\us23\/_0102_ ), .C(\us23\/_0109_ ), .Y(\us23\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1220_ ( .A(\us23\/_0077_ ), .B(\us23\/_0017_ ), .X(\us23\/_0428_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1221_ ( .A(\us23\/_0077_ ), .B(\us23\/_0554_ ), .X(\us23\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us23/_1222_ ( .A1(\us23\/_0050_ ), .A2(\us23\/_0205_ ), .B1(\us23\/_0380_ ), .C1(\us23\/_0078_ ), .X(\us23\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us23/_1223_ ( .A(\us23\/_0428_ ), .B(\us23\/_0429_ ), .C(\us23\/_0430_ ), .Y(\us23\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us23/_1224_ ( .A_N(\us23\/_0209_ ), .B(\us23\/_0431_ ), .X(\us23\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us23/_1225_ ( .A1(\us23\/_0215_ ), .A2(\us23\/_0404_ ), .B1(\us23\/_0427_ ), .C1(\us23\/_0432_ ), .X(\us23\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1226_ ( .A(\us23\/_0043_ ), .B(\us23\/_0058_ ), .Y(\us23\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1227_ ( .A(\us23\/_0195_ ), .B(\us23\/_0233_ ), .C(\us23\/_0320_ ), .D(\us23\/_0435_ ), .X(\us23\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1228_ ( .A(\us23\/_0261_ ), .B(\us23\/_0738_ ), .Y(\us23\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1229_ ( .A1(\us23\/_0218_ ), .A2(\us23\/_0640_ ), .B1(\us23\/_0261_ ), .B2(\us23\/_0056_ ), .Y(\us23\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1230_ ( .A(\us23\/_0436_ ), .B(\us23\/_0394_ ), .C(\us23\/_0437_ ), .D(\us23\/_0438_ ), .X(\us23\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1231_ ( .A(\us23\/_0410_ ), .B(\us23\/_0426_ ), .C(\us23\/_0433_ ), .D(\us23\/_0439_ ), .X(\us23\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us23/_1232_ ( .A(\us23\/_0135_ ), .SLEEP(\us23\/_0273_ ), .X(\us23\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1233_ ( .A1(\us23\/_0279_ ), .A2(\us23\/_0134_ ), .B1(\us23\/_0099_ ), .Y(\us23\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1234_ ( .A(\us23\/_0441_ ), .B(\us23\/_0164_ ), .C(\us23\/_0270_ ), .D(\us23\/_0442_ ), .X(\us23\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1235_ ( .A(\us23\/_0051_ ), .B(\us23\/_0662_ ), .Y(\us23\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1236_ ( .A(\us23\/_0051_ ), .B(\us23\/_0271_ ), .Y(\us23\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1237_ ( .A(\us23\/_0444_ ), .B(\us23\/_0446_ ), .X(\us23\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1238_ ( .A(\us23\/_0193_ ), .B(\us23\/_0304_ ), .X(\us23\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1239_ ( .A(\us23\/_0448_ ), .Y(\us23\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1240_ ( .A(\us23\/_0162_ ), .B(\us23\/_0130_ ), .X(\us23\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1241_ ( .A(\us23\/_0450_ ), .Y(\us23\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1242_ ( .A1(\us23\/_0129_ ), .A2(\us23\/_0554_ ), .B1(\us23\/_0043_ ), .Y(\us23\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1243_ ( .A(\us23\/_0447_ ), .B(\us23\/_0449_ ), .C(\us23\/_0451_ ), .D(\us23\/_0452_ ), .X(\us23\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1244_ ( .A(\us23\/_0056_ ), .B(\us23\/_0064_ ), .Y(\us23\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us23/_1245_ ( .A_N(\us23\/_0248_ ), .B(\us23\/_0454_ ), .C(\us23\/_0254_ ), .D(\us23\/_0256_ ), .X(\us23\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1246_ ( .A1(\us23\/_0330_ ), .A2(\us23\/_0099_ ), .B1(\us23\/_0134_ ), .B2(\us23\/_0705_ ), .Y(\us23\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1247_ ( .A1(\us23\/_0748_ ), .A2(\us23\/_0738_ ), .B1(\us23\/_0092_ ), .B2(\us23\/_0752_ ), .Y(\us23\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1248_ ( .A1(\us23\/_0072_ ), .A2(\us23\/_0035_ ), .B1(\us23\/_0748_ ), .B2(\us23\/_0056_ ), .Y(\us23\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1249_ ( .A1(\us23\/_0748_ ), .A2(\us23\/_0251_ ), .B1(\us23\/_0247_ ), .Y(\us23\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1250_ ( .A(\us23\/_0457_ ), .B(\us23\/_0458_ ), .C(\us23\/_0459_ ), .D(\us23\/_0460_ ), .X(\us23\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1251_ ( .A(\us23\/_0443_ ), .B(\us23\/_0453_ ), .C(\us23\/_0455_ ), .D(\us23\/_0461_ ), .X(\us23\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1252_ ( .A(\us23\/_0705_ ), .B(\us23\/_0079_ ), .X(\us23\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1253_ ( .A(\us23\/_0586_ ), .B(\us23\/_0124_ ), .Y(\us23\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1254_ ( .A(\us23\/_0218_ ), .B(\us23\/_0746_ ), .Y(\us23\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us23/_1255_ ( .A_N(\us23\/_0463_ ), .B(\us23\/_0464_ ), .C(\us23\/_0465_ ), .X(\us23\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us23/_1256_ ( .A1(\us23\/_0271_ ), .A2(\us23\/_0072_ ), .B1(\us23\/_0142_ ), .B2(\us23\/_0027_ ), .X(\us23\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1257_ ( .A1(\us23\/_0144_ ), .A2(\us23\/_0099_ ), .B1(\us23\/_0360_ ), .C1(\us23\/_0468_ ), .Y(\us23\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us23/_1258_ ( .A1(\us23\/_0662_ ), .A2(\us23\/_0251_ ), .B1(\us23\/_0218_ ), .X(\us23\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1259_ ( .A1(\us23\/_0575_ ), .A2(\us23\/_0056_ ), .B1(\us23\/_0379_ ), .C1(\us23\/_0470_ ), .Y(\us23\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1260_ ( .A(\us23\/_0466_ ), .B(\us23\/_0469_ ), .C(\us23\/_0471_ ), .D(\us23\/_0305_ ), .X(\us23\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us23/_1261_ ( .A1(\us23\/_0247_ ), .A2(\us23\/_0683_ ), .B1(\us23\/_0324_ ), .B2(\us23\/_0056_ ), .X(\us23\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1262_ ( .A(\us23\/_0280_ ), .B(\us23\/_0099_ ), .X(\us23\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us23/_1263_ ( .A1(\us23\/_0092_ ), .A2(\us23\/_0247_ ), .B1(\us23\/_0474_ ), .X(\us23\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us23/_1264_ ( .A(\us23\/_0075_ ), .B(\us23\/_0473_ ), .C(\us23\/_0475_ ), .Y(\us23\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1265_ ( .A1(\us23\/_0279_ ), .A2(\us23\/_0255_ ), .B1(\us23\/_0280_ ), .B2(\us23\/_0060_ ), .Y(\us23\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1266_ ( .A1(\us23\/_0093_ ), .A2(\us23\/_0056_ ), .B1(\us23\/_0134_ ), .B2(\us23\/_0114_ ), .Y(\us23\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1267_ ( .A1(\us23\/_0161_ ), .A2(\us23\/_0032_ ), .B1(\us23\/_0324_ ), .B2(\us23\/_0147_ ), .Y(\us23\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1268_ ( .A1(\us23\/_0054_ ), .A2(\us23\/_0731_ ), .B1(\us23\/_0748_ ), .B2(\us23\/_0304_ ), .Y(\us23\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1269_ ( .A(\us23\/_0477_ ), .B(\us23\/_0479_ ), .C(\us23\/_0480_ ), .D(\us23\/_0481_ ), .X(\us23\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1270_ ( .A(\us23\/_0161_ ), .B(\us23\/_0064_ ), .Y(\us23\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us23/_1271_ ( .A(\us23\/_0731_ ), .B(\us23\/_0123_ ), .C(\us23\/_0467_ ), .Y(\us23\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1272_ ( .A(\us23\/_0483_ ), .B(\us23\/_0484_ ), .Y(\us23\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1273_ ( .A(\us23\/_0297_ ), .Y(\us23\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us23/_1274_ ( .A_N(\us23\/_0485_ ), .B(\us23\/_0181_ ), .C(\us23\/_0486_ ), .D(\us23\/_0386_ ), .X(\us23\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1275_ ( .A(\us23\/_0472_ ), .B(\us23\/_0476_ ), .C(\us23\/_0482_ ), .D(\us23\/_0487_ ), .X(\us23\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \us23/_1276_ ( .A(\us23\/_0440_ ), .B(\us23\/_0462_ ), .C(\us23\/_0488_ ), .Y(\us23\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1277_ ( .A(\us23\/_0403_ ), .B(\us23\/_0230_ ), .C(\us23\/_0451_ ), .D(\us23\/_0361_ ), .X(\us23\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1278_ ( .A1(\us23\/_0118_ ), .A2(\us23\/_0050_ ), .B1(\us23\/_0109_ ), .C1(\us23\/_0139_ ), .Y(\us23\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1279_ ( .A(\us23\/_0447_ ), .B(\us23\/_0437_ ), .C(\us23\/_0491_ ), .D(\us23\/_0427_ ), .X(\us23\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1280_ ( .A1(\us23\/_0280_ ), .A2(\us23\/_0255_ ), .B1(\us23\/_0608_ ), .B2(\us23\/_0247_ ), .Y(\us23\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1281_ ( .A1(\us23\/_0144_ ), .A2(\us23\/_0147_ ), .B1(\us23\/_0355_ ), .B2(\us23\/_0093_ ), .Y(\us23\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1282_ ( .A1(\us23\/_0705_ ), .A2(\us23\/_0279_ ), .B1(\us23\/_0330_ ), .B2(\us23\/_0247_ ), .Y(\us23\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1283_ ( .A1(\us23\/_0279_ ), .A2(\us23\/_0280_ ), .B1(\us23\/_0114_ ), .Y(\us23\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1284_ ( .A(\us23\/_0493_ ), .B(\us23\/_0494_ ), .C(\us23\/_0495_ ), .D(\us23\/_0496_ ), .X(\us23\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1285_ ( .A1(\us23\/_0134_ ), .A2(\us23\/_0137_ ), .B1(\us23\/_0355_ ), .B2(\us23\/_0575_ ), .Y(\us23\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1286_ ( .A1(\us23\/_0099_ ), .A2(\us23\/_0733_ ), .B1(\us23\/_0093_ ), .B2(\us23\/_0218_ ), .Y(\us23\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1287_ ( .A(\us23\/_0147_ ), .B(\us23\/_0640_ ), .Y(\us23\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1288_ ( .A1(\us23\/_0153_ ), .A2(\us23\/_0056_ ), .B1(\us23\/_0748_ ), .Y(\us23\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1289_ ( .A(\us23\/_0498_ ), .B(\us23\/_0500_ ), .C(\us23\/_0501_ ), .D(\us23\/_0502_ ), .X(\us23\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1290_ ( .A(\us23\/_0490_ ), .B(\us23\/_0492_ ), .C(\us23\/_0497_ ), .D(\us23\/_0503_ ), .X(\us23\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us23/_1291_ ( .A_N(\us23\/_0275_ ), .B(\us23\/_0705_ ), .X(\us23\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1292_ ( .A(\us23\/_0505_ ), .Y(\us23\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1293_ ( .A(\us23\/_0380_ ), .B(\us23\/_0347_ ), .X(\us23\/_0507_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1294_ ( .A1(\us23\/_0507_ ), .A2(\us23\/_0093_ ), .B1(\us23\/_0056_ ), .Y(\us23\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1295_ ( .A(\us23\/_0322_ ), .B(\us23\/_0277_ ), .C(\us23\/_0506_ ), .D(\us23\/_0508_ ), .X(\us23\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1296_ ( .A(\us23\/_0280_ ), .B(\us23\/_0705_ ), .X(\us23\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1297_ ( .A1(\us23\/_0733_ ), .A2(\us23\/_0114_ ), .B1(\us23\/_0429_ ), .C1(\us23\/_0511_ ), .Y(\us23\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_1298_ ( .A(\us23\/_0019_ ), .B(\us23\/_0024_ ), .Y(\us23\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1299_ ( .A(\us23\/_0512_ ), .B(\us23\/_0513_ ), .C(\us23\/_0742_ ), .D(\us23\/_0306_ ), .X(\us23\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1300_ ( .A1(\us23\/_0532_ ), .A2(\us23\/_0089_ ), .B1(\us23\/_0154_ ), .C1(\us23\/_0169_ ), .Y(\us23\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us23/_1301_ ( .A1(\us23\/_0749_ ), .A2(\us23\/_0026_ ), .B1(\us23\/_0069_ ), .C1(\us23\/_0032_ ), .X(\us23\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us23/_1302_ ( .A1(\us23\/_0324_ ), .A2(\us23\/_0355_ ), .B1(\us23\/_0330_ ), .B2(\us23\/_0727_ ), .X(\us23\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us23/_1303_ ( .A(\us23\/_0133_ ), .B(\us23\/_0516_ ), .C(\us23\/_0517_ ), .Y(\us23\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1304_ ( .A(\us23\/_0509_ ), .B(\us23\/_0514_ ), .C(\us23\/_0515_ ), .D(\us23\/_0518_ ), .X(\us23\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1305_ ( .A(\us23\/_0746_ ), .B(\us23\/_0072_ ), .Y(\us23\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1306_ ( .A1(\us23\/_0082_ ), .A2(\us23\/_0070_ ), .B1(\us23\/_0043_ ), .B2(\us23\/_0193_ ), .Y(\us23\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1307_ ( .A(\us23\/_0311_ ), .B(\us23\/_0520_ ), .C(\us23\/_0332_ ), .D(\us23\/_0522_ ), .X(\us23\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1308_ ( .A(\us23\/_0129_ ), .B(\us23\/_0218_ ), .X(\us23\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_1309_ ( .A(\us23\/_0235_ ), .B(\us23\/_0524_ ), .Y(\us23\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us23/_1310_ ( .A(\us23\/_0081_ ), .B(\us23\/_0085_ ), .Y(\us23\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1311_ ( .A1(\us23\/_0051_ ), .A2(\us23\/_0045_ ), .B1(\us23\/_0130_ ), .B2(\us23\/_0094_ ), .Y(\us23\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1312_ ( .A(\us23\/_0523_ ), .B(\us23\/_0525_ ), .C(\us23\/_0526_ ), .D(\us23\/_0527_ ), .X(\us23\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us23/_1313_ ( .A_N(\us23\/_0250_ ), .B(\us23\/_0521_ ), .Y(\us23\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1314_ ( .A(\us23\/_0128_ ), .B(\us23\/_0020_ ), .X(\us23\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1315_ ( .A(\us23\/_0530_ ), .Y(\us23\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1316_ ( .A(\us23\/_0099_ ), .B(\us23\/_0058_ ), .X(\us23\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1317_ ( .A(\us23\/_0533_ ), .Y(\us23\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us23/_1318_ ( .A_N(\us23\/_0529_ ), .B(\us23\/_0531_ ), .C(\us23\/_0534_ ), .D(\us23\/_0192_ ), .X(\us23\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1319_ ( .A(\us23\/_0434_ ), .B(\us23\/_0078_ ), .X(\us23\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us23/_1320_ ( .A1(\us23\/_0750_ ), .A2(\us23\/_0079_ ), .B1(\us23\/_0129_ ), .B2(\us23\/_0705_ ), .X(\us23\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1321_ ( .A1(\us23\/_0161_ ), .A2(\us23\/_0032_ ), .B1(\us23\/_0536_ ), .C1(\us23\/_0537_ ), .Y(\us23\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us23/_1322_ ( .A1(\us23\/_0746_ ), .A2(\us23\/_0162_ ), .B1(\us23\/_0079_ ), .B2(\us23\/_0043_ ), .X(\us23\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1323_ ( .A1(\us23\/_0093_ ), .A2(\us23\/_0247_ ), .B1(\us23\/_0240_ ), .C1(\us23\/_0539_ ), .Y(\us23\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1324_ ( .A(\us23\/_0434_ ), .B(\us23\/_0043_ ), .X(\us23\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us23/_1325_ ( .A1(\us23\/_0142_ ), .A2(\us23\/_0150_ ), .B1(\us23\/_0022_ ), .B2(\us23\/_0137_ ), .X(\us23\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1326_ ( .A1(\us23\/_0279_ ), .A2(\us23\/_0051_ ), .B1(\us23\/_0541_ ), .C1(\us23\/_0542_ ), .Y(\us23\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1327_ ( .A(\us23\/_0159_ ), .B(\us23\/_0035_ ), .X(\us23\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us23/_1328_ ( .A1(\us23\/_0271_ ), .A2(\us23\/_0434_ ), .B1(\us23\/_0027_ ), .X(\us23\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1329_ ( .A1(\us23\/_0091_ ), .A2(\us23\/_0128_ ), .B1(\us23\/_0545_ ), .C1(\us23\/_0546_ ), .Y(\us23\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1330_ ( .A(\us23\/_0538_ ), .B(\us23\/_0540_ ), .C(\us23\/_0544_ ), .D(\us23\/_0547_ ), .X(\us23\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1331_ ( .A(\us23\/_0099_ ), .B(\us23\/_0193_ ), .X(\us23\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us23/_1332_ ( .A(\us23\/_0549_ ), .B(\us23\/_0186_ ), .C(\us23\/_0187_ ), .Y(\us23\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1333_ ( .A(\us23\/_0062_ ), .B(\us23\/_0347_ ), .C(\us23\/_0749_ ), .D(\us23\/_0694_ ), .X(\us23\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1334_ ( .A1(\us23\/_0130_ ), .A2(\us23\/_0218_ ), .B1(\us23\/_0551_ ), .C1(\us23\/_0101_ ), .Y(\us23\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1335_ ( .A(\us23\/_0139_ ), .B(\us23\/_0640_ ), .Y(\us23\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1336_ ( .A1(\us23\/_0752_ ), .A2(\us23\/_0662_ ), .B1(\us23\/_0280_ ), .B2(\us23\/_0099_ ), .Y(\us23\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1337_ ( .A(\us23\/_0550_ ), .B(\us23\/_0552_ ), .C(\us23\/_0553_ ), .D(\us23\/_0555_ ), .X(\us23\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1338_ ( .A(\us23\/_0528_ ), .B(\us23\/_0535_ ), .C(\us23\/_0548_ ), .D(\us23\/_0556_ ), .X(\us23\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us23/_1339_ ( .A(\us23\/_0504_ ), .B(\us23\/_0519_ ), .C(\us23\/_0557_ ), .Y(\us23\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1340_ ( .A(\us23\/_0054_ ), .B(\us23\/_0507_ ), .X(\us23\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us23/_1341_ ( .A_N(\us23\/_0558_ ), .B(\us23\/_0408_ ), .C(\us23\/_0451_ ), .D(\us23\/_0452_ ), .X(\us23\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1342_ ( .A(\us23\/_0549_ ), .Y(\us23\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1343_ ( .A(\us23\/_0559_ ), .B(\us23\/_0403_ ), .C(\us23\/_0560_ ), .D(\us23\/_0371_ ), .X(\us23\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1344_ ( .A(\us23\/_0181_ ), .B(\us23\/_0178_ ), .X(\us23\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1345_ ( .A(\us23\/_0562_ ), .B(\us23\/_0552_ ), .C(\us23\/_0553_ ), .D(\us23\/_0555_ ), .X(\us23\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1346_ ( .A(\us23\/_0247_ ), .B(\us23\/_0020_ ), .Y(\us23\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1347_ ( .A(\us23\/_0051_ ), .B(\us23\/_0130_ ), .X(\us23\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1348_ ( .A(\us23\/_0566_ ), .Y(\us23\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1349_ ( .A(\us23\/_0159_ ), .B(\us23\/_0423_ ), .X(\us23\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1350_ ( .A1(\us23\/_0752_ ), .A2(\us23\/_0640_ ), .B1(\us23\/_0568_ ), .B2(\us23\/_0175_ ), .Y(\us23\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1351_ ( .A(\us23\/_0076_ ), .B(\us23\/_0565_ ), .C(\us23\/_0567_ ), .D(\us23\/_0569_ ), .X(\us23\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us23/_1352_ ( .A1(\us23\/_0035_ ), .A2(\us23\/_0142_ ), .B1(\us23\/_0161_ ), .X(\us23\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1353_ ( .A(\us23\/_0099_ ), .B(\us23\/_0662_ ), .Y(\us23\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us23/_1354_ ( .A(\us23\/_0420_ ), .B(\us23\/_0571_ ), .C_N(\us23\/_0572_ ), .Y(\us23\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1355_ ( .A(\us23\/_0051_ ), .B(\us23\/_0746_ ), .Y(\us23\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1356_ ( .A(\us23\/_0574_ ), .B(\us23\/_0319_ ), .C(\us23\/_0320_ ), .D(\us23\/_0411_ ), .X(\us23\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1357_ ( .A(\us23\/_0736_ ), .B(\us23\/_0035_ ), .Y(\us23\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1358_ ( .A(\us23\/_0736_ ), .B(\us23\/_0030_ ), .Y(\us23\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1359_ ( .A(\us23\/_0298_ ), .B(\us23\/_0208_ ), .C(\us23\/_0577_ ), .D(\us23\/_0578_ ), .X(\us23\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1360_ ( .A1(\us23\/_0020_ ), .A2(\us23\/_0137_ ), .B1(\us23\/_0261_ ), .B2(\us23\/_0128_ ), .Y(\us23\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1361_ ( .A(\us23\/_0573_ ), .B(\us23\/_0576_ ), .C(\us23\/_0579_ ), .D(\us23\/_0580_ ), .X(\us23\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1362_ ( .A(\us23\/_0561_ ), .B(\us23\/_0563_ ), .C(\us23\/_0570_ ), .D(\us23\/_0581_ ), .X(\us23\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1363_ ( .A(\us23\/_0128_ ), .B(\us23\/_0193_ ), .X(\us23\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1364_ ( .A(\us23\/_0082_ ), .B(\us23\/_0162_ ), .X(\us23\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us23/_1365_ ( .A(\us23\/_0583_ ), .B(\us23\/_0584_ ), .C_N(\us23\/_0437_ ), .Y(\us23\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us23/_1366_ ( .A(\us23\/_0150_ ), .B(\us23\/_0118_ ), .C(\us23\/_0380_ ), .Y(\us23\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us23/_1367_ ( .A_N(\us23\/_0182_ ), .B(\us23\/_0587_ ), .C(\us23\/_0323_ ), .X(\us23\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1368_ ( .A1(\us23\/_0575_ ), .A2(\us23\/_0153_ ), .B1(\us23\/_0727_ ), .B2(\us23\/_0058_ ), .Y(\us23\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1369_ ( .A1(\us23\/_0218_ ), .A2(\us23\/_0064_ ), .B1(\us23\/_0134_ ), .B2(\us23\/_0255_ ), .Y(\us23\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1370_ ( .A(\us23\/_0585_ ), .B(\us23\/_0588_ ), .C(\us23\/_0589_ ), .D(\us23\/_0590_ ), .X(\us23\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us23/_1371_ ( .A1(\us23\/_0091_ ), .A2(\us23\/_0139_ ), .B1(\us23\/_0250_ ), .Y(\us23\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1372_ ( .A1(\us23\/_0092_ ), .A2(\us23\/_0739_ ), .B1(\us23\/_0324_ ), .B2(\us23\/_0247_ ), .Y(\us23\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1373_ ( .A1(\us23\/_0144_ ), .A2(\us23\/_0153_ ), .B1(\us23\/_0683_ ), .B2(\us23\/_0056_ ), .Y(\us23\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1374_ ( .A1(\us23\/_0091_ ), .A2(\us23\/_0218_ ), .B1(\us23\/_0330_ ), .B2(\us23\/_0056_ ), .Y(\us23\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1375_ ( .A(\us23\/_0592_ ), .B(\us23\/_0593_ ), .C(\us23\/_0594_ ), .D(\us23\/_0595_ ), .X(\us23\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1376_ ( .A(\us23\/_0218_ ), .B(\us23\/_0144_ ), .Y(\us23\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1377_ ( .A(\us23\/_0312_ ), .B(\us23\/_0598_ ), .Y(\us23\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1378_ ( .A(\us23\/_0575_ ), .B(\us23\/_0147_ ), .Y(\us23\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1379_ ( .A1(\us23\/_0293_ ), .A2(\us23\/_0137_ ), .B1(\us23\/_0093_ ), .B2(\us23\/_0739_ ), .Y(\us23\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1380_ ( .A1(\us23\/_0734_ ), .A2(\us23\/_0531_ ), .B1(\us23\/_0600_ ), .C1(\us23\/_0601_ ), .Y(\us23\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1381_ ( .A1(\us23\/_0153_ ), .A2(\us23\/_0261_ ), .B1(\us23\/_0599_ ), .C1(\us23\/_0602_ ), .Y(\us23\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1382_ ( .A(\us23\/_0591_ ), .B(\us23\/_0596_ ), .C(\us23\/_0174_ ), .D(\us23\/_0603_ ), .X(\us23\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1383_ ( .A(\us23\/_0247_ ), .B(\us23\/_0144_ ), .Y(\us23\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1384_ ( .A(\us23\/_0113_ ), .B(\us23\/_0017_ ), .Y(\us23\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1385_ ( .A(\us23\/_0381_ ), .B(\us23\/_0605_ ), .C(\us23\/_0361_ ), .D(\us23\/_0606_ ), .X(\us23\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1386_ ( .A1(\us23\/_0016_ ), .A2(\us23\/_0727_ ), .B1(\us23\/_0733_ ), .Y(\us23\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1387_ ( .A1(\us23\/_0586_ ), .A2(\us23\/_0159_ ), .B1(\us23\/_0082_ ), .B2(\us23\/_0750_ ), .Y(\us23\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1388_ ( .A1(\us23\/_0142_ ), .A2(\us23\/_0162_ ), .B1(\us23\/_0079_ ), .B2(\us23\/_0054_ ), .Y(\us23\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1389_ ( .A(\us23\/_0610_ ), .B(\us23\/_0611_ ), .C(\us23\/_0105_ ), .D(\us23\/_0106_ ), .X(\us23\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1390_ ( .A1(\us23\/_0094_ ), .A2(\us23\/_0302_ ), .B1(\us23\/_0324_ ), .B2(\us23\/_0089_ ), .Y(\us23\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1391_ ( .A(\us23\/_0607_ ), .B(\us23\/_0609_ ), .C(\us23\/_0612_ ), .D(\us23\/_0613_ ), .X(\us23\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1392_ ( .A(\us23\/_0041_ ), .B(\us23\/_0170_ ), .X(\us23\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1393_ ( .A(\us23\/_0554_ ), .B(\us23\/_0027_ ), .X(\us23\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1394_ ( .A(\us23\/_0027_ ), .B(\us23\/_0261_ ), .Y(\us23\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us23/_1395_ ( .A_N(\us23\/_0616_ ), .B(\us23\/_0617_ ), .Y(\us23\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1396_ ( .A1(\us23\/_0147_ ), .A2(\us23\/_0302_ ), .B1(\us23\/_0342_ ), .C1(\us23\/_0618_ ), .Y(\us23\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1397_ ( .A(\us23\/_0614_ ), .B(\us23\/_0272_ ), .C(\us23\/_0615_ ), .D(\us23\/_0620_ ), .X(\us23\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us23/_1398_ ( .A(\us23\/_0582_ ), .B(\us23\/_0604_ ), .C(\us23\/_0621_ ), .Y(\us23\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1399_ ( .A1(\us23\/_0280_ ), .A2(\us23\/_0134_ ), .B1(\us23\/_0089_ ), .Y(\us23\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1400_ ( .A1(\us23\/_0144_ ), .A2(\us23\/_0608_ ), .A3(\us23\/_0330_ ), .B1(\us23\/_0089_ ), .Y(\us23\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1401_ ( .A1(\us23\/_0197_ ), .A2(\us23\/_0130_ ), .A3(\us23\/_0110_ ), .B1(\us23\/_0094_ ), .Y(\us23\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1402_ ( .A(\us23\/_0432_ ), .B(\us23\/_0622_ ), .C(\us23\/_0623_ ), .D(\us23\/_0624_ ), .X(\us23\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us23/_1403_ ( .A1(\us23\/_0554_ ), .A2(\us23\/_0017_ ), .A3(\us23\/_0022_ ), .B1(\us23\/_0161_ ), .X(\us23\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us23/_1404_ ( .A_N(\us23\/_0269_ ), .B(\us23\/_0170_ ), .X(\us23\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1405_ ( .A1(\us23\/_0109_ ), .A2(\us23\/_0064_ ), .A3(\us23\/_0733_ ), .B1(\us23\/_0355_ ), .Y(\us23\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us23/_1406_ ( .A_N(\us23\/_0626_ ), .B(\us23\/_0627_ ), .C(\us23\/_0353_ ), .D(\us23\/_0628_ ), .X(\us23\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1407_ ( .A1(\us23\/_0091_ ), .A2(\us23\/_0110_ ), .A3(\us23\/_0176_ ), .B1(\us23\/_0139_ ), .Y(\us23\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1408_ ( .A1(\us23\/_0020_ ), .A2(\us23\/_0261_ ), .B1(\us23\/_0147_ ), .Y(\us23\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1409_ ( .A(\us23\/_0631_ ), .B(\us23\/_0344_ ), .C(\us23\/_0421_ ), .D(\us23\/_0632_ ), .X(\us23\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us23/_1410_ ( .A1(\us23\/_0325_ ), .A2(\us23\/_0734_ ), .B1(\us23\/_0038_ ), .C1(\us23\/_0113_ ), .X(\us23\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1411_ ( .A1(\us23\/_0134_ ), .A2(\us23\/_0114_ ), .B1(\us23\/_0221_ ), .C1(\us23\/_0634_ ), .Y(\us23\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us23/_1412_ ( .A(\us23\/_0119_ ), .B_N(\us23\/_0111_ ), .Y(\us23\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1413_ ( .A1(\us23\/_0032_ ), .A2(\us23\/_0113_ ), .B1(\us23\/_0636_ ), .C1(\us23\/_0400_ ), .Y(\us23\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1414_ ( .A1(\us23\/_0731_ ), .A2(\us23\/_0293_ ), .A3(\us23\/_0251_ ), .B1(\us23\/_0099_ ), .Y(\us23\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1415_ ( .A(\us23\/_0189_ ), .B(\us23\/_0635_ ), .C(\us23\/_0637_ ), .D(\us23\/_0638_ ), .X(\us23\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1416_ ( .A(\us23\/_0625_ ), .B(\us23\/_0630_ ), .C(\us23\/_0633_ ), .D(\us23\/_0639_ ), .X(\us23\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1417_ ( .A(\us23\/_0746_ ), .B(\us23\/_0738_ ), .X(\us23\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1418_ ( .A(\us23\/_0736_ ), .B(\us23\/_0731_ ), .X(\us23\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us23/_1419_ ( .A_N(\us23\/_0643_ ), .B(\us23\/_0577_ ), .Y(\us23\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1420_ ( .A1(\us23\/_0280_ ), .A2(\us23\/_0739_ ), .B1(\us23\/_0642_ ), .C1(\us23\/_0644_ ), .Y(\us23\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1421_ ( .A1(\us23\/_0050_ ), .A2(\us23\/_0543_ ), .B1(\us23\/_0194_ ), .C1(\us23\/_0738_ ), .Y(\us23\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1422_ ( .A(\us23\/_0646_ ), .B(\us23\/_0232_ ), .C(\us23\/_0417_ ), .D(\us23\/_0578_ ), .X(\us23\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1423_ ( .A1(\us23\/_0064_ ), .A2(\us23\/_0733_ ), .B1(\us23\/_0727_ ), .Y(\us23\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1424_ ( .A1(\us23\/_0193_ ), .A2(\us23\/_0276_ ), .B1(\us23\/_0727_ ), .Y(\us23\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1425_ ( .A(\us23\/_0645_ ), .B(\us23\/_0647_ ), .C(\us23\/_0648_ ), .D(\us23\/_0649_ ), .X(\us23\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1426_ ( .A1(\us23\/_0325_ ), .A2(\us23\/_0734_ ), .B1(\us23\/_0038_ ), .C1(\us23\/_0247_ ), .Y(\us23\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1427_ ( .A1(\us23\/_0543_ ), .A2(\us23\/_0205_ ), .B1(\us23\/_0423_ ), .C1(\us23\/_0247_ ), .Y(\us23\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1428_ ( .A(\us23\/_0652_ ), .B(\us23\/_0653_ ), .X(\us23\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1429_ ( .A1(\us23\/_0733_ ), .A2(\us23\/_0748_ ), .A3(\us23\/_0324_ ), .B1(\us23\/_0016_ ), .Y(\us23\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1430_ ( .A1(\us23\/_0640_ ), .A2(\us23\/_0193_ ), .A3(\us23\/_0091_ ), .B1(\us23\/_0016_ ), .Y(\us23\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1431_ ( .A1(\us23\/_0102_ ), .A2(\us23\/_0301_ ), .B1(\sa23\[3\] ), .C1(\us23\/_0247_ ), .Y(\us23\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1432_ ( .A(\us23\/_0654_ ), .B(\us23\/_0655_ ), .C(\us23\/_0656_ ), .D(\us23\/_0657_ ), .X(\us23\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1433_ ( .A1(\us23\/_0118_ ), .A2(\us23\/_0050_ ), .B1(\us23\/_0038_ ), .C1(\us23\/_0478_ ), .Y(\us23\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us23/_1434_ ( .A_N(\us23\/_0250_ ), .B(\us23\/_0465_ ), .C(\us23\/_0659_ ), .X(\us23\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1435_ ( .A1(\us23\/_0683_ ), .A2(\us23\/_0324_ ), .B1(\us23\/_0255_ ), .Y(\us23\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1436_ ( .A1(\us23\/_0032_ ), .A2(\us23\/_0193_ ), .A3(\us23\/_0047_ ), .B1(\us23\/_0255_ ), .Y(\us23\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1437_ ( .A1(\us23\/_0144_ ), .A2(\us23\/_0586_ ), .A3(\us23\/_0047_ ), .B1(\us23\/_0218_ ), .Y(\us23\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1438_ ( .A(\us23\/_0660_ ), .B(\us23\/_0661_ ), .C(\us23\/_0663_ ), .D(\us23\/_0664_ ), .X(\us23\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1439_ ( .A1(\us23\/_0091_ ), .A2(\us23\/_0276_ ), .B1(\us23\/_0060_ ), .Y(\us23\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1440_ ( .A1(\us23\/_0144_ ), .A2(\us23\/_0608_ ), .B1(\us23\/_0056_ ), .Y(\us23\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1441_ ( .A1(\us23\/_0423_ ), .A2(\us23\/_0038_ ), .B1(\us23\/_0102_ ), .C1(\us23\/_0060_ ), .Y(\us23\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1442_ ( .A1(\sa23\[1\] ), .A2(\us23\/_0734_ ), .B1(\us23\/_0109_ ), .C1(\us23\/_0056_ ), .Y(\us23\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1443_ ( .A(\us23\/_0666_ ), .B(\us23\/_0667_ ), .C(\us23\/_0668_ ), .D(\us23\/_0669_ ), .X(\us23\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1444_ ( .A(\us23\/_0650_ ), .B(\us23\/_0658_ ), .C(\us23\/_0665_ ), .D(\us23\/_0670_ ), .X(\us23\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us23/_1445_ ( .A(\us23\/_0641_ ), .B(\us23\/_0174_ ), .C(\us23\/_0671_ ), .Y(\us23\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us23/_1446_ ( .A(\us23\/_0049_ ), .B(\us23\/_0618_ ), .C_N(\us23\/_0052_ ), .Y(\us23\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us23/_1447_ ( .A(\us23\/_0239_ ), .Y(\us23\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1448_ ( .A(\us23\/_0705_ ), .B(\us23\/_0032_ ), .Y(\us23\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1449_ ( .A1(\us23\/_0054_ ), .A2(\us23\/_0731_ ), .B1(\us23\/_0035_ ), .B2(\us23\/_0705_ ), .Y(\us23\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1450_ ( .A1(\us23\/_0304_ ), .A2(\us23\/_0731_ ), .B1(\us23\/_0047_ ), .B2(\us23\/_0750_ ), .Y(\us23\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1451_ ( .A(\us23\/_0674_ ), .B(\us23\/_0675_ ), .C(\us23\/_0676_ ), .D(\us23\/_0677_ ), .X(\us23\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us23/_1452_ ( .A_N(\us23\/_0584_ ), .B(\us23\/_0283_ ), .X(\us23\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1453_ ( .A(\us23\/_0673_ ), .B(\us23\/_0678_ ), .C(\us23\/_0679_ ), .D(\us23\/_0508_ ), .X(\us23\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1454_ ( .A1(\us23\/_0016_ ), .A2(\us23\/_0733_ ), .B1(\us23\/_0355_ ), .B2(\us23\/_0092_ ), .Y(\us23\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1455_ ( .A(\us23\/_0681_ ), .B(\us23\/_0034_ ), .X(\us23\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us23/_1456_ ( .A1(\us23\/_0330_ ), .A2(\us23\/_0139_ ), .B1(\us23\/_0324_ ), .B2(\us23\/_0089_ ), .X(\us23\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1457_ ( .A1(\us23\/_0146_ ), .A2(\us23\/_0147_ ), .B1(\us23\/_0133_ ), .C1(\us23\/_0684_ ), .Y(\us23\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1458_ ( .A(\us23\/_0113_ ), .B(\us23\/_0251_ ), .Y(\us23\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us23/_1459_ ( .A_N(\us23\/_0463_ ), .B(\us23\/_0686_ ), .C(\us23\/_0383_ ), .D(\us23\/_0464_ ), .X(\us23\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1460_ ( .A1(\us23\/_0051_ ), .A2(\us23\/_0293_ ), .B1(\us23\/_0280_ ), .B2(\us23\/_0705_ ), .Y(\us23\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1461_ ( .A1(\us23\/_0017_ ), .A2(\us23\/_0072_ ), .B1(\us23\/_0134_ ), .B2(\us23\/_0078_ ), .Y(\us23\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1462_ ( .A(\us23\/_0687_ ), .B(\us23\/_0236_ ), .C(\us23\/_0688_ ), .D(\us23\/_0689_ ), .X(\us23\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1463_ ( .A(\us23\/_0680_ ), .B(\us23\/_0682_ ), .C(\us23\/_0685_ ), .D(\us23\/_0690_ ), .X(\us23\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us23/_1464_ ( .A1(\us23\/_0532_ ), .A2(\us23\/_0380_ ), .B1(\us23\/_0102_ ), .C1(\us23\/_0355_ ), .X(\us23\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us23/_1465_ ( .A(\us23\/_0692_ ), .B(\us23\/_0338_ ), .C(\us23\/_0644_ ), .Y(\us23\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1466_ ( .A(\us23\/_0016_ ), .B(\us23\/_0020_ ), .Y(\us23\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1467_ ( .A1(\us23\/_0032_ ), .A2(\us23\/_0137_ ), .B1(\us23\/_0279_ ), .B2(\us23\/_0094_ ), .Y(\us23\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1468_ ( .A1(\us23\/_0575_ ), .A2(\us23\/_0153_ ), .B1(\us23\/_0161_ ), .B2(\us23\/_0293_ ), .Y(\us23\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1469_ ( .A(\us23\/_0259_ ), .B(\us23\/_0695_ ), .C(\us23\/_0696_ ), .D(\us23\/_0697_ ), .X(\us23\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us23/_1470_ ( .A1(\us23\/_0255_ ), .A2(\us23\/_0640_ ), .B1(\us23\/_0016_ ), .B2(\us23\/_0193_ ), .X(\us23\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1471_ ( .A1(\us23\/_0060_ ), .A2(\us23\/_0176_ ), .B1(\us23\/_0699_ ), .C1(\us23\/_0177_ ), .Y(\us23\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1472_ ( .A1(\us23\/_0091_ ), .A2(\us23\/_0218_ ), .B1(\us23\/_0092_ ), .B2(\us23\/_0705_ ), .Y(\us23\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us23/_1473_ ( .A1(\us23\/_0705_ ), .A2(\us23\/_0683_ ), .B1(\us23\/_0093_ ), .B2(\us23\/_0114_ ), .Y(\us23\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us23/_1474_ ( .A1(\us23\/_0683_ ), .A2(\us23\/_0280_ ), .B1(\us23\/_0094_ ), .Y(\us23\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us23/_1475_ ( .A1(\us23\/_0543_ ), .A2(\us23\/_0205_ ), .B1(\us23\/_0038_ ), .C1(\us23\/_0056_ ), .Y(\us23\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1476_ ( .A(\us23\/_0701_ ), .B(\us23\/_0702_ ), .C(\us23\/_0703_ ), .D(\us23\/_0704_ ), .X(\us23\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1477_ ( .A(\us23\/_0693_ ), .B(\us23\/_0698_ ), .C(\us23\/_0700_ ), .D(\us23\/_0706_ ), .X(\us23\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us23/_1478_ ( .A1(\us23\/_0113_ ), .A2(\us23\/_0640_ ), .B1(\us23\/_0099_ ), .B2(\us23\/_0058_ ), .X(\us23\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us23/_1479_ ( .A(\us23\/_0407_ ), .B(\us23\/_0708_ ), .C(\us23\/_0529_ ), .Y(\us23\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1480_ ( .A(\us23\/_0568_ ), .B(\us23\/_0175_ ), .Y(\us23\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us23/_1481_ ( .A1(\us23\/_0247_ ), .A2(\us23\/_0114_ ), .A3(\us23\/_0051_ ), .B1(\us23\/_0130_ ), .Y(\us23\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1482_ ( .A(\us23\/_0709_ ), .B(\us23\/_0550_ ), .C(\us23\/_0710_ ), .D(\us23\/_0711_ ), .X(\us23\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us23/_1483_ ( .A1(\us23\/_0114_ ), .A2(\us23\/_0064_ ), .B1(\us23\/_0261_ ), .B2(\us23\/_0089_ ), .X(\us23\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1484_ ( .A1(\us23\/_0355_ ), .A2(\us23\/_0261_ ), .B1(\us23\/_0198_ ), .C1(\us23\/_0713_ ), .Y(\us23\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1485_ ( .A(\us23\/_0586_ ), .B(\us23\/_0478_ ), .Y(\us23\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us23/_1486_ ( .A_N(\us23\/_0541_ ), .B(\us23\/_0267_ ), .C(\us23\/_0715_ ), .D(\us23\/_0320_ ), .X(\us23\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1487_ ( .A(\us23\/_0586_ ), .B(\us23\/_0070_ ), .Y(\us23\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us23/_1488_ ( .A_N(\us23\/_0211_ ), .B(\us23\/_0155_ ), .C(\us23\/_0202_ ), .D(\us23\/_0718_ ), .X(\us23\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us23/_1489_ ( .A(\us23\/_0150_ ), .B(\us23\/_0205_ ), .C(\us23\/_0380_ ), .Y(\us23\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us23/_1490_ ( .A(\us23\/_0411_ ), .B(\us23\/_0720_ ), .X(\us23\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us23/_1491_ ( .A1(\us23\/_0017_ ), .A2(\us23\/_0022_ ), .B1(\us23\/_0078_ ), .X(\us23\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us23/_1492_ ( .A1(\us23\/_0134_ ), .A2(\us23\/_0738_ ), .B1(\us23\/_0101_ ), .C1(\us23\/_0722_ ), .Y(\us23\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1493_ ( .A(\us23\/_0717_ ), .B(\us23\/_0719_ ), .C(\us23\/_0721_ ), .D(\us23\/_0723_ ), .X(\us23\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us23/_1494_ ( .A(\us23\/_0739_ ), .B(\us23\/_0193_ ), .Y(\us23\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1495_ ( .A(\us23\/_0344_ ), .B(\us23\/_0184_ ), .C(\us23\/_0449_ ), .D(\us23\/_0725_ ), .X(\us23\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us23/_1496_ ( .A(\us23\/_0712_ ), .B(\us23\/_0714_ ), .C(\us23\/_0724_ ), .D(\us23\/_0726_ ), .X(\us23\/_0728_ ) );
sky130_fd_sc_hd__nand3_2 \us23/_1497_ ( .A(\us23\/_0691_ ), .B(\us23\/_0707_ ), .C(\us23\/_0728_ ), .Y(\us23\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \us30/_0753_ ( .A(\sa30\[2\] ), .B_N(\sa30\[3\] ), .Y(\us30\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \us30/_0755_ ( .A(\sa30\[1\] ), .B(\sa30\[0\] ), .X(\us30\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us30/_0756_ ( .A(\us30\/_0096_ ), .B(\us30\/_0118_ ), .X(\us30\/_0129_ ) );
sky130_fd_sc_hd__and2_1 \us30/_0757_ ( .A(\sa30\[7\] ), .B(\sa30\[6\] ), .X(\us30\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_0758_ ( .A(\sa30\[4\] ), .B(\sa30\[5\] ), .Y(\us30\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0759_ ( .A(\us30\/_0140_ ), .B(\us30\/_0151_ ), .X(\us30\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0761_ ( .A(\us30\/_0129_ ), .B(\us30\/_0162_ ), .X(\us30\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0762_ ( .A(\us30\/_0096_ ), .X(\us30\/_0194_ ) );
sky130_fd_sc_hd__nor2b_2 \us30/_0763_ ( .A(\sa30\[1\] ), .B_N(\sa30\[0\] ), .Y(\us30\/_0205_ ) );
sky130_fd_sc_hd__and3_1 \us30/_0765_ ( .A(\us30\/_0162_ ), .B(\us30\/_0194_ ), .C(\us30\/_0205_ ), .X(\us30\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us30/_0766_ ( .A(\us30\/_0183_ ), .SLEEP(\us30\/_0227_ ), .X(\us30\/_0238_ ) );
sky130_fd_sc_hd__nor2b_2 \us30/_0767_ ( .A(\sa30\[0\] ), .B_N(\sa30\[1\] ), .Y(\us30\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_0768_ ( .A(\sa30\[2\] ), .B(\sa30\[3\] ), .Y(\us30\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0769_ ( .A(\us30\/_0249_ ), .B(\us30\/_0260_ ), .X(\us30\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0771_ ( .A(\us30\/_0271_ ), .X(\us30\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0772_ ( .A(\us30\/_0162_ ), .X(\us30\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_0773_ ( .A(\us30\/_0293_ ), .B(\us30\/_0304_ ), .Y(\us30\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us30/_0774_ ( .A(\sa30\[1\] ), .Y(\us30\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us30/_0776_ ( .A(\sa30\[0\] ), .Y(\us30\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0777_ ( .A(\sa30\[2\] ), .B(\sa30\[3\] ), .X(\us30\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0779_ ( .A(\us30\/_0358_ ), .X(\us30\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_0780_ ( .A1(\us30\/_0325_ ), .A2(\us30\/_0347_ ), .B1(\us30\/_0380_ ), .C1(\us30\/_0304_ ), .Y(\us30\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us30/_0781_ ( .A_N(\us30\/_0238_ ), .B(\us30\/_0314_ ), .C(\us30\/_0391_ ), .X(\us30\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us30/_0782_ ( .A(\sa30\[3\] ), .B_N(\sa30\[2\] ), .Y(\us30\/_0412_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0784_ ( .A(\us30\/_0412_ ), .B(\us30\/_0205_ ), .X(\us30\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \us30/_0787_ ( .A(\sa30\[5\] ), .B_N(\sa30\[4\] ), .Y(\us30\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0788_ ( .A(\us30\/_0467_ ), .B(\us30\/_0140_ ), .X(\us30\/_0478_ ) );
sky130_fd_sc_hd__buf_2 \us30/_0790_ ( .A(\us30\/_0478_ ), .X(\us30\/_0499_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_0791_ ( .A(\us30\/_0134_ ), .B(\us30\/_0499_ ), .Y(\us30\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_0792_ ( .A(\us30\/_0478_ ), .B(\us30\/_0271_ ), .Y(\us30\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0793_ ( .A(\us30\/_0194_ ), .X(\us30\/_0532_ ) );
sky130_fd_sc_hd__and2_1 \us30/_0795_ ( .A(\us30\/_0249_ ), .B(\us30\/_0358_ ), .X(\us30\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0797_ ( .A(\us30\/_0554_ ), .X(\us30\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us30/_0798_ ( .A(\us30\/_0205_ ), .B(\us30\/_0358_ ), .X(\us30\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0800_ ( .A(\us30\/_0586_ ), .X(\us30\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_0801_ ( .A1(\us30\/_0532_ ), .A2(\us30\/_0575_ ), .A3(\us30\/_0608_ ), .B1(\us30\/_0499_ ), .Y(\us30\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us30/_0802_ ( .A(\us30\/_0401_ ), .B(\us30\/_0510_ ), .C(\us30\/_0521_ ), .D(\us30\/_0619_ ), .X(\us30\/_0629_ ) );
sky130_fd_sc_hd__and2_1 \us30/_0803_ ( .A(\us30\/_0358_ ), .B(\sa30\[1\] ), .X(\us30\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0805_ ( .A(\us30\/_0205_ ), .B(\us30\/_0260_ ), .X(\us30\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0807_ ( .A(\us30\/_0662_ ), .X(\us30\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us30/_0808_ ( .A(\sa30\[6\] ), .B_N(\sa30\[7\] ), .Y(\us30\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \us30/_0809_ ( .A(\us30\/_0467_ ), .B(\us30\/_0694_ ), .X(\us30\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0811_ ( .A(\us30\/_0705_ ), .X(\us30\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_0812_ ( .A1(\us30\/_0640_ ), .A2(\us30\/_0293_ ), .A3(\us30\/_0683_ ), .B1(\us30\/_0727_ ), .Y(\us30\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_0813_ ( .A(\sa30\[1\] ), .B(\sa30\[0\] ), .Y(\us30\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0814_ ( .A(\us30\/_0730_ ), .B(\us30\/_0260_ ), .X(\us30\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0816_ ( .A(\us30\/_0731_ ), .X(\us30\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0817_ ( .A(\sa30\[0\] ), .X(\us30\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us30/_0818_ ( .A1(\us30\/_0325_ ), .A2(\us30\/_0734_ ), .B1(\us30\/_0412_ ), .X(\us30\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0819_ ( .A(\us30\/_0694_ ), .B(\us30\/_0151_ ), .X(\us30\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0821_ ( .A(\us30\/_0736_ ), .X(\us30\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0822_ ( .A(\us30\/_0738_ ), .X(\us30\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_0823_ ( .A1(\us30\/_0733_ ), .A2(\us30\/_0735_ ), .A3(\us30\/_0293_ ), .B1(\us30\/_0739_ ), .Y(\us30\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us30/_0824_ ( .A(\us30\/_0730_ ), .B_N(\us30\/_0358_ ), .Y(\us30\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_0825_ ( .A(\us30\/_0741_ ), .B(\us30\/_0739_ ), .Y(\us30\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_0827_ ( .A1(\us30\/_0118_ ), .A2(\us30\/_0205_ ), .B1(\us30\/_0532_ ), .C1(\us30\/_0739_ ), .Y(\us30\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us30/_0828_ ( .A(\us30\/_0729_ ), .B(\us30\/_0740_ ), .C(\us30\/_0742_ ), .D(\us30\/_0744_ ), .X(\us30\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0829_ ( .A(\us30\/_0412_ ), .B(\us30\/_0730_ ), .X(\us30\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0831_ ( .A(\us30\/_0746_ ), .X(\us30\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us30/_0832_ ( .A(\sa30\[4\] ), .B_N(\sa30\[5\] ), .Y(\us30\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0833_ ( .A(\us30\/_0749_ ), .B(\us30\/_0694_ ), .X(\us30\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0835_ ( .A(\us30\/_0750_ ), .X(\us30\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0836_ ( .A(\us30\/_0752_ ), .X(\us30\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0837_ ( .A(\us30\/_0118_ ), .B(\us30\/_0358_ ), .X(\us30\/_0017_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0839_ ( .A(\us30\/_0752_ ), .B(\us30\/_0017_ ), .X(\us30\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0840_ ( .A(\us30\/_0358_ ), .B(\us30\/_0325_ ), .X(\us30\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0842_ ( .A(\us30\/_0096_ ), .B(\us30\/_0205_ ), .X(\us30\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \us30/_0844_ ( .A1(\us30\/_0020_ ), .A2(\us30\/_0022_ ), .B1(\us30\/_0752_ ), .X(\us30\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_0845_ ( .A1(\us30\/_0748_ ), .A2(\us30\/_0016_ ), .B1(\us30\/_0019_ ), .C1(\us30\/_0024_ ), .Y(\us30\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \us30/_0846_ ( .A(\sa30\[4\] ), .B(\sa30\[5\] ), .X(\us30\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0847_ ( .A(\us30\/_0694_ ), .B(\us30\/_0026_ ), .X(\us30\/_0027_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0850_ ( .A(\us30\/_0358_ ), .B(\us30\/_0730_ ), .X(\us30\/_0030_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0852_ ( .A(\us30\/_0030_ ), .X(\us30\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_0853_ ( .A(\us30\/_0247_ ), .B(\us30\/_0032_ ), .Y(\us30\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_0854_ ( .A(\us30\/_0247_ ), .B(\us30\/_0735_ ), .Y(\us30\/_0034_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0855_ ( .A(\us30\/_0118_ ), .B(\us30\/_0260_ ), .X(\us30\/_0035_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0857_ ( .A(\us30\/_0027_ ), .B(\us30\/_0035_ ), .X(\us30\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0858_ ( .A(\us30\/_0260_ ), .X(\us30\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_0859_ ( .A(\us30\/_0038_ ), .B(\us30\/_0347_ ), .Y(\us30\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us30/_0860_ ( .A_N(\us30\/_0039_ ), .B(\us30\/_0027_ ), .X(\us30\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_0861_ ( .A(\us30\/_0037_ ), .B(\us30\/_0040_ ), .Y(\us30\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us30/_0862_ ( .A(\us30\/_0025_ ), .B(\us30\/_0033_ ), .C(\us30\/_0034_ ), .D(\us30\/_0041_ ), .X(\us30\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0863_ ( .A(\us30\/_0749_ ), .B(\us30\/_0140_ ), .X(\us30\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us30/_0865_ ( .A(\sa30\[0\] ), .B(\sa30\[2\] ), .C(\sa30\[3\] ), .X(\us30\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0866_ ( .A(\us30\/_0043_ ), .B(\us30\/_0045_ ), .X(\us30\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0867_ ( .A(\us30\/_0096_ ), .B(\us30\/_0249_ ), .X(\us30\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0869_ ( .A(\us30\/_0047_ ), .B(\us30\/_0043_ ), .X(\us30\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0870_ ( .A(\us30\/_0730_ ), .X(\us30\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0871_ ( .A(\us30\/_0043_ ), .X(\us30\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_0872_ ( .A1(\us30\/_0118_ ), .A2(\us30\/_0050_ ), .B1(\us30\/_0194_ ), .C1(\us30\/_0051_ ), .Y(\us30\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us30/_0873_ ( .A(\us30\/_0046_ ), .B(\us30\/_0049_ ), .C_N(\us30\/_0052_ ), .Y(\us30\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0874_ ( .A(\us30\/_0026_ ), .B(\us30\/_0140_ ), .X(\us30\/_0054_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_0877_ ( .A1(\us30\/_0532_ ), .A2(\us30\/_0575_ ), .B1(\us30\/_0292_ ), .Y(\us30\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0878_ ( .A(\us30\/_0412_ ), .B(\us30\/_0325_ ), .X(\us30\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0880_ ( .A(\us30\/_0051_ ), .X(\us30\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_0881_ ( .A1(\us30\/_0731_ ), .A2(\us30\/_0035_ ), .A3(\us30\/_0058_ ), .B1(\us30\/_0060_ ), .Y(\us30\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0882_ ( .A(\us30\/_0260_ ), .B(\sa30\[1\] ), .X(\us30\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0884_ ( .A(\us30\/_0062_ ), .X(\us30\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_0885_ ( .A1(\us30\/_0064_ ), .A2(\us30\/_0748_ ), .A3(\us30\/_0683_ ), .B1(\us30\/_0292_ ), .Y(\us30\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us30/_0886_ ( .A(\us30\/_0053_ ), .B(\us30\/_0057_ ), .C(\us30\/_0061_ ), .D(\us30\/_0065_ ), .X(\us30\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us30/_0887_ ( .A(\us30\/_0629_ ), .B(\us30\/_0745_ ), .C(\us30\/_0042_ ), .D(\us30\/_0066_ ), .X(\us30\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us30/_0889_ ( .A(\sa30\[7\] ), .B_N(\sa30\[6\] ), .Y(\us30\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0890_ ( .A(\us30\/_0069_ ), .B(\us30\/_0151_ ), .X(\us30\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0892_ ( .A(\us30\/_0070_ ), .X(\us30\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_0893_ ( .A1(\us30\/_0129_ ), .A2(\us30\/_0586_ ), .B1(\us30\/_0072_ ), .Y(\us30\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_0894_ ( .A1(\us30\/_0380_ ), .A2(\us30\/_0347_ ), .B1(\us30\/_0194_ ), .B2(\us30\/_0205_ ), .Y(\us30\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us30/_0895_ ( .A(\us30\/_0074_ ), .B_N(\us30\/_0070_ ), .Y(\us30\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us30/_0896_ ( .A(\us30\/_0073_ ), .SLEEP(\us30\/_0075_ ), .X(\us30\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us30/_0897_ ( .A(\us30\/_0467_ ), .B(\us30\/_0069_ ), .X(\us30\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0898_ ( .A(\us30\/_0077_ ), .X(\us30\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0899_ ( .A(\us30\/_0412_ ), .B(\us30\/_0118_ ), .X(\us30\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0901_ ( .A(\us30\/_0078_ ), .B(\us30\/_0079_ ), .X(\us30\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0902_ ( .A(\us30\/_0412_ ), .B(\us30\/_0249_ ), .X(\us30\/_0082_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0905_ ( .A(\us30\/_0280_ ), .B(\us30\/_0078_ ), .X(\us30\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us30/_0906_ ( .A1(\sa30\[0\] ), .A2(\us30\/_0325_ ), .B1(\us30\/_0260_ ), .Y(\us30\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us30/_0907_ ( .A_N(\us30\/_0086_ ), .B(\us30\/_0078_ ), .X(\us30\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us30/_0908_ ( .A(\us30\/_0081_ ), .B(\us30\/_0085_ ), .C(\us30\/_0087_ ), .Y(\us30\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0909_ ( .A(\us30\/_0072_ ), .X(\us30\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_0910_ ( .A1(\us30\/_0733_ ), .A2(\us30\/_0748_ ), .A3(\us30\/_0683_ ), .B1(\us30\/_0089_ ), .Y(\us30\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0911_ ( .A(\us30\/_0129_ ), .X(\us30\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0912_ ( .A(\us30\/_0017_ ), .X(\us30\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0913_ ( .A(\us30\/_0022_ ), .X(\us30\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0914_ ( .A(\us30\/_0078_ ), .X(\us30\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_0915_ ( .A1(\us30\/_0091_ ), .A2(\us30\/_0092_ ), .A3(\us30\/_0093_ ), .B1(\us30\/_0094_ ), .Y(\us30\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us30/_0916_ ( .A(\us30\/_0076_ ), .B(\us30\/_0088_ ), .C(\us30\/_0090_ ), .D(\us30\/_0095_ ), .X(\us30\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us30/_0917_ ( .A(\us30\/_0069_ ), .B(\us30\/_0026_ ), .X(\us30\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \us30/_0918_ ( .A(\us30\/_0098_ ), .X(\us30\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0919_ ( .A(\us30\/_0434_ ), .B(\us30\/_0099_ ), .X(\us30\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0920_ ( .A(\us30\/_0079_ ), .B(\us30\/_0098_ ), .X(\us30\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0921_ ( .A(\us30\/_0325_ ), .X(\us30\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_0922_ ( .A1(\us30\/_0102_ ), .A2(\us30\/_0734_ ), .B1(\us30\/_0038_ ), .C1(\us30\/_0099_ ), .Y(\us30\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us30/_0923_ ( .A(\us30\/_0100_ ), .B(\us30\/_0101_ ), .C_N(\us30\/_0103_ ), .Y(\us30\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_0924_ ( .A1(\us30\/_0554_ ), .A2(\us30\/_0586_ ), .B1(\us30\/_0099_ ), .Y(\us30\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_0925_ ( .A(\us30\/_0129_ ), .B(\us30\/_0099_ ), .Y(\us30\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0926_ ( .A(\us30\/_0105_ ), .B(\us30\/_0106_ ), .X(\us30\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0927_ ( .A(\us30\/_0412_ ), .X(\us30\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us30/_0928_ ( .A(\us30\/_0260_ ), .B(\sa30\[0\] ), .X(\us30\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0929_ ( .A(\us30\/_0069_ ), .B(\us30\/_0749_ ), .X(\us30\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0931_ ( .A(\us30\/_0111_ ), .X(\us30\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0932_ ( .A(\us30\/_0113_ ), .X(\us30\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_0933_ ( .A1(\us30\/_0109_ ), .A2(\us30\/_0110_ ), .B1(\us30\/_0114_ ), .Y(\us30\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us30/_0934_ ( .A(\us30\/_0022_ ), .Y(\us30\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us30/_0935_ ( .A(\us30\/_0554_ ), .Y(\us30\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us30/_0936_ ( .A1(\us30\/_0050_ ), .A2(\us30\/_0118_ ), .B1(\us30\/_0194_ ), .Y(\us30\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us30/_0937_ ( .A(\us30\/_0113_ ), .Y(\us30\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us30/_0938_ ( .A1(\us30\/_0116_ ), .A2(\us30\/_0117_ ), .A3(\us30\/_0119_ ), .B1(\us30\/_0120_ ), .X(\us30\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us30/_0939_ ( .A(\us30\/_0104_ ), .B(\us30\/_0108_ ), .C(\us30\/_0115_ ), .D(\us30\/_0121_ ), .X(\us30\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_0940_ ( .A(\sa30\[7\] ), .B(\sa30\[6\] ), .Y(\us30\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0941_ ( .A(\us30\/_0749_ ), .B(\us30\/_0123_ ), .X(\us30\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0943_ ( .A(\us30\/_0082_ ), .B(\us30\/_0124_ ), .X(\us30\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_0944_ ( .A(\us30\/_0271_ ), .B(\us30\/_0124_ ), .Y(\us30\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0945_ ( .A(\us30\/_0124_ ), .X(\us30\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0946_ ( .A(\us30\/_0260_ ), .B(\us30\/_0325_ ), .X(\us30\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_0948_ ( .A(\us30\/_0128_ ), .B(\us30\/_0130_ ), .Y(\us30\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_0949_ ( .A(\us30\/_0127_ ), .B(\us30\/_0132_ ), .Y(\us30\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us30/_0950_ ( .A(\us30\/_0434_ ), .X(\us30\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_0951_ ( .A(\us30\/_0134_ ), .B(\us30\/_0128_ ), .Y(\us30\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us30/_0952_ ( .A(\us30\/_0126_ ), .B(\us30\/_0133_ ), .C_N(\us30\/_0135_ ), .Y(\us30\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us30/_0953_ ( .A(\us30\/_0026_ ), .B(\us30\/_0123_ ), .X(\us30\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0955_ ( .A(\us30\/_0137_ ), .X(\us30\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_0956_ ( .A1(\us30\/_0110_ ), .A2(\us30\/_0293_ ), .A3(\us30\/_0280_ ), .B1(\us30\/_0139_ ), .Y(\us30\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0957_ ( .A(\us30\/_0096_ ), .B(\us30\/_0730_ ), .X(\us30\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0959_ ( .A(\us30\/_0142_ ), .X(\us30\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_0960_ ( .A1(\us30\/_0020_ ), .A2(\us30\/_0144_ ), .A3(\us30\/_0017_ ), .B1(\us30\/_0139_ ), .Y(\us30\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \us30/_0961_ ( .A(\sa30\[2\] ), .B(\us30\/_0050_ ), .C_N(\sa30\[3\] ), .Y(\us30\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0962_ ( .A(\us30\/_0128_ ), .X(\us30\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_0963_ ( .A1(\us30\/_0146_ ), .A2(\us30\/_0032_ ), .A3(\us30\/_0640_ ), .B1(\us30\/_0147_ ), .Y(\us30\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us30/_0964_ ( .A(\us30\/_0136_ ), .B(\us30\/_0141_ ), .C(\us30\/_0145_ ), .D(\us30\/_0148_ ), .X(\us30\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0965_ ( .A(\us30\/_0123_ ), .B(\us30\/_0151_ ), .X(\us30\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0967_ ( .A(\us30\/_0150_ ), .X(\us30\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \us30/_0968_ ( .A(\us30\/_0150_ ), .B(\us30\/_0062_ ), .X(\us30\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_0969_ ( .A(\us30\/_0079_ ), .B(\us30\/_0150_ ), .Y(\us30\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us30/_0970_ ( .A(\us30\/_0150_ ), .B(\us30\/_0412_ ), .C(\us30\/_0249_ ), .Y(\us30\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_0971_ ( .A(\us30\/_0155_ ), .B(\us30\/_0156_ ), .Y(\us30\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_0972_ ( .A1(\us30\/_0153_ ), .A2(\us30\/_0134_ ), .B1(\us30\/_0154_ ), .C1(\us30\/_0157_ ), .Y(\us30\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0973_ ( .A(\us30\/_0467_ ), .B(\us30\/_0123_ ), .X(\us30\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_0975_ ( .A(\us30\/_0159_ ), .X(\us30\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us30/_0976_ ( .A_N(\us30\/_0119_ ), .B(\us30\/_0161_ ), .X(\us30\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us30/_0977_ ( .A(\us30\/_0163_ ), .Y(\us30\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_0978_ ( .A1(\us30\/_0146_ ), .A2(\us30\/_0575_ ), .A3(\us30\/_0608_ ), .B1(\us30\/_0153_ ), .Y(\us30\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_0979_ ( .A1(\us30\/_0062_ ), .A2(\us30\/_0280_ ), .A3(\us30\/_0134_ ), .B1(\us30\/_0161_ ), .Y(\us30\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us30/_0980_ ( .A(\us30\/_0158_ ), .B(\us30\/_0164_ ), .C(\us30\/_0165_ ), .D(\us30\/_0166_ ), .X(\us30\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us30/_0981_ ( .A(\us30\/_0097_ ), .B(\us30\/_0122_ ), .C(\us30\/_0149_ ), .D(\us30\/_0167_ ), .X(\us30\/_0168_ ) );
sky130_fd_sc_hd__and2_1 \us30/_0982_ ( .A(\us30\/_0662_ ), .B(\us30\/_0150_ ), .X(\us30\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_0983_ ( .A(\us30\/_0154_ ), .B(\us30\/_0169_ ), .Y(\us30\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us30/_0984_ ( .A(\us30\/_0123_ ), .B(\us30\/_0151_ ), .C(\us30\/_0038_ ), .X(\us30\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0985_ ( .A(\us30\/_0170_ ), .B(\us30\/_0171_ ), .X(\us30\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \us30/_0986_ ( .A(\us30\/_0172_ ), .Y(\us30\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \us30/_0987_ ( .A(\us30\/_0067_ ), .B(\us30\/_0168_ ), .C(\us30\/_0174_ ), .Y(\us30\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us30/_0988_ ( .A(\sa30\[1\] ), .B(\sa30\[0\] ), .Y(\us30\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us30/_0989_ ( .A(\us30\/_0175_ ), .B(\us30\/_0358_ ), .X(\us30\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0990_ ( .A(\us30\/_0176_ ), .B(\us30\/_0478_ ), .X(\us30\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_0991_ ( .A(\us30\/_0280_ ), .B(\us30\/_0113_ ), .Y(\us30\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0992_ ( .A(\us30\/_0111_ ), .B(\us30\/_0062_ ), .X(\us30\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0993_ ( .A(\us30\/_0111_ ), .B(\us30\/_0662_ ), .X(\us30\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_0994_ ( .A(\us30\/_0179_ ), .B(\us30\/_0180_ ), .Y(\us30\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0995_ ( .A(\us30\/_0054_ ), .B(\us30\/_0058_ ), .X(\us30\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us30/_0996_ ( .A(\us30\/_0182_ ), .Y(\us30\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us30/_0997_ ( .A_N(\us30\/_0177_ ), .B(\us30\/_0178_ ), .C(\us30\/_0181_ ), .D(\us30\/_0184_ ), .X(\us30\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0998_ ( .A(\us30\/_0098_ ), .B(\us30\/_0741_ ), .X(\us30\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us30/_0999_ ( .A(\us30\/_0047_ ), .B(\us30\/_0098_ ), .X(\us30\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us30/_1000_ ( .A(\us30\/_0186_ ), .B(\us30\/_0187_ ), .X(\us30\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1001_ ( .A(\us30\/_0188_ ), .Y(\us30\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1002_ ( .A(\us30\/_0738_ ), .B(\us30\/_0735_ ), .X(\us30\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1003_ ( .A(\us30\/_0271_ ), .B(\us30\/_0736_ ), .X(\us30\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_1004_ ( .A(\us30\/_0190_ ), .B(\us30\/_0191_ ), .Y(\us30\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us30/_1005_ ( .A(\us30\/_0096_ ), .B(\us30\/_0325_ ), .X(\us30\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1006_ ( .A1(\us30\/_0193_ ), .A2(\us30\/_0176_ ), .B1(\us30\/_0043_ ), .Y(\us30\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1007_ ( .A(\us30\/_0185_ ), .B(\us30\/_0189_ ), .C(\us30\/_0192_ ), .D(\us30\/_0195_ ), .X(\us30\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us30/_1008_ ( .A_N(\sa30\[3\] ), .B(\us30\/_0734_ ), .C(\sa30\[2\] ), .X(\us30\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1009_ ( .A(\us30\/_0137_ ), .B(\us30\/_0197_ ), .X(\us30\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_1010_ ( .A(\us30\/_0198_ ), .B(\us30\/_0040_ ), .Y(\us30\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1011_ ( .A(\us30\/_0293_ ), .B(\us30\/_0137_ ), .X(\us30\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1012_ ( .A(\us30\/_0200_ ), .Y(\us30\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1013_ ( .A(\us30\/_0137_ ), .B(\us30\/_0110_ ), .Y(\us30\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1014_ ( .A(\us30\/_0139_ ), .B(\us30\/_0020_ ), .Y(\us30\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1015_ ( .A(\us30\/_0199_ ), .B(\us30\/_0201_ ), .C(\us30\/_0202_ ), .D(\us30\/_0203_ ), .X(\us30\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us30/_1016_ ( .A1(\us30\/_0532_ ), .A2(\us30\/_0109_ ), .B1(\us30\/_0102_ ), .C1(\us30\/_0727_ ), .X(\us30\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1017_ ( .A(\us30\/_0022_ ), .B(\us30\/_0078_ ), .Y(\us30\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1018_ ( .A(\us30\/_0078_ ), .B(\us30\/_0142_ ), .Y(\us30\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1019_ ( .A(\us30\/_0207_ ), .B(\us30\/_0208_ ), .Y(\us30\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1020_ ( .A1(\us30\/_0094_ ), .A2(\us30\/_0176_ ), .B1(\us30\/_0206_ ), .C1(\us30\/_0209_ ), .Y(\us30\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1021_ ( .A(\us30\/_0662_ ), .B(\us30\/_0070_ ), .X(\us30\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us30/_1022_ ( .A(\us30\/_0731_ ), .B(\us30\/_0123_ ), .C(\us30\/_0749_ ), .Y(\us30\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us30/_1023_ ( .A(\us30\/_0731_ ), .B(\us30\/_0467_ ), .C(\us30\/_0069_ ), .Y(\us30\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us30/_1024_ ( .A_N(\us30\/_0211_ ), .B(\us30\/_0127_ ), .C(\us30\/_0212_ ), .D(\us30\/_0213_ ), .X(\us30\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1025_ ( .A(\us30\/_0137_ ), .Y(\us30\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1026_ ( .A(\us30\/_0128_ ), .B(\us30\/_0035_ ), .Y(\us30\/_0217_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1028_ ( .A1(\us30\/_0159_ ), .A2(\us30\/_0746_ ), .B1(\us30\/_0434_ ), .B2(\us30\/_0499_ ), .Y(\us30\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us30/_1029_ ( .A1(\us30\/_0116_ ), .A2(\us30\/_0215_ ), .B1(\us30\/_0217_ ), .C1(\us30\/_0219_ ), .X(\us30\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1030_ ( .A(\us30\/_0113_ ), .B(\us30\/_0746_ ), .X(\us30\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us30/_1031_ ( .A1(\us30\/_0098_ ), .A2(\us30\/_0746_ ), .B1(\us30\/_0434_ ), .B2(\us30\/_0750_ ), .X(\us30\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1032_ ( .A1(\us30\/_0047_ ), .A2(\us30\/_0113_ ), .B1(\us30\/_0221_ ), .C1(\us30\/_0222_ ), .Y(\us30\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us30/_1033_ ( .A1(\us30\/_0129_ ), .A2(\us30\/_0162_ ), .B1(\us30\/_0271_ ), .B2(\us30\/_0705_ ), .X(\us30\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1034_ ( .A1(\us30\/_0093_ ), .A2(\us30\/_0738_ ), .B1(\us30\/_0081_ ), .C1(\us30\/_0224_ ), .Y(\us30\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1035_ ( .A(\us30\/_0214_ ), .B(\us30\/_0220_ ), .C(\us30\/_0223_ ), .D(\us30\/_0225_ ), .X(\us30\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1036_ ( .A(\us30\/_0196_ ), .B(\us30\/_0204_ ), .C(\us30\/_0210_ ), .D(\us30\/_0226_ ), .X(\us30\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1037_ ( .A(\us30\/_0111_ ), .B(\us30\/_0554_ ), .X(\us30\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1038_ ( .A(\us30\/_0229_ ), .Y(\us30\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1039_ ( .A(\us30\/_0111_ ), .B(\us30\/_0129_ ), .Y(\us30\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1040_ ( .A(\us30\/_0017_ ), .B(\us30\/_0738_ ), .Y(\us30\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1041_ ( .A(\us30\/_0030_ ), .B(\us30\/_0304_ ), .Y(\us30\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1042_ ( .A(\us30\/_0230_ ), .B(\us30\/_0231_ ), .C(\us30\/_0232_ ), .D(\us30\/_0233_ ), .X(\us30\/_0234_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1043_ ( .A(\us30\/_0047_ ), .B(\us30\/_0478_ ), .X(\us30\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1044_ ( .A1(\us30\/_0129_ ), .A2(\us30\/_0554_ ), .B1(\us30\/_0137_ ), .Y(\us30\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us30/_1045_ ( .A(\us30\/_0235_ ), .B(\us30\/_0049_ ), .C_N(\us30\/_0236_ ), .Y(\us30\/_0237_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1046_ ( .A(\us30\/_0047_ ), .B(\us30\/_0077_ ), .X(\us30\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1047_ ( .A(\us30\/_0070_ ), .B(\us30\/_0035_ ), .X(\us30\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us30/_1048_ ( .A1(\us30\/_0047_ ), .A2(\us30\/_0736_ ), .B1(\us30\/_0022_ ), .B2(\us30\/_0099_ ), .X(\us30\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us30/_1049_ ( .A(\us30\/_0239_ ), .B(\us30\/_0240_ ), .C(\us30\/_0241_ ), .Y(\us30\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1050_ ( .A(\us30\/_0554_ ), .B(\us30\/_0072_ ), .X(\us30\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us30/_1051_ ( .A1(\us30\/_0142_ ), .A2(\us30\/_0137_ ), .B1(\us30\/_0159_ ), .B2(\us30\/_0082_ ), .X(\us30\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1052_ ( .A1(\us30\/_0608_ ), .A2(\us30\/_0072_ ), .B1(\us30\/_0243_ ), .C1(\us30\/_0244_ ), .Y(\us30\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1053_ ( .A(\us30\/_0234_ ), .B(\us30\/_0237_ ), .C(\us30\/_0242_ ), .D(\us30\/_0245_ ), .X(\us30\/_0246_ ) );
sky130_fd_sc_hd__buf_2 \us30/_1054_ ( .A(\us30\/_0027_ ), .X(\us30\/_0247_ ) );
sky130_fd_sc_hd__o21a_1 \us30/_1055_ ( .A1(\us30\/_0554_ ), .A2(\us30\/_0586_ ), .B1(\us30\/_0247_ ), .X(\us30\/_0248_ ) );
sky130_fd_sc_hd__and2_1 \us30/_1056_ ( .A(\us30\/_0082_ ), .B(\us30\/_0478_ ), .X(\us30\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_1057_ ( .A(\us30\/_0079_ ), .X(\us30\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1058_ ( .A(\us30\/_0251_ ), .B(\us30\/_0478_ ), .X(\us30\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_1059_ ( .A(\us30\/_0250_ ), .B(\us30\/_0252_ ), .Y(\us30\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1060_ ( .A(\us30\/_0016_ ), .B(\us30\/_0064_ ), .Y(\us30\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_1061_ ( .A(\us30\/_0304_ ), .X(\us30\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1062_ ( .A(\us30\/_0255_ ), .B(\us30\/_0640_ ), .Y(\us30\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us30/_1063_ ( .A_N(\us30\/_0248_ ), .B(\us30\/_0253_ ), .C(\us30\/_0254_ ), .D(\us30\/_0256_ ), .X(\us30\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1064_ ( .A(\us30\/_0099_ ), .B(\us30\/_0110_ ), .X(\us30\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us30/_1065_ ( .A1(\us30\/_0161_ ), .A2(\us30\/_0130_ ), .B1(\us30\/_0258_ ), .Y(\us30\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1066_ ( .A(\us30\/_0194_ ), .B(\sa30\[1\] ), .X(\us30\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1068_ ( .A(\us30\/_0261_ ), .B(\us30\/_0153_ ), .Y(\us30\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us30/_1069_ ( .A_N(\us30\/_0154_ ), .B(\us30\/_0259_ ), .C(\us30\/_0263_ ), .X(\us30\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1070_ ( .A(\us30\/_0246_ ), .B(\us30\/_0174_ ), .C(\us30\/_0257_ ), .D(\us30\/_0264_ ), .X(\us30\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us30/_1071_ ( .A1(\us30\/_0261_ ), .A2(\us30\/_0554_ ), .B1(\us30\/_0159_ ), .X(\us30\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1072_ ( .A(\us30\/_0746_ ), .B(\us30\/_0150_ ), .Y(\us30\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1073_ ( .A(\us30\/_0175_ ), .Y(\us30\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us30/_1074_ ( .A(\us30\/_0412_ ), .B(\us30\/_0123_ ), .C(\us30\/_0151_ ), .X(\us30\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1075_ ( .A(\us30\/_0268_ ), .B(\us30\/_0269_ ), .Y(\us30\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us30/_1076_ ( .A_N(\us30\/_0266_ ), .B(\us30\/_0267_ ), .C(\us30\/_0270_ ), .X(\us30\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1077_ ( .A(\us30\/_0554_ ), .B(\us30\/_0150_ ), .X(\us30\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1078_ ( .A(\us30\/_0273_ ), .Y(\us30\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1079_ ( .A1(\us30\/_0734_ ), .A2(\us30\/_0325_ ), .B1(\us30\/_0380_ ), .Y(\us30\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1080_ ( .A(\us30\/_0275_ ), .Y(\us30\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1081_ ( .A(\us30\/_0276_ ), .B(\us30\/_0153_ ), .Y(\us30\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us30/_1082_ ( .A(\us30\/_0272_ ), .B(\us30\/_0274_ ), .C(\us30\/_0277_ ), .X(\us30\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_1083_ ( .A(\us30\/_0035_ ), .X(\us30\/_0279_ ) );
sky130_fd_sc_hd__buf_2 \us30/_1084_ ( .A(\us30\/_0082_ ), .X(\us30\/_0280_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1085_ ( .A1(\us30\/_0499_ ), .A2(\us30\/_0279_ ), .B1(\us30\/_0280_ ), .B2(\us30\/_0060_ ), .Y(\us30\/_0281_ ) );
sky130_fd_sc_hd__o21ai_1 \us30/_1086_ ( .A1(\us30\/_0251_ ), .A2(\us30\/_0434_ ), .B1(\us30\/_0304_ ), .Y(\us30\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1087_ ( .A(\us30\/_0091_ ), .B(\us30\/_0292_ ), .Y(\us30\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1088_ ( .A1(\us30\/_0118_ ), .A2(\us30\/_0050_ ), .B1(\us30\/_0038_ ), .C1(\us30\/_0255_ ), .Y(\us30\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1089_ ( .A(\us30\/_0281_ ), .B(\us30\/_0283_ ), .C(\us30\/_0284_ ), .D(\us30\/_0285_ ), .X(\us30\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1090_ ( .A(\us30\/_0082_ ), .B(\us30\/_0027_ ), .X(\us30\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1091_ ( .A(\us30\/_0129_ ), .B(\us30\/_0027_ ), .X(\us30\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_1092_ ( .A(\us30\/_0287_ ), .B(\us30\/_0288_ ), .Y(\us30\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1093_ ( .A1(\us30\/_0752_ ), .A2(\us30\/_0683_ ), .B1(\us30\/_0093_ ), .B2(\us30\/_0247_ ), .Y(\us30\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1094_ ( .A1(\us30\/_0092_ ), .A2(\us30\/_0575_ ), .B1(\us30\/_0292_ ), .Y(\us30\/_0291_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_1095_ ( .A(\us30\/_0054_ ), .X(\us30\/_0292_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1096_ ( .A1(\us30\/_0499_ ), .A2(\us30\/_0662_ ), .B1(\us30\/_0280_ ), .B2(\us30\/_0292_ ), .Y(\us30\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1097_ ( .A(\us30\/_0289_ ), .B(\us30\/_0290_ ), .C(\us30\/_0291_ ), .D(\us30\/_0294_ ), .X(\us30\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1098_ ( .A(\us30\/_0750_ ), .B(\us30\/_0193_ ), .X(\us30\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1099_ ( .A(\us30\/_0705_ ), .B(\us30\/_0380_ ), .X(\us30\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1100_ ( .A(\us30\/_0752_ ), .B(\us30\/_0129_ ), .Y(\us30\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us30/_1101_ ( .A(\us30\/_0296_ ), .B(\us30\/_0297_ ), .C_N(\us30\/_0298_ ), .Y(\us30\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1102_ ( .A(\us30\/_0089_ ), .B(\us30\/_0532_ ), .Y(\us30\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1103_ ( .A(\sa30\[2\] ), .Y(\us30\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \us30/_1104_ ( .A(\us30\/_0301_ ), .B(\sa30\[3\] ), .C(\us30\/_0118_ ), .Y(\us30\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1105_ ( .A(\us30\/_0072_ ), .B(\us30\/_0302_ ), .X(\us30\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1106_ ( .A(\us30\/_0303_ ), .Y(\us30\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1107_ ( .A(\us30\/_0147_ ), .B(\us30\/_0302_ ), .Y(\us30\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1108_ ( .A(\us30\/_0299_ ), .B(\us30\/_0300_ ), .C(\us30\/_0305_ ), .D(\us30\/_0306_ ), .X(\us30\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1109_ ( .A(\us30\/_0278_ ), .B(\us30\/_0286_ ), .C(\us30\/_0295_ ), .D(\us30\/_0307_ ), .X(\us30\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us30/_1110_ ( .A(\us30\/_0228_ ), .B(\us30\/_0265_ ), .C(\us30\/_0308_ ), .Y(\us30\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1111_ ( .A(\us30\/_0235_ ), .Y(\us30\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1112_ ( .A(\us30\/_0478_ ), .B(\us30\/_0640_ ), .X(\us30\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1113_ ( .A(\us30\/_0310_ ), .Y(\us30\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1114_ ( .A(\us30\/_0022_ ), .B(\us30\/_0499_ ), .Y(\us30\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1115_ ( .A(\us30\/_0499_ ), .B(\us30\/_0032_ ), .Y(\us30\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1116_ ( .A(\us30\/_0309_ ), .B(\us30\/_0311_ ), .C(\us30\/_0312_ ), .D(\us30\/_0313_ ), .X(\us30\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1117_ ( .A(\us30\/_0499_ ), .B(\us30\/_0064_ ), .Y(\us30\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1118_ ( .A(\us30\/_0499_ ), .B(\us30\/_0683_ ), .Y(\us30\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1119_ ( .A(\us30\/_0315_ ), .B(\us30\/_0316_ ), .C(\us30\/_0317_ ), .D(\us30\/_0253_ ), .X(\us30\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1120_ ( .A(\us30\/_0047_ ), .B(\us30\/_0304_ ), .Y(\us30\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1121_ ( .A(\us30\/_0586_ ), .B(\us30\/_0162_ ), .Y(\us30\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1122_ ( .A(\us30\/_0319_ ), .B(\us30\/_0320_ ), .Y(\us30\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_1123_ ( .A(\us30\/_0321_ ), .B(\us30\/_0238_ ), .Y(\us30\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1124_ ( .A(\us30\/_0304_ ), .B(\us30\/_0062_ ), .Y(\us30\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_1125_ ( .A(\us30\/_0251_ ), .X(\us30\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1126_ ( .A1(\us30\/_0324_ ), .A2(\us30\/_0280_ ), .B1(\us30\/_0255_ ), .Y(\us30\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1127_ ( .A1(\us30\/_0050_ ), .A2(\us30\/_0205_ ), .B1(\us30\/_0109_ ), .C1(\us30\/_0255_ ), .Y(\us30\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1128_ ( .A(\us30\/_0322_ ), .B(\us30\/_0323_ ), .C(\us30\/_0326_ ), .D(\us30\/_0327_ ), .X(\us30\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1129_ ( .A1(\us30\/_0733_ ), .A2(\us30\/_0279_ ), .A3(\us30\/_0058_ ), .B1(\us30\/_0292_ ), .Y(\us30\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_1130_ ( .A(\us30\/_0047_ ), .X(\us30\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1131_ ( .A(\us30\/_0330_ ), .B(\us30\/_0292_ ), .Y(\us30\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1132_ ( .A(\us30\/_0054_ ), .B(\us30\/_0045_ ), .Y(\us30\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1133_ ( .A(\us30\/_0329_ ), .B(\us30\/_0331_ ), .C(\us30\/_0284_ ), .D(\us30\/_0332_ ), .X(\us30\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us30/_1134_ ( .A1(\us30\/_0249_ ), .A2(\us30\/_0205_ ), .B1(\us30\/_0532_ ), .C1(\us30\/_0060_ ), .X(\us30\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1135_ ( .A(\us30\/_0280_ ), .B(\us30\/_0060_ ), .Y(\us30\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1136_ ( .A(\us30\/_0324_ ), .B(\us30\/_0060_ ), .Y(\us30\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1137_ ( .A(\us30\/_0335_ ), .B(\us30\/_0337_ ), .Y(\us30\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1138_ ( .A1(\us30\/_0276_ ), .A2(\us30\/_0060_ ), .B1(\us30\/_0334_ ), .C1(\us30\/_0338_ ), .Y(\us30\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1139_ ( .A(\us30\/_0318_ ), .B(\us30\/_0328_ ), .C(\us30\/_0333_ ), .D(\us30\/_0339_ ), .X(\us30\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us30/_1140_ ( .A1(\us30\/_0746_ ), .A2(\us30\/_0134_ ), .B1(\us30\/_0128_ ), .X(\us30\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us30/_1141_ ( .A_N(\us30\/_0086_ ), .B(\us30\/_0128_ ), .X(\us30\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1142_ ( .A(\us30\/_0079_ ), .B(\us30\/_0124_ ), .X(\us30\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_1143_ ( .A(\us30\/_0126_ ), .B(\us30\/_0343_ ), .Y(\us30\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us30/_1144_ ( .A(\us30\/_0341_ ), .B(\us30\/_0342_ ), .C_N(\us30\/_0344_ ), .Y(\us30\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1146_ ( .A1(\us30\/_0193_ ), .A2(\us30\/_0092_ ), .A3(\us30\/_0330_ ), .B1(\us30\/_0147_ ), .Y(\us30\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1147_ ( .A1(\us30\/_0130_ ), .A2(\us30\/_0280_ ), .A3(\us30\/_0134_ ), .B1(\us30\/_0139_ ), .Y(\us30\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1148_ ( .A1(\us30\/_0144_ ), .A2(\us30\/_0608_ ), .A3(\us30\/_0092_ ), .B1(\us30\/_0139_ ), .Y(\us30\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1149_ ( .A(\us30\/_0345_ ), .B(\us30\/_0348_ ), .C(\us30\/_0349_ ), .D(\us30\/_0350_ ), .X(\us30\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us30/_1150_ ( .A(\us30\/_0150_ ), .B(\us30\/_0194_ ), .C(\us30\/_0249_ ), .X(\us30\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us30/_1151_ ( .A(\us30\/_0277_ ), .SLEEP(\us30\/_0352_ ), .X(\us30\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us30/_1152_ ( .A1(\us30\/_0268_ ), .A2(\us30\/_0171_ ), .B1(\us30\/_0157_ ), .Y(\us30\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us30/_1153_ ( .A(\us30\/_0161_ ), .X(\us30\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1154_ ( .A1(\us30\/_0279_ ), .A2(\us30\/_0280_ ), .B1(\us30\/_0355_ ), .Y(\us30\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1155_ ( .A1(\us30\/_0020_ ), .A2(\us30\/_0193_ ), .A3(\us30\/_0091_ ), .B1(\us30\/_0355_ ), .Y(\us30\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1156_ ( .A(\us30\/_0353_ ), .B(\us30\/_0354_ ), .C(\us30\/_0356_ ), .D(\us30\/_0357_ ), .X(\us30\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1157_ ( .A(\us30\/_0111_ ), .B(\us30\/_0586_ ), .X(\us30\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1158_ ( .A(\us30\/_0360_ ), .Y(\us30\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us30/_1159_ ( .A1(\us30\/_0119_ ), .A2(\us30\/_0120_ ), .B1(\us30\/_0230_ ), .C1(\us30\/_0361_ ), .X(\us30\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1160_ ( .A1(\us30\/_0662_ ), .A2(\us30\/_0251_ ), .A3(\us30\/_0134_ ), .B1(\us30\/_0114_ ), .Y(\us30\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1162_ ( .A1(\us30\/_0035_ ), .A2(\us30\/_0251_ ), .A3(\us30\/_0134_ ), .B1(\us30\/_0099_ ), .Y(\us30\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1163_ ( .A1(\us30\/_0193_ ), .A2(\us30\/_0608_ ), .B1(\us30\/_0099_ ), .Y(\us30\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1164_ ( .A(\us30\/_0362_ ), .B(\us30\/_0363_ ), .C(\us30\/_0365_ ), .D(\us30\/_0366_ ), .X(\us30\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1165_ ( .A1(\us30\/_0575_ ), .A2(\us30\/_0092_ ), .A3(\us30\/_0330_ ), .B1(\us30\/_0089_ ), .Y(\us30\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1166_ ( .A1(\us30\/_0586_ ), .A2(\us30\/_0017_ ), .A3(\us30\/_0330_ ), .B1(\us30\/_0094_ ), .Y(\us30\/_0370_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1167_ ( .A1(\us30\/_0293_ ), .A2(\us30\/_0134_ ), .B1(\us30\/_0089_ ), .Y(\us30\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1168_ ( .A1(\us30\/_0279_ ), .A2(\us30\/_0134_ ), .B1(\us30\/_0094_ ), .Y(\us30\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1169_ ( .A(\us30\/_0368_ ), .B(\us30\/_0370_ ), .C(\us30\/_0371_ ), .D(\us30\/_0372_ ), .X(\us30\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1170_ ( .A(\us30\/_0351_ ), .B(\us30\/_0359_ ), .C(\us30\/_0367_ ), .D(\us30\/_0373_ ), .X(\us30\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1171_ ( .A1(\us30\/_0102_ ), .A2(\us30\/_0347_ ), .B1(\us30\/_0109_ ), .C1(\us30\/_0247_ ), .Y(\us30\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1172_ ( .A1(\us30\/_0102_ ), .A2(\us30\/_0347_ ), .B1(\us30\/_0532_ ), .C1(\us30\/_0247_ ), .Y(\us30\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1173_ ( .A1(\us30\/_0050_ ), .A2(\us30\/_0249_ ), .B1(\us30\/_0380_ ), .C1(\us30\/_0247_ ), .Y(\us30\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1174_ ( .A(\us30\/_0041_ ), .B(\us30\/_0375_ ), .C(\us30\/_0376_ ), .D(\us30\/_0377_ ), .X(\us30\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1175_ ( .A(\us30\/_0047_ ), .B(\us30\/_0750_ ), .X(\us30\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1176_ ( .A(\us30\/_0379_ ), .Y(\us30\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1177_ ( .A(\us30\/_0016_ ), .B(\us30\/_0608_ ), .Y(\us30\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1178_ ( .A(\us30\/_0752_ ), .B(\us30\/_0554_ ), .Y(\us30\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1179_ ( .A1(\sa30\[1\] ), .A2(\us30\/_0734_ ), .B1(\us30\/_0109_ ), .C1(\us30\/_0016_ ), .Y(\us30\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1180_ ( .A(\us30\/_0381_ ), .B(\us30\/_0382_ ), .C(\us30\/_0383_ ), .D(\us30\/_0384_ ), .X(\us30\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us30/_1181_ ( .A(\us30\/_0086_ ), .B_N(\us30\/_0736_ ), .X(\us30\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1182_ ( .A1(\us30\/_0748_ ), .A2(\us30\/_0134_ ), .B1(\us30\/_0739_ ), .Y(\us30\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1183_ ( .A1(\us30\/_0118_ ), .A2(\us30\/_0249_ ), .B1(\us30\/_0109_ ), .C1(\us30\/_0739_ ), .Y(\us30\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1184_ ( .A1(\us30\/_0102_ ), .A2(\us30\/_0301_ ), .B1(\sa30\[3\] ), .C1(\us30\/_0739_ ), .Y(\us30\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1185_ ( .A(\us30\/_0386_ ), .B(\us30\/_0387_ ), .C(\us30\/_0388_ ), .D(\us30\/_0389_ ), .X(\us30\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1186_ ( .A(\us30\/_0020_ ), .Y(\us30\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1187_ ( .A(\us30\/_0727_ ), .Y(\us30\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1188_ ( .A(\us30\/_0727_ ), .B(\us30\/_0064_ ), .Y(\us30\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1189_ ( .A1(\us30\/_0102_ ), .A2(\us30\/_0734_ ), .B1(\us30\/_0532_ ), .C1(\us30\/_0727_ ), .Y(\us30\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us30/_1190_ ( .A1(\us30\/_0392_ ), .A2(\us30\/_0393_ ), .B1(\us30\/_0394_ ), .C1(\us30\/_0395_ ), .X(\us30\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1191_ ( .A(\us30\/_0378_ ), .B(\us30\/_0385_ ), .C(\us30\/_0390_ ), .D(\us30\/_0396_ ), .X(\us30\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us30/_1192_ ( .A(\us30\/_0340_ ), .B(\us30\/_0374_ ), .C(\us30\/_0397_ ), .Y(\us30\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1193_ ( .A(\us30\/_0077_ ), .B(\us30\/_0129_ ), .X(\us30\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_1194_ ( .A(\us30\/_0398_ ), .B(\us30\/_0239_ ), .Y(\us30\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1195_ ( .A(\us30\/_0022_ ), .B(\us30\/_0111_ ), .X(\us30\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us30/_1196_ ( .A_N(\us30\/_0400_ ), .B(\us30\/_0231_ ), .Y(\us30\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us30/_1197_ ( .A(\us30\/_0399_ ), .SLEEP(\us30\/_0402_ ), .X(\us30\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_1198_ ( .A(\us30\/_0746_ ), .B(\us30\/_0251_ ), .Y(\us30\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us30/_1199_ ( .A_N(\us30\/_0404_ ), .B(\us30\/_0752_ ), .Y(\us30\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us30/_1200_ ( .A(\us30\/_0467_ ), .B(\us30\/_0194_ ), .C(\us30\/_0694_ ), .X(\us30\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us30/_1201_ ( .A_N(\us30\/_0175_ ), .B(\us30\/_0406_ ), .X(\us30\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1202_ ( .A(\us30\/_0407_ ), .Y(\us30\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1203_ ( .A1(\us30\/_0094_ ), .A2(\us30\/_0197_ ), .B1(\us30\/_0114_ ), .B2(\us30\/_0640_ ), .Y(\us30\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1204_ ( .A(\us30\/_0403_ ), .B(\us30\/_0405_ ), .C(\us30\/_0408_ ), .D(\us30\/_0409_ ), .X(\us30\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1205_ ( .A(\us30\/_0030_ ), .B(\us30\/_0150_ ), .Y(\us30\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us30/_1206_ ( .A_N(\us30\/_0169_ ), .B(\us30\/_0289_ ), .C(\us30\/_0411_ ), .X(\us30\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us30/_1207_ ( .A1(\us30\/_0467_ ), .A2(\us30\/_0151_ ), .B1(\us30\/_0140_ ), .C1(\us30\/_0129_ ), .X(\us30\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1208_ ( .A1(\us30\/_0608_ ), .A2(\us30\/_0099_ ), .B1(\us30\/_0037_ ), .C1(\us30\/_0414_ ), .Y(\us30\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1209_ ( .A(\us30\/_0738_ ), .Y(\us30\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1210_ ( .A(\us30\/_0586_ ), .B(\us30\/_0736_ ), .Y(\us30\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1211_ ( .A1(\us30\/_0194_ ), .A2(\us30\/_0038_ ), .B1(\us30\/_0118_ ), .C1(\us30\/_0153_ ), .Y(\us30\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us30/_1212_ ( .A1(\us30\/_0416_ ), .A2(\us30\/_0117_ ), .B1(\us30\/_0417_ ), .C1(\us30\/_0418_ ), .X(\us30\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1213_ ( .A(\us30\/_0077_ ), .B(\us30\/_0035_ ), .X(\us30\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1214_ ( .A(\us30\/_0662_ ), .B(\us30\/_0124_ ), .Y(\us30\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1215_ ( .A(\us30\/_0030_ ), .B(\us30\/_0137_ ), .Y(\us30\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1216_ ( .A(\us30\/_0072_ ), .B(\us30\/_0731_ ), .Y(\us30\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us30/_1217_ ( .A_N(\us30\/_0420_ ), .B(\us30\/_0421_ ), .C(\us30\/_0422_ ), .D(\us30\/_0424_ ), .X(\us30\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1218_ ( .A(\us30\/_0413_ ), .B(\us30\/_0415_ ), .C(\us30\/_0419_ ), .D(\us30\/_0425_ ), .X(\us30\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us30/_1219_ ( .A(\us30\/_0355_ ), .B(\us30\/_0102_ ), .C(\us30\/_0109_ ), .Y(\us30\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1220_ ( .A(\us30\/_0077_ ), .B(\us30\/_0017_ ), .X(\us30\/_0428_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1221_ ( .A(\us30\/_0077_ ), .B(\us30\/_0554_ ), .X(\us30\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us30/_1222_ ( .A1(\us30\/_0050_ ), .A2(\us30\/_0205_ ), .B1(\us30\/_0380_ ), .C1(\us30\/_0078_ ), .X(\us30\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us30/_1223_ ( .A(\us30\/_0428_ ), .B(\us30\/_0429_ ), .C(\us30\/_0430_ ), .Y(\us30\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us30/_1224_ ( .A_N(\us30\/_0209_ ), .B(\us30\/_0431_ ), .X(\us30\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us30/_1225_ ( .A1(\us30\/_0215_ ), .A2(\us30\/_0404_ ), .B1(\us30\/_0427_ ), .C1(\us30\/_0432_ ), .X(\us30\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1226_ ( .A(\us30\/_0043_ ), .B(\us30\/_0058_ ), .Y(\us30\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1227_ ( .A(\us30\/_0195_ ), .B(\us30\/_0233_ ), .C(\us30\/_0320_ ), .D(\us30\/_0435_ ), .X(\us30\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1228_ ( .A(\us30\/_0261_ ), .B(\us30\/_0738_ ), .Y(\us30\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1229_ ( .A1(\us30\/_0499_ ), .A2(\us30\/_0640_ ), .B1(\us30\/_0261_ ), .B2(\us30\/_0292_ ), .Y(\us30\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1230_ ( .A(\us30\/_0436_ ), .B(\us30\/_0394_ ), .C(\us30\/_0437_ ), .D(\us30\/_0438_ ), .X(\us30\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1231_ ( .A(\us30\/_0410_ ), .B(\us30\/_0426_ ), .C(\us30\/_0433_ ), .D(\us30\/_0439_ ), .X(\us30\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us30/_1232_ ( .A(\us30\/_0135_ ), .SLEEP(\us30\/_0273_ ), .X(\us30\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1233_ ( .A1(\us30\/_0279_ ), .A2(\us30\/_0134_ ), .B1(\us30\/_0099_ ), .Y(\us30\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1234_ ( .A(\us30\/_0441_ ), .B(\us30\/_0164_ ), .C(\us30\/_0270_ ), .D(\us30\/_0442_ ), .X(\us30\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1235_ ( .A(\us30\/_0051_ ), .B(\us30\/_0662_ ), .Y(\us30\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1236_ ( .A(\us30\/_0051_ ), .B(\us30\/_0271_ ), .Y(\us30\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1237_ ( .A(\us30\/_0444_ ), .B(\us30\/_0446_ ), .X(\us30\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1238_ ( .A(\us30\/_0193_ ), .B(\us30\/_0304_ ), .X(\us30\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1239_ ( .A(\us30\/_0448_ ), .Y(\us30\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1240_ ( .A(\us30\/_0162_ ), .B(\us30\/_0130_ ), .X(\us30\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1241_ ( .A(\us30\/_0450_ ), .Y(\us30\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1242_ ( .A1(\us30\/_0129_ ), .A2(\us30\/_0554_ ), .B1(\us30\/_0043_ ), .Y(\us30\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1243_ ( .A(\us30\/_0447_ ), .B(\us30\/_0449_ ), .C(\us30\/_0451_ ), .D(\us30\/_0452_ ), .X(\us30\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1244_ ( .A(\us30\/_0292_ ), .B(\us30\/_0064_ ), .Y(\us30\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us30/_1245_ ( .A_N(\us30\/_0248_ ), .B(\us30\/_0454_ ), .C(\us30\/_0254_ ), .D(\us30\/_0256_ ), .X(\us30\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1246_ ( .A1(\us30\/_0330_ ), .A2(\us30\/_0099_ ), .B1(\us30\/_0134_ ), .B2(\us30\/_0705_ ), .Y(\us30\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1247_ ( .A1(\us30\/_0748_ ), .A2(\us30\/_0738_ ), .B1(\us30\/_0092_ ), .B2(\us30\/_0752_ ), .Y(\us30\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1248_ ( .A1(\us30\/_0072_ ), .A2(\us30\/_0035_ ), .B1(\us30\/_0748_ ), .B2(\us30\/_0292_ ), .Y(\us30\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1249_ ( .A1(\us30\/_0748_ ), .A2(\us30\/_0251_ ), .B1(\us30\/_0247_ ), .Y(\us30\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1250_ ( .A(\us30\/_0457_ ), .B(\us30\/_0458_ ), .C(\us30\/_0459_ ), .D(\us30\/_0460_ ), .X(\us30\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1251_ ( .A(\us30\/_0443_ ), .B(\us30\/_0453_ ), .C(\us30\/_0455_ ), .D(\us30\/_0461_ ), .X(\us30\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1252_ ( .A(\us30\/_0705_ ), .B(\us30\/_0079_ ), .X(\us30\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1253_ ( .A(\us30\/_0586_ ), .B(\us30\/_0124_ ), .Y(\us30\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1254_ ( .A(\us30\/_0499_ ), .B(\us30\/_0746_ ), .Y(\us30\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us30/_1255_ ( .A_N(\us30\/_0463_ ), .B(\us30\/_0464_ ), .C(\us30\/_0465_ ), .X(\us30\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us30/_1256_ ( .A1(\us30\/_0271_ ), .A2(\us30\/_0072_ ), .B1(\us30\/_0142_ ), .B2(\us30\/_0027_ ), .X(\us30\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1257_ ( .A1(\us30\/_0144_ ), .A2(\us30\/_0099_ ), .B1(\us30\/_0360_ ), .C1(\us30\/_0468_ ), .Y(\us30\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us30/_1258_ ( .A1(\us30\/_0662_ ), .A2(\us30\/_0251_ ), .B1(\us30\/_0499_ ), .X(\us30\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1259_ ( .A1(\us30\/_0575_ ), .A2(\us30\/_0292_ ), .B1(\us30\/_0379_ ), .C1(\us30\/_0470_ ), .Y(\us30\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1260_ ( .A(\us30\/_0466_ ), .B(\us30\/_0469_ ), .C(\us30\/_0471_ ), .D(\us30\/_0305_ ), .X(\us30\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us30/_1261_ ( .A1(\us30\/_0247_ ), .A2(\us30\/_0683_ ), .B1(\us30\/_0324_ ), .B2(\us30\/_0292_ ), .X(\us30\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1262_ ( .A(\us30\/_0280_ ), .B(\us30\/_0099_ ), .X(\us30\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us30/_1263_ ( .A1(\us30\/_0092_ ), .A2(\us30\/_0247_ ), .B1(\us30\/_0474_ ), .X(\us30\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us30/_1264_ ( .A(\us30\/_0075_ ), .B(\us30\/_0473_ ), .C(\us30\/_0475_ ), .Y(\us30\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1265_ ( .A1(\us30\/_0279_ ), .A2(\us30\/_0255_ ), .B1(\us30\/_0280_ ), .B2(\us30\/_0060_ ), .Y(\us30\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1266_ ( .A1(\us30\/_0093_ ), .A2(\us30\/_0292_ ), .B1(\us30\/_0134_ ), .B2(\us30\/_0114_ ), .Y(\us30\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1267_ ( .A1(\us30\/_0161_ ), .A2(\us30\/_0032_ ), .B1(\us30\/_0324_ ), .B2(\us30\/_0147_ ), .Y(\us30\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1268_ ( .A1(\us30\/_0054_ ), .A2(\us30\/_0731_ ), .B1(\us30\/_0748_ ), .B2(\us30\/_0304_ ), .Y(\us30\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1269_ ( .A(\us30\/_0477_ ), .B(\us30\/_0479_ ), .C(\us30\/_0480_ ), .D(\us30\/_0481_ ), .X(\us30\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1270_ ( .A(\us30\/_0161_ ), .B(\us30\/_0064_ ), .Y(\us30\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us30/_1271_ ( .A(\us30\/_0731_ ), .B(\us30\/_0123_ ), .C(\us30\/_0467_ ), .Y(\us30\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1272_ ( .A(\us30\/_0483_ ), .B(\us30\/_0484_ ), .Y(\us30\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1273_ ( .A(\us30\/_0297_ ), .Y(\us30\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us30/_1274_ ( .A_N(\us30\/_0485_ ), .B(\us30\/_0181_ ), .C(\us30\/_0486_ ), .D(\us30\/_0386_ ), .X(\us30\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1275_ ( .A(\us30\/_0472_ ), .B(\us30\/_0476_ ), .C(\us30\/_0482_ ), .D(\us30\/_0487_ ), .X(\us30\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \us30/_1276_ ( .A(\us30\/_0440_ ), .B(\us30\/_0462_ ), .C(\us30\/_0488_ ), .Y(\us30\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1277_ ( .A(\us30\/_0403_ ), .B(\us30\/_0230_ ), .C(\us30\/_0451_ ), .D(\us30\/_0361_ ), .X(\us30\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1278_ ( .A1(\us30\/_0118_ ), .A2(\us30\/_0050_ ), .B1(\us30\/_0109_ ), .C1(\us30\/_0139_ ), .Y(\us30\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1279_ ( .A(\us30\/_0447_ ), .B(\us30\/_0437_ ), .C(\us30\/_0491_ ), .D(\us30\/_0427_ ), .X(\us30\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1280_ ( .A1(\us30\/_0280_ ), .A2(\us30\/_0255_ ), .B1(\us30\/_0608_ ), .B2(\us30\/_0247_ ), .Y(\us30\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1281_ ( .A1(\us30\/_0144_ ), .A2(\us30\/_0147_ ), .B1(\us30\/_0355_ ), .B2(\us30\/_0093_ ), .Y(\us30\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1282_ ( .A1(\us30\/_0705_ ), .A2(\us30\/_0279_ ), .B1(\us30\/_0330_ ), .B2(\us30\/_0247_ ), .Y(\us30\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1283_ ( .A1(\us30\/_0279_ ), .A2(\us30\/_0280_ ), .B1(\us30\/_0114_ ), .Y(\us30\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1284_ ( .A(\us30\/_0493_ ), .B(\us30\/_0494_ ), .C(\us30\/_0495_ ), .D(\us30\/_0496_ ), .X(\us30\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1285_ ( .A1(\us30\/_0134_ ), .A2(\us30\/_0137_ ), .B1(\us30\/_0355_ ), .B2(\us30\/_0575_ ), .Y(\us30\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1286_ ( .A1(\us30\/_0099_ ), .A2(\us30\/_0733_ ), .B1(\us30\/_0093_ ), .B2(\us30\/_0499_ ), .Y(\us30\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1287_ ( .A(\us30\/_0147_ ), .B(\us30\/_0640_ ), .Y(\us30\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1288_ ( .A1(\us30\/_0153_ ), .A2(\us30\/_0292_ ), .B1(\us30\/_0748_ ), .Y(\us30\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1289_ ( .A(\us30\/_0498_ ), .B(\us30\/_0500_ ), .C(\us30\/_0501_ ), .D(\us30\/_0502_ ), .X(\us30\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1290_ ( .A(\us30\/_0490_ ), .B(\us30\/_0492_ ), .C(\us30\/_0497_ ), .D(\us30\/_0503_ ), .X(\us30\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us30/_1291_ ( .A_N(\us30\/_0275_ ), .B(\us30\/_0705_ ), .X(\us30\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1292_ ( .A(\us30\/_0505_ ), .Y(\us30\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1293_ ( .A(\us30\/_0380_ ), .B(\us30\/_0347_ ), .X(\us30\/_0507_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1294_ ( .A1(\us30\/_0507_ ), .A2(\us30\/_0093_ ), .B1(\us30\/_0292_ ), .Y(\us30\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1295_ ( .A(\us30\/_0322_ ), .B(\us30\/_0277_ ), .C(\us30\/_0506_ ), .D(\us30\/_0508_ ), .X(\us30\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1296_ ( .A(\us30\/_0280_ ), .B(\us30\/_0705_ ), .X(\us30\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1297_ ( .A1(\us30\/_0733_ ), .A2(\us30\/_0114_ ), .B1(\us30\/_0429_ ), .C1(\us30\/_0511_ ), .Y(\us30\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_1298_ ( .A(\us30\/_0019_ ), .B(\us30\/_0024_ ), .Y(\us30\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1299_ ( .A(\us30\/_0512_ ), .B(\us30\/_0513_ ), .C(\us30\/_0742_ ), .D(\us30\/_0306_ ), .X(\us30\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1300_ ( .A1(\us30\/_0532_ ), .A2(\us30\/_0089_ ), .B1(\us30\/_0154_ ), .C1(\us30\/_0169_ ), .Y(\us30\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us30/_1301_ ( .A1(\us30\/_0749_ ), .A2(\us30\/_0026_ ), .B1(\us30\/_0069_ ), .C1(\us30\/_0032_ ), .X(\us30\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us30/_1302_ ( .A1(\us30\/_0324_ ), .A2(\us30\/_0355_ ), .B1(\us30\/_0330_ ), .B2(\us30\/_0727_ ), .X(\us30\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us30/_1303_ ( .A(\us30\/_0133_ ), .B(\us30\/_0516_ ), .C(\us30\/_0517_ ), .Y(\us30\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1304_ ( .A(\us30\/_0509_ ), .B(\us30\/_0514_ ), .C(\us30\/_0515_ ), .D(\us30\/_0518_ ), .X(\us30\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1305_ ( .A(\us30\/_0746_ ), .B(\us30\/_0072_ ), .Y(\us30\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1306_ ( .A1(\us30\/_0082_ ), .A2(\us30\/_0070_ ), .B1(\us30\/_0043_ ), .B2(\us30\/_0193_ ), .Y(\us30\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1307_ ( .A(\us30\/_0311_ ), .B(\us30\/_0520_ ), .C(\us30\/_0332_ ), .D(\us30\/_0522_ ), .X(\us30\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1308_ ( .A(\us30\/_0129_ ), .B(\us30\/_0499_ ), .X(\us30\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_1309_ ( .A(\us30\/_0235_ ), .B(\us30\/_0524_ ), .Y(\us30\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us30/_1310_ ( .A(\us30\/_0081_ ), .B(\us30\/_0085_ ), .Y(\us30\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1311_ ( .A1(\us30\/_0051_ ), .A2(\us30\/_0045_ ), .B1(\us30\/_0130_ ), .B2(\us30\/_0094_ ), .Y(\us30\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1312_ ( .A(\us30\/_0523_ ), .B(\us30\/_0525_ ), .C(\us30\/_0526_ ), .D(\us30\/_0527_ ), .X(\us30\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us30/_1313_ ( .A_N(\us30\/_0250_ ), .B(\us30\/_0521_ ), .Y(\us30\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1314_ ( .A(\us30\/_0128_ ), .B(\us30\/_0020_ ), .X(\us30\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1315_ ( .A(\us30\/_0530_ ), .Y(\us30\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1316_ ( .A(\us30\/_0099_ ), .B(\us30\/_0058_ ), .X(\us30\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1317_ ( .A(\us30\/_0533_ ), .Y(\us30\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us30/_1318_ ( .A_N(\us30\/_0529_ ), .B(\us30\/_0531_ ), .C(\us30\/_0534_ ), .D(\us30\/_0192_ ), .X(\us30\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1319_ ( .A(\us30\/_0434_ ), .B(\us30\/_0078_ ), .X(\us30\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us30/_1320_ ( .A1(\us30\/_0750_ ), .A2(\us30\/_0079_ ), .B1(\us30\/_0129_ ), .B2(\us30\/_0705_ ), .X(\us30\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1321_ ( .A1(\us30\/_0161_ ), .A2(\us30\/_0032_ ), .B1(\us30\/_0536_ ), .C1(\us30\/_0537_ ), .Y(\us30\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us30/_1322_ ( .A1(\us30\/_0746_ ), .A2(\us30\/_0162_ ), .B1(\us30\/_0079_ ), .B2(\us30\/_0043_ ), .X(\us30\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1323_ ( .A1(\us30\/_0093_ ), .A2(\us30\/_0247_ ), .B1(\us30\/_0240_ ), .C1(\us30\/_0539_ ), .Y(\us30\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1324_ ( .A(\us30\/_0434_ ), .B(\us30\/_0043_ ), .X(\us30\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us30/_1325_ ( .A1(\us30\/_0142_ ), .A2(\us30\/_0150_ ), .B1(\us30\/_0022_ ), .B2(\us30\/_0137_ ), .X(\us30\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1326_ ( .A1(\us30\/_0279_ ), .A2(\us30\/_0051_ ), .B1(\us30\/_0541_ ), .C1(\us30\/_0542_ ), .Y(\us30\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1327_ ( .A(\us30\/_0159_ ), .B(\us30\/_0035_ ), .X(\us30\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us30/_1328_ ( .A1(\us30\/_0271_ ), .A2(\us30\/_0434_ ), .B1(\us30\/_0027_ ), .X(\us30\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1329_ ( .A1(\us30\/_0091_ ), .A2(\us30\/_0128_ ), .B1(\us30\/_0545_ ), .C1(\us30\/_0546_ ), .Y(\us30\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1330_ ( .A(\us30\/_0538_ ), .B(\us30\/_0540_ ), .C(\us30\/_0544_ ), .D(\us30\/_0547_ ), .X(\us30\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1331_ ( .A(\us30\/_0099_ ), .B(\us30\/_0193_ ), .X(\us30\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us30/_1332_ ( .A(\us30\/_0549_ ), .B(\us30\/_0186_ ), .C(\us30\/_0187_ ), .Y(\us30\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1333_ ( .A(\us30\/_0062_ ), .B(\us30\/_0347_ ), .C(\us30\/_0749_ ), .D(\us30\/_0694_ ), .X(\us30\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1334_ ( .A1(\us30\/_0130_ ), .A2(\us30\/_0499_ ), .B1(\us30\/_0551_ ), .C1(\us30\/_0101_ ), .Y(\us30\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1335_ ( .A(\us30\/_0139_ ), .B(\us30\/_0640_ ), .Y(\us30\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1336_ ( .A1(\us30\/_0752_ ), .A2(\us30\/_0662_ ), .B1(\us30\/_0280_ ), .B2(\us30\/_0099_ ), .Y(\us30\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1337_ ( .A(\us30\/_0550_ ), .B(\us30\/_0552_ ), .C(\us30\/_0553_ ), .D(\us30\/_0555_ ), .X(\us30\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1338_ ( .A(\us30\/_0528_ ), .B(\us30\/_0535_ ), .C(\us30\/_0548_ ), .D(\us30\/_0556_ ), .X(\us30\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us30/_1339_ ( .A(\us30\/_0504_ ), .B(\us30\/_0519_ ), .C(\us30\/_0557_ ), .Y(\us30\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1340_ ( .A(\us30\/_0054_ ), .B(\us30\/_0507_ ), .X(\us30\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us30/_1341_ ( .A_N(\us30\/_0558_ ), .B(\us30\/_0408_ ), .C(\us30\/_0451_ ), .D(\us30\/_0452_ ), .X(\us30\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1342_ ( .A(\us30\/_0549_ ), .Y(\us30\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1343_ ( .A(\us30\/_0559_ ), .B(\us30\/_0403_ ), .C(\us30\/_0560_ ), .D(\us30\/_0371_ ), .X(\us30\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1344_ ( .A(\us30\/_0181_ ), .B(\us30\/_0178_ ), .X(\us30\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1345_ ( .A(\us30\/_0562_ ), .B(\us30\/_0552_ ), .C(\us30\/_0553_ ), .D(\us30\/_0555_ ), .X(\us30\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1346_ ( .A(\us30\/_0247_ ), .B(\us30\/_0020_ ), .Y(\us30\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1347_ ( .A(\us30\/_0051_ ), .B(\us30\/_0130_ ), .X(\us30\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1348_ ( .A(\us30\/_0566_ ), .Y(\us30\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1349_ ( .A(\us30\/_0159_ ), .B(\us30\/_0412_ ), .X(\us30\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1350_ ( .A1(\us30\/_0752_ ), .A2(\us30\/_0640_ ), .B1(\us30\/_0568_ ), .B2(\us30\/_0175_ ), .Y(\us30\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1351_ ( .A(\us30\/_0076_ ), .B(\us30\/_0565_ ), .C(\us30\/_0567_ ), .D(\us30\/_0569_ ), .X(\us30\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us30/_1352_ ( .A1(\us30\/_0035_ ), .A2(\us30\/_0142_ ), .B1(\us30\/_0161_ ), .X(\us30\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1353_ ( .A(\us30\/_0099_ ), .B(\us30\/_0662_ ), .Y(\us30\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us30/_1354_ ( .A(\us30\/_0420_ ), .B(\us30\/_0571_ ), .C_N(\us30\/_0572_ ), .Y(\us30\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1355_ ( .A(\us30\/_0051_ ), .B(\us30\/_0746_ ), .Y(\us30\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1356_ ( .A(\us30\/_0574_ ), .B(\us30\/_0319_ ), .C(\us30\/_0320_ ), .D(\us30\/_0411_ ), .X(\us30\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1357_ ( .A(\us30\/_0736_ ), .B(\us30\/_0035_ ), .Y(\us30\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1358_ ( .A(\us30\/_0736_ ), .B(\us30\/_0030_ ), .Y(\us30\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1359_ ( .A(\us30\/_0298_ ), .B(\us30\/_0208_ ), .C(\us30\/_0577_ ), .D(\us30\/_0578_ ), .X(\us30\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1360_ ( .A1(\us30\/_0020_ ), .A2(\us30\/_0137_ ), .B1(\us30\/_0261_ ), .B2(\us30\/_0128_ ), .Y(\us30\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1361_ ( .A(\us30\/_0573_ ), .B(\us30\/_0576_ ), .C(\us30\/_0579_ ), .D(\us30\/_0580_ ), .X(\us30\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1362_ ( .A(\us30\/_0561_ ), .B(\us30\/_0563_ ), .C(\us30\/_0570_ ), .D(\us30\/_0581_ ), .X(\us30\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1363_ ( .A(\us30\/_0128_ ), .B(\us30\/_0193_ ), .X(\us30\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1364_ ( .A(\us30\/_0082_ ), .B(\us30\/_0162_ ), .X(\us30\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us30/_1365_ ( .A(\us30\/_0583_ ), .B(\us30\/_0584_ ), .C_N(\us30\/_0437_ ), .Y(\us30\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us30/_1366_ ( .A(\us30\/_0150_ ), .B(\us30\/_0118_ ), .C(\us30\/_0380_ ), .Y(\us30\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us30/_1367_ ( .A_N(\us30\/_0182_ ), .B(\us30\/_0587_ ), .C(\us30\/_0323_ ), .X(\us30\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1368_ ( .A1(\us30\/_0575_ ), .A2(\us30\/_0153_ ), .B1(\us30\/_0727_ ), .B2(\us30\/_0058_ ), .Y(\us30\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1369_ ( .A1(\us30\/_0499_ ), .A2(\us30\/_0064_ ), .B1(\us30\/_0134_ ), .B2(\us30\/_0255_ ), .Y(\us30\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1370_ ( .A(\us30\/_0585_ ), .B(\us30\/_0588_ ), .C(\us30\/_0589_ ), .D(\us30\/_0590_ ), .X(\us30\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us30/_1371_ ( .A1(\us30\/_0091_ ), .A2(\us30\/_0139_ ), .B1(\us30\/_0250_ ), .Y(\us30\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1372_ ( .A1(\us30\/_0092_ ), .A2(\us30\/_0739_ ), .B1(\us30\/_0324_ ), .B2(\us30\/_0247_ ), .Y(\us30\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1373_ ( .A1(\us30\/_0144_ ), .A2(\us30\/_0153_ ), .B1(\us30\/_0683_ ), .B2(\us30\/_0292_ ), .Y(\us30\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1374_ ( .A1(\us30\/_0091_ ), .A2(\us30\/_0499_ ), .B1(\us30\/_0330_ ), .B2(\us30\/_0292_ ), .Y(\us30\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1375_ ( .A(\us30\/_0592_ ), .B(\us30\/_0593_ ), .C(\us30\/_0594_ ), .D(\us30\/_0595_ ), .X(\us30\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1376_ ( .A(\us30\/_0499_ ), .B(\us30\/_0144_ ), .Y(\us30\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1377_ ( .A(\us30\/_0312_ ), .B(\us30\/_0598_ ), .Y(\us30\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1378_ ( .A(\us30\/_0575_ ), .B(\us30\/_0147_ ), .Y(\us30\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1379_ ( .A1(\us30\/_0293_ ), .A2(\us30\/_0137_ ), .B1(\us30\/_0093_ ), .B2(\us30\/_0739_ ), .Y(\us30\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1380_ ( .A1(\us30\/_0734_ ), .A2(\us30\/_0531_ ), .B1(\us30\/_0600_ ), .C1(\us30\/_0601_ ), .Y(\us30\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1381_ ( .A1(\us30\/_0153_ ), .A2(\us30\/_0261_ ), .B1(\us30\/_0599_ ), .C1(\us30\/_0602_ ), .Y(\us30\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1382_ ( .A(\us30\/_0591_ ), .B(\us30\/_0596_ ), .C(\us30\/_0174_ ), .D(\us30\/_0603_ ), .X(\us30\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1383_ ( .A(\us30\/_0247_ ), .B(\us30\/_0144_ ), .Y(\us30\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1384_ ( .A(\us30\/_0113_ ), .B(\us30\/_0017_ ), .Y(\us30\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1385_ ( .A(\us30\/_0381_ ), .B(\us30\/_0605_ ), .C(\us30\/_0361_ ), .D(\us30\/_0606_ ), .X(\us30\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1386_ ( .A1(\us30\/_0016_ ), .A2(\us30\/_0727_ ), .B1(\us30\/_0733_ ), .Y(\us30\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1387_ ( .A1(\us30\/_0586_ ), .A2(\us30\/_0159_ ), .B1(\us30\/_0082_ ), .B2(\us30\/_0750_ ), .Y(\us30\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1388_ ( .A1(\us30\/_0142_ ), .A2(\us30\/_0162_ ), .B1(\us30\/_0079_ ), .B2(\us30\/_0054_ ), .Y(\us30\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1389_ ( .A(\us30\/_0610_ ), .B(\us30\/_0611_ ), .C(\us30\/_0105_ ), .D(\us30\/_0106_ ), .X(\us30\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1390_ ( .A1(\us30\/_0094_ ), .A2(\us30\/_0302_ ), .B1(\us30\/_0324_ ), .B2(\us30\/_0089_ ), .Y(\us30\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1391_ ( .A(\us30\/_0607_ ), .B(\us30\/_0609_ ), .C(\us30\/_0612_ ), .D(\us30\/_0613_ ), .X(\us30\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1392_ ( .A(\us30\/_0041_ ), .B(\us30\/_0170_ ), .X(\us30\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1393_ ( .A(\us30\/_0554_ ), .B(\us30\/_0027_ ), .X(\us30\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1394_ ( .A(\us30\/_0027_ ), .B(\us30\/_0261_ ), .Y(\us30\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us30/_1395_ ( .A_N(\us30\/_0616_ ), .B(\us30\/_0617_ ), .Y(\us30\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1396_ ( .A1(\us30\/_0147_ ), .A2(\us30\/_0302_ ), .B1(\us30\/_0342_ ), .C1(\us30\/_0618_ ), .Y(\us30\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1397_ ( .A(\us30\/_0614_ ), .B(\us30\/_0272_ ), .C(\us30\/_0615_ ), .D(\us30\/_0620_ ), .X(\us30\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us30/_1398_ ( .A(\us30\/_0582_ ), .B(\us30\/_0604_ ), .C(\us30\/_0621_ ), .Y(\us30\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1399_ ( .A1(\us30\/_0280_ ), .A2(\us30\/_0134_ ), .B1(\us30\/_0089_ ), .Y(\us30\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1400_ ( .A1(\us30\/_0144_ ), .A2(\us30\/_0608_ ), .A3(\us30\/_0330_ ), .B1(\us30\/_0089_ ), .Y(\us30\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1401_ ( .A1(\us30\/_0197_ ), .A2(\us30\/_0130_ ), .A3(\us30\/_0110_ ), .B1(\us30\/_0094_ ), .Y(\us30\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1402_ ( .A(\us30\/_0432_ ), .B(\us30\/_0622_ ), .C(\us30\/_0623_ ), .D(\us30\/_0624_ ), .X(\us30\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us30/_1403_ ( .A1(\us30\/_0554_ ), .A2(\us30\/_0017_ ), .A3(\us30\/_0022_ ), .B1(\us30\/_0161_ ), .X(\us30\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us30/_1404_ ( .A_N(\us30\/_0269_ ), .B(\us30\/_0170_ ), .X(\us30\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1405_ ( .A1(\us30\/_0109_ ), .A2(\us30\/_0064_ ), .A3(\us30\/_0733_ ), .B1(\us30\/_0355_ ), .Y(\us30\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us30/_1406_ ( .A_N(\us30\/_0626_ ), .B(\us30\/_0627_ ), .C(\us30\/_0353_ ), .D(\us30\/_0628_ ), .X(\us30\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1407_ ( .A1(\us30\/_0091_ ), .A2(\us30\/_0110_ ), .A3(\us30\/_0176_ ), .B1(\us30\/_0139_ ), .Y(\us30\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1408_ ( .A1(\us30\/_0020_ ), .A2(\us30\/_0261_ ), .B1(\us30\/_0147_ ), .Y(\us30\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1409_ ( .A(\us30\/_0631_ ), .B(\us30\/_0344_ ), .C(\us30\/_0421_ ), .D(\us30\/_0632_ ), .X(\us30\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us30/_1410_ ( .A1(\us30\/_0325_ ), .A2(\us30\/_0734_ ), .B1(\us30\/_0038_ ), .C1(\us30\/_0113_ ), .X(\us30\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1411_ ( .A1(\us30\/_0134_ ), .A2(\us30\/_0114_ ), .B1(\us30\/_0221_ ), .C1(\us30\/_0634_ ), .Y(\us30\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us30/_1412_ ( .A(\us30\/_0119_ ), .B_N(\us30\/_0111_ ), .Y(\us30\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1413_ ( .A1(\us30\/_0032_ ), .A2(\us30\/_0113_ ), .B1(\us30\/_0636_ ), .C1(\us30\/_0400_ ), .Y(\us30\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1414_ ( .A1(\us30\/_0731_ ), .A2(\us30\/_0293_ ), .A3(\us30\/_0251_ ), .B1(\us30\/_0099_ ), .Y(\us30\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1415_ ( .A(\us30\/_0189_ ), .B(\us30\/_0635_ ), .C(\us30\/_0637_ ), .D(\us30\/_0638_ ), .X(\us30\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1416_ ( .A(\us30\/_0625_ ), .B(\us30\/_0630_ ), .C(\us30\/_0633_ ), .D(\us30\/_0639_ ), .X(\us30\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1417_ ( .A(\us30\/_0746_ ), .B(\us30\/_0738_ ), .X(\us30\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1418_ ( .A(\us30\/_0736_ ), .B(\us30\/_0731_ ), .X(\us30\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us30/_1419_ ( .A_N(\us30\/_0643_ ), .B(\us30\/_0577_ ), .Y(\us30\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1420_ ( .A1(\us30\/_0280_ ), .A2(\us30\/_0739_ ), .B1(\us30\/_0642_ ), .C1(\us30\/_0644_ ), .Y(\us30\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1421_ ( .A1(\us30\/_0050_ ), .A2(\us30\/_0249_ ), .B1(\us30\/_0194_ ), .C1(\us30\/_0738_ ), .Y(\us30\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1422_ ( .A(\us30\/_0646_ ), .B(\us30\/_0232_ ), .C(\us30\/_0417_ ), .D(\us30\/_0578_ ), .X(\us30\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1423_ ( .A1(\us30\/_0064_ ), .A2(\us30\/_0733_ ), .B1(\us30\/_0727_ ), .Y(\us30\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1424_ ( .A1(\us30\/_0193_ ), .A2(\us30\/_0276_ ), .B1(\us30\/_0727_ ), .Y(\us30\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1425_ ( .A(\us30\/_0645_ ), .B(\us30\/_0647_ ), .C(\us30\/_0648_ ), .D(\us30\/_0649_ ), .X(\us30\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1426_ ( .A1(\us30\/_0325_ ), .A2(\us30\/_0734_ ), .B1(\us30\/_0038_ ), .C1(\us30\/_0247_ ), .Y(\us30\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1427_ ( .A1(\us30\/_0249_ ), .A2(\us30\/_0205_ ), .B1(\us30\/_0412_ ), .C1(\us30\/_0247_ ), .Y(\us30\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1428_ ( .A(\us30\/_0652_ ), .B(\us30\/_0653_ ), .X(\us30\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1429_ ( .A1(\us30\/_0733_ ), .A2(\us30\/_0748_ ), .A3(\us30\/_0324_ ), .B1(\us30\/_0016_ ), .Y(\us30\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1430_ ( .A1(\us30\/_0640_ ), .A2(\us30\/_0193_ ), .A3(\us30\/_0091_ ), .B1(\us30\/_0016_ ), .Y(\us30\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1431_ ( .A1(\us30\/_0102_ ), .A2(\us30\/_0301_ ), .B1(\sa30\[3\] ), .C1(\us30\/_0247_ ), .Y(\us30\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1432_ ( .A(\us30\/_0654_ ), .B(\us30\/_0655_ ), .C(\us30\/_0656_ ), .D(\us30\/_0657_ ), .X(\us30\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1433_ ( .A1(\us30\/_0118_ ), .A2(\us30\/_0050_ ), .B1(\us30\/_0038_ ), .C1(\us30\/_0478_ ), .Y(\us30\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us30/_1434_ ( .A_N(\us30\/_0250_ ), .B(\us30\/_0465_ ), .C(\us30\/_0659_ ), .X(\us30\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1435_ ( .A1(\us30\/_0683_ ), .A2(\us30\/_0324_ ), .B1(\us30\/_0255_ ), .Y(\us30\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1436_ ( .A1(\us30\/_0032_ ), .A2(\us30\/_0193_ ), .A3(\us30\/_0047_ ), .B1(\us30\/_0255_ ), .Y(\us30\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1437_ ( .A1(\us30\/_0144_ ), .A2(\us30\/_0586_ ), .A3(\us30\/_0047_ ), .B1(\us30\/_0499_ ), .Y(\us30\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1438_ ( .A(\us30\/_0660_ ), .B(\us30\/_0661_ ), .C(\us30\/_0663_ ), .D(\us30\/_0664_ ), .X(\us30\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1439_ ( .A1(\us30\/_0091_ ), .A2(\us30\/_0276_ ), .B1(\us30\/_0060_ ), .Y(\us30\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1440_ ( .A1(\us30\/_0144_ ), .A2(\us30\/_0608_ ), .B1(\us30\/_0292_ ), .Y(\us30\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1441_ ( .A1(\us30\/_0412_ ), .A2(\us30\/_0038_ ), .B1(\us30\/_0102_ ), .C1(\us30\/_0060_ ), .Y(\us30\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1442_ ( .A1(\sa30\[1\] ), .A2(\us30\/_0734_ ), .B1(\us30\/_0109_ ), .C1(\us30\/_0292_ ), .Y(\us30\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1443_ ( .A(\us30\/_0666_ ), .B(\us30\/_0667_ ), .C(\us30\/_0668_ ), .D(\us30\/_0669_ ), .X(\us30\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1444_ ( .A(\us30\/_0650_ ), .B(\us30\/_0658_ ), .C(\us30\/_0665_ ), .D(\us30\/_0670_ ), .X(\us30\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us30/_1445_ ( .A(\us30\/_0641_ ), .B(\us30\/_0174_ ), .C(\us30\/_0671_ ), .Y(\us30\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us30/_1446_ ( .A(\us30\/_0049_ ), .B(\us30\/_0618_ ), .C_N(\us30\/_0052_ ), .Y(\us30\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us30/_1447_ ( .A(\us30\/_0239_ ), .Y(\us30\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1448_ ( .A(\us30\/_0705_ ), .B(\us30\/_0032_ ), .Y(\us30\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1449_ ( .A1(\us30\/_0054_ ), .A2(\us30\/_0731_ ), .B1(\us30\/_0035_ ), .B2(\us30\/_0705_ ), .Y(\us30\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1450_ ( .A1(\us30\/_0304_ ), .A2(\us30\/_0731_ ), .B1(\us30\/_0047_ ), .B2(\us30\/_0750_ ), .Y(\us30\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1451_ ( .A(\us30\/_0674_ ), .B(\us30\/_0675_ ), .C(\us30\/_0676_ ), .D(\us30\/_0677_ ), .X(\us30\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us30/_1452_ ( .A_N(\us30\/_0584_ ), .B(\us30\/_0283_ ), .X(\us30\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1453_ ( .A(\us30\/_0673_ ), .B(\us30\/_0678_ ), .C(\us30\/_0679_ ), .D(\us30\/_0508_ ), .X(\us30\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1454_ ( .A1(\us30\/_0016_ ), .A2(\us30\/_0733_ ), .B1(\us30\/_0355_ ), .B2(\us30\/_0092_ ), .Y(\us30\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1455_ ( .A(\us30\/_0681_ ), .B(\us30\/_0034_ ), .X(\us30\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us30/_1456_ ( .A1(\us30\/_0330_ ), .A2(\us30\/_0139_ ), .B1(\us30\/_0324_ ), .B2(\us30\/_0089_ ), .X(\us30\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1457_ ( .A1(\us30\/_0146_ ), .A2(\us30\/_0147_ ), .B1(\us30\/_0133_ ), .C1(\us30\/_0684_ ), .Y(\us30\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1458_ ( .A(\us30\/_0113_ ), .B(\us30\/_0251_ ), .Y(\us30\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us30/_1459_ ( .A_N(\us30\/_0463_ ), .B(\us30\/_0686_ ), .C(\us30\/_0383_ ), .D(\us30\/_0464_ ), .X(\us30\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1460_ ( .A1(\us30\/_0051_ ), .A2(\us30\/_0293_ ), .B1(\us30\/_0280_ ), .B2(\us30\/_0705_ ), .Y(\us30\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1461_ ( .A1(\us30\/_0017_ ), .A2(\us30\/_0072_ ), .B1(\us30\/_0134_ ), .B2(\us30\/_0078_ ), .Y(\us30\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1462_ ( .A(\us30\/_0687_ ), .B(\us30\/_0236_ ), .C(\us30\/_0688_ ), .D(\us30\/_0689_ ), .X(\us30\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1463_ ( .A(\us30\/_0680_ ), .B(\us30\/_0682_ ), .C(\us30\/_0685_ ), .D(\us30\/_0690_ ), .X(\us30\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us30/_1464_ ( .A1(\us30\/_0532_ ), .A2(\us30\/_0380_ ), .B1(\us30\/_0102_ ), .C1(\us30\/_0355_ ), .X(\us30\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us30/_1465_ ( .A(\us30\/_0692_ ), .B(\us30\/_0338_ ), .C(\us30\/_0644_ ), .Y(\us30\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1466_ ( .A(\us30\/_0016_ ), .B(\us30\/_0020_ ), .Y(\us30\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1467_ ( .A1(\us30\/_0032_ ), .A2(\us30\/_0137_ ), .B1(\us30\/_0279_ ), .B2(\us30\/_0094_ ), .Y(\us30\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1468_ ( .A1(\us30\/_0575_ ), .A2(\us30\/_0153_ ), .B1(\us30\/_0161_ ), .B2(\us30\/_0293_ ), .Y(\us30\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1469_ ( .A(\us30\/_0259_ ), .B(\us30\/_0695_ ), .C(\us30\/_0696_ ), .D(\us30\/_0697_ ), .X(\us30\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us30/_1470_ ( .A1(\us30\/_0255_ ), .A2(\us30\/_0640_ ), .B1(\us30\/_0016_ ), .B2(\us30\/_0193_ ), .X(\us30\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1471_ ( .A1(\us30\/_0060_ ), .A2(\us30\/_0176_ ), .B1(\us30\/_0699_ ), .C1(\us30\/_0177_ ), .Y(\us30\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1472_ ( .A1(\us30\/_0091_ ), .A2(\us30\/_0499_ ), .B1(\us30\/_0092_ ), .B2(\us30\/_0705_ ), .Y(\us30\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us30/_1473_ ( .A1(\us30\/_0705_ ), .A2(\us30\/_0683_ ), .B1(\us30\/_0093_ ), .B2(\us30\/_0114_ ), .Y(\us30\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us30/_1474_ ( .A1(\us30\/_0683_ ), .A2(\us30\/_0280_ ), .B1(\us30\/_0094_ ), .Y(\us30\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us30/_1475_ ( .A1(\us30\/_0249_ ), .A2(\us30\/_0205_ ), .B1(\us30\/_0038_ ), .C1(\us30\/_0292_ ), .Y(\us30\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1476_ ( .A(\us30\/_0701_ ), .B(\us30\/_0702_ ), .C(\us30\/_0703_ ), .D(\us30\/_0704_ ), .X(\us30\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1477_ ( .A(\us30\/_0693_ ), .B(\us30\/_0698_ ), .C(\us30\/_0700_ ), .D(\us30\/_0706_ ), .X(\us30\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us30/_1478_ ( .A1(\us30\/_0113_ ), .A2(\us30\/_0640_ ), .B1(\us30\/_0099_ ), .B2(\us30\/_0058_ ), .X(\us30\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us30/_1479_ ( .A(\us30\/_0407_ ), .B(\us30\/_0708_ ), .C(\us30\/_0529_ ), .Y(\us30\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1480_ ( .A(\us30\/_0568_ ), .B(\us30\/_0175_ ), .Y(\us30\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us30/_1481_ ( .A1(\us30\/_0247_ ), .A2(\us30\/_0114_ ), .A3(\us30\/_0051_ ), .B1(\us30\/_0130_ ), .Y(\us30\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1482_ ( .A(\us30\/_0709_ ), .B(\us30\/_0550_ ), .C(\us30\/_0710_ ), .D(\us30\/_0711_ ), .X(\us30\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us30/_1483_ ( .A1(\us30\/_0114_ ), .A2(\us30\/_0064_ ), .B1(\us30\/_0261_ ), .B2(\us30\/_0089_ ), .X(\us30\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1484_ ( .A1(\us30\/_0355_ ), .A2(\us30\/_0261_ ), .B1(\us30\/_0198_ ), .C1(\us30\/_0713_ ), .Y(\us30\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1485_ ( .A(\us30\/_0586_ ), .B(\us30\/_0478_ ), .Y(\us30\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us30/_1486_ ( .A_N(\us30\/_0541_ ), .B(\us30\/_0267_ ), .C(\us30\/_0715_ ), .D(\us30\/_0320_ ), .X(\us30\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1487_ ( .A(\us30\/_0586_ ), .B(\us30\/_0070_ ), .Y(\us30\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us30/_1488_ ( .A_N(\us30\/_0211_ ), .B(\us30\/_0155_ ), .C(\us30\/_0202_ ), .D(\us30\/_0718_ ), .X(\us30\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us30/_1489_ ( .A(\us30\/_0150_ ), .B(\us30\/_0205_ ), .C(\us30\/_0380_ ), .Y(\us30\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us30/_1490_ ( .A(\us30\/_0411_ ), .B(\us30\/_0720_ ), .X(\us30\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us30/_1491_ ( .A1(\us30\/_0017_ ), .A2(\us30\/_0022_ ), .B1(\us30\/_0078_ ), .X(\us30\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us30/_1492_ ( .A1(\us30\/_0134_ ), .A2(\us30\/_0738_ ), .B1(\us30\/_0101_ ), .C1(\us30\/_0722_ ), .Y(\us30\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1493_ ( .A(\us30\/_0717_ ), .B(\us30\/_0719_ ), .C(\us30\/_0721_ ), .D(\us30\/_0723_ ), .X(\us30\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us30/_1494_ ( .A(\us30\/_0739_ ), .B(\us30\/_0193_ ), .Y(\us30\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1495_ ( .A(\us30\/_0344_ ), .B(\us30\/_0184_ ), .C(\us30\/_0449_ ), .D(\us30\/_0725_ ), .X(\us30\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us30/_1496_ ( .A(\us30\/_0712_ ), .B(\us30\/_0714_ ), .C(\us30\/_0724_ ), .D(\us30\/_0726_ ), .X(\us30\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \us30/_1497_ ( .A(\us30\/_0691_ ), .B(\us30\/_0707_ ), .C(\us30\/_0728_ ), .Y(\us30\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \us31/_0753_ ( .A(\sa31\[2\] ), .B_N(\sa31\[3\] ), .Y(\us31\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \us31/_0755_ ( .A(\sa31\[1\] ), .B(\sa31\[0\] ), .X(\us31\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us31/_0756_ ( .A(\us31\/_0096_ ), .B(\us31\/_0118_ ), .X(\us31\/_0129_ ) );
sky130_fd_sc_hd__and2_1 \us31/_0757_ ( .A(\sa31\[7\] ), .B(\sa31\[6\] ), .X(\us31\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_0758_ ( .A(\sa31\[4\] ), .B(\sa31\[5\] ), .Y(\us31\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0759_ ( .A(\us31\/_0140_ ), .B(\us31\/_0151_ ), .X(\us31\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0761_ ( .A(\us31\/_0129_ ), .B(\us31\/_0162_ ), .X(\us31\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0762_ ( .A(\us31\/_0096_ ), .X(\us31\/_0194_ ) );
sky130_fd_sc_hd__nor2b_2 \us31/_0763_ ( .A(\sa31\[1\] ), .B_N(\sa31\[0\] ), .Y(\us31\/_0205_ ) );
sky130_fd_sc_hd__and3_1 \us31/_0765_ ( .A(\us31\/_0162_ ), .B(\us31\/_0194_ ), .C(\us31\/_0205_ ), .X(\us31\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us31/_0766_ ( .A(\us31\/_0183_ ), .SLEEP(\us31\/_0227_ ), .X(\us31\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \us31/_0767_ ( .A(\sa31\[0\] ), .B_N(\sa31\[1\] ), .Y(\us31\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_0768_ ( .A(\sa31\[2\] ), .B(\sa31\[3\] ), .Y(\us31\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0769_ ( .A(\us31\/_0249_ ), .B(\us31\/_0260_ ), .X(\us31\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0771_ ( .A(\us31\/_0271_ ), .X(\us31\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0772_ ( .A(\us31\/_0162_ ), .X(\us31\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_0773_ ( .A(\us31\/_0293_ ), .B(\us31\/_0304_ ), .Y(\us31\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us31/_0774_ ( .A(\sa31\[1\] ), .Y(\us31\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us31/_0776_ ( .A(\sa31\[0\] ), .Y(\us31\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0777_ ( .A(\sa31\[2\] ), .B(\sa31\[3\] ), .X(\us31\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0779_ ( .A(\us31\/_0358_ ), .X(\us31\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_0780_ ( .A1(\us31\/_0325_ ), .A2(\us31\/_0347_ ), .B1(\us31\/_0380_ ), .C1(\us31\/_0304_ ), .Y(\us31\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us31/_0781_ ( .A_N(\us31\/_0238_ ), .B(\us31\/_0314_ ), .C(\us31\/_0391_ ), .X(\us31\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us31/_0782_ ( .A(\sa31\[3\] ), .B_N(\sa31\[2\] ), .Y(\us31\/_0412_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0783_ ( .A(\us31\/_0412_ ), .X(\us31\/_0423_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0784_ ( .A(\us31\/_0423_ ), .B(\us31\/_0205_ ), .X(\us31\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \us31/_0787_ ( .A(\sa31\[5\] ), .B_N(\sa31\[4\] ), .Y(\us31\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0788_ ( .A(\us31\/_0467_ ), .B(\us31\/_0140_ ), .X(\us31\/_0478_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_0791_ ( .A(\us31\/_0134_ ), .B(\us31\/_0218_ ), .Y(\us31\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_0792_ ( .A(\us31\/_0478_ ), .B(\us31\/_0271_ ), .Y(\us31\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0793_ ( .A(\us31\/_0194_ ), .X(\us31\/_0532_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0794_ ( .A(\us31\/_0249_ ), .X(\us31\/_0543_ ) );
sky130_fd_sc_hd__and2_1 \us31/_0795_ ( .A(\us31\/_0543_ ), .B(\us31\/_0358_ ), .X(\us31\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0797_ ( .A(\us31\/_0554_ ), .X(\us31\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us31/_0798_ ( .A(\us31\/_0205_ ), .B(\us31\/_0358_ ), .X(\us31\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0800_ ( .A(\us31\/_0586_ ), .X(\us31\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_0801_ ( .A1(\us31\/_0532_ ), .A2(\us31\/_0575_ ), .A3(\us31\/_0608_ ), .B1(\us31\/_0218_ ), .Y(\us31\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us31/_0802_ ( .A(\us31\/_0401_ ), .B(\us31\/_0510_ ), .C(\us31\/_0521_ ), .D(\us31\/_0619_ ), .X(\us31\/_0629_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0803_ ( .A(\us31\/_0358_ ), .B(\sa31\[1\] ), .X(\us31\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0805_ ( .A(\us31\/_0205_ ), .B(\us31\/_0260_ ), .X(\us31\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0807_ ( .A(\us31\/_0662_ ), .X(\us31\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us31/_0808_ ( .A(\sa31\[6\] ), .B_N(\sa31\[7\] ), .Y(\us31\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \us31/_0809_ ( .A(\us31\/_0467_ ), .B(\us31\/_0694_ ), .X(\us31\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0811_ ( .A(\us31\/_0705_ ), .X(\us31\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_0812_ ( .A1(\us31\/_0640_ ), .A2(\us31\/_0293_ ), .A3(\us31\/_0683_ ), .B1(\us31\/_0727_ ), .Y(\us31\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_0813_ ( .A(\sa31\[1\] ), .B(\sa31\[0\] ), .Y(\us31\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0814_ ( .A(\us31\/_0730_ ), .B(\us31\/_0260_ ), .X(\us31\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0816_ ( .A(\us31\/_0731_ ), .X(\us31\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0817_ ( .A(\sa31\[0\] ), .X(\us31\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us31/_0818_ ( .A1(\us31\/_0325_ ), .A2(\us31\/_0734_ ), .B1(\us31\/_0423_ ), .X(\us31\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0819_ ( .A(\us31\/_0694_ ), .B(\us31\/_0151_ ), .X(\us31\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0821_ ( .A(\us31\/_0736_ ), .X(\us31\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0822_ ( .A(\us31\/_0738_ ), .X(\us31\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_0823_ ( .A1(\us31\/_0733_ ), .A2(\us31\/_0735_ ), .A3(\us31\/_0293_ ), .B1(\us31\/_0739_ ), .Y(\us31\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us31/_0824_ ( .A(\us31\/_0730_ ), .B_N(\us31\/_0358_ ), .Y(\us31\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_0825_ ( .A(\us31\/_0741_ ), .B(\us31\/_0739_ ), .Y(\us31\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_0827_ ( .A1(\us31\/_0118_ ), .A2(\us31\/_0205_ ), .B1(\us31\/_0532_ ), .C1(\us31\/_0739_ ), .Y(\us31\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us31/_0828_ ( .A(\us31\/_0729_ ), .B(\us31\/_0740_ ), .C(\us31\/_0742_ ), .D(\us31\/_0744_ ), .X(\us31\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0829_ ( .A(\us31\/_0423_ ), .B(\us31\/_0730_ ), .X(\us31\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0831_ ( .A(\us31\/_0746_ ), .X(\us31\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us31/_0832_ ( .A(\sa31\[4\] ), .B_N(\sa31\[5\] ), .Y(\us31\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0833_ ( .A(\us31\/_0749_ ), .B(\us31\/_0694_ ), .X(\us31\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0835_ ( .A(\us31\/_0750_ ), .X(\us31\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0836_ ( .A(\us31\/_0752_ ), .X(\us31\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0837_ ( .A(\us31\/_0118_ ), .B(\us31\/_0358_ ), .X(\us31\/_0017_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0839_ ( .A(\us31\/_0752_ ), .B(\us31\/_0017_ ), .X(\us31\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0840_ ( .A(\us31\/_0358_ ), .B(\us31\/_0325_ ), .X(\us31\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0842_ ( .A(\us31\/_0096_ ), .B(\us31\/_0205_ ), .X(\us31\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \us31/_0844_ ( .A1(\us31\/_0020_ ), .A2(\us31\/_0022_ ), .B1(\us31\/_0752_ ), .X(\us31\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_0845_ ( .A1(\us31\/_0748_ ), .A2(\us31\/_0016_ ), .B1(\us31\/_0019_ ), .C1(\us31\/_0024_ ), .Y(\us31\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \us31/_0846_ ( .A(\sa31\[4\] ), .B(\sa31\[5\] ), .X(\us31\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0847_ ( .A(\us31\/_0694_ ), .B(\us31\/_0026_ ), .X(\us31\/_0027_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0850_ ( .A(\us31\/_0358_ ), .B(\us31\/_0730_ ), .X(\us31\/_0030_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0852_ ( .A(\us31\/_0030_ ), .X(\us31\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_0853_ ( .A(\us31\/_0247_ ), .B(\us31\/_0032_ ), .Y(\us31\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_0854_ ( .A(\us31\/_0247_ ), .B(\us31\/_0735_ ), .Y(\us31\/_0034_ ) );
sky130_fd_sc_hd__and2_1 \us31/_0855_ ( .A(\us31\/_0118_ ), .B(\us31\/_0260_ ), .X(\us31\/_0035_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0857_ ( .A(\us31\/_0027_ ), .B(\us31\/_0035_ ), .X(\us31\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0858_ ( .A(\us31\/_0260_ ), .X(\us31\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_0859_ ( .A(\us31\/_0038_ ), .B(\us31\/_0347_ ), .Y(\us31\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us31/_0860_ ( .A_N(\us31\/_0039_ ), .B(\us31\/_0027_ ), .X(\us31\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_0861_ ( .A(\us31\/_0037_ ), .B(\us31\/_0040_ ), .Y(\us31\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us31/_0862_ ( .A(\us31\/_0025_ ), .B(\us31\/_0033_ ), .C(\us31\/_0034_ ), .D(\us31\/_0041_ ), .X(\us31\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0863_ ( .A(\us31\/_0749_ ), .B(\us31\/_0140_ ), .X(\us31\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us31/_0865_ ( .A(\sa31\[0\] ), .B(\sa31\[2\] ), .C(\sa31\[3\] ), .X(\us31\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0866_ ( .A(\us31\/_0043_ ), .B(\us31\/_0045_ ), .X(\us31\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0867_ ( .A(\us31\/_0096_ ), .B(\us31\/_0543_ ), .X(\us31\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0869_ ( .A(\us31\/_0047_ ), .B(\us31\/_0043_ ), .X(\us31\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0870_ ( .A(\us31\/_0730_ ), .X(\us31\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0871_ ( .A(\us31\/_0043_ ), .X(\us31\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_0872_ ( .A1(\us31\/_0118_ ), .A2(\us31\/_0050_ ), .B1(\us31\/_0194_ ), .C1(\us31\/_0051_ ), .Y(\us31\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us31/_0873_ ( .A(\us31\/_0046_ ), .B(\us31\/_0049_ ), .C_N(\us31\/_0052_ ), .Y(\us31\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0874_ ( .A(\us31\/_0026_ ), .B(\us31\/_0140_ ), .X(\us31\/_0054_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_0877_ ( .A1(\us31\/_0532_ ), .A2(\us31\/_0575_ ), .B1(\us31\/_0292_ ), .Y(\us31\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0878_ ( .A(\us31\/_0423_ ), .B(\us31\/_0325_ ), .X(\us31\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0880_ ( .A(\us31\/_0051_ ), .X(\us31\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_0881_ ( .A1(\us31\/_0731_ ), .A2(\us31\/_0035_ ), .A3(\us31\/_0058_ ), .B1(\us31\/_0060_ ), .Y(\us31\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0882_ ( .A(\us31\/_0260_ ), .B(\sa31\[1\] ), .X(\us31\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0884_ ( .A(\us31\/_0062_ ), .X(\us31\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_0885_ ( .A1(\us31\/_0064_ ), .A2(\us31\/_0748_ ), .A3(\us31\/_0683_ ), .B1(\us31\/_0292_ ), .Y(\us31\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us31/_0886_ ( .A(\us31\/_0053_ ), .B(\us31\/_0057_ ), .C(\us31\/_0061_ ), .D(\us31\/_0065_ ), .X(\us31\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us31/_0887_ ( .A(\us31\/_0629_ ), .B(\us31\/_0745_ ), .C(\us31\/_0042_ ), .D(\us31\/_0066_ ), .X(\us31\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us31/_0889_ ( .A(\sa31\[7\] ), .B_N(\sa31\[6\] ), .Y(\us31\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0890_ ( .A(\us31\/_0069_ ), .B(\us31\/_0151_ ), .X(\us31\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0892_ ( .A(\us31\/_0070_ ), .X(\us31\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_0893_ ( .A1(\us31\/_0129_ ), .A2(\us31\/_0586_ ), .B1(\us31\/_0072_ ), .Y(\us31\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_0894_ ( .A1(\us31\/_0380_ ), .A2(\us31\/_0347_ ), .B1(\us31\/_0194_ ), .B2(\us31\/_0205_ ), .Y(\us31\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us31/_0895_ ( .A(\us31\/_0074_ ), .B_N(\us31\/_0070_ ), .Y(\us31\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us31/_0896_ ( .A(\us31\/_0073_ ), .SLEEP(\us31\/_0075_ ), .X(\us31\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us31/_0897_ ( .A(\us31\/_0467_ ), .B(\us31\/_0069_ ), .X(\us31\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0898_ ( .A(\us31\/_0077_ ), .X(\us31\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0899_ ( .A(\us31\/_0412_ ), .B(\us31\/_0118_ ), .X(\us31\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0901_ ( .A(\us31\/_0078_ ), .B(\us31\/_0079_ ), .X(\us31\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0902_ ( .A(\us31\/_0412_ ), .B(\us31\/_0249_ ), .X(\us31\/_0082_ ) );
sky130_fd_sc_hd__buf_2 \us31/_0904_ ( .A(\us31\/_0082_ ), .X(\us31\/_0084_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0905_ ( .A(\us31\/_0084_ ), .B(\us31\/_0078_ ), .X(\us31\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us31/_0906_ ( .A1(\sa31\[0\] ), .A2(\us31\/_0325_ ), .B1(\us31\/_0260_ ), .Y(\us31\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us31/_0907_ ( .A_N(\us31\/_0086_ ), .B(\us31\/_0078_ ), .X(\us31\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us31/_0908_ ( .A(\us31\/_0081_ ), .B(\us31\/_0085_ ), .C(\us31\/_0087_ ), .Y(\us31\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0909_ ( .A(\us31\/_0072_ ), .X(\us31\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_0910_ ( .A1(\us31\/_0733_ ), .A2(\us31\/_0748_ ), .A3(\us31\/_0683_ ), .B1(\us31\/_0089_ ), .Y(\us31\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0911_ ( .A(\us31\/_0129_ ), .X(\us31\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0912_ ( .A(\us31\/_0017_ ), .X(\us31\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0913_ ( .A(\us31\/_0022_ ), .X(\us31\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0914_ ( .A(\us31\/_0078_ ), .X(\us31\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_0915_ ( .A1(\us31\/_0091_ ), .A2(\us31\/_0092_ ), .A3(\us31\/_0093_ ), .B1(\us31\/_0094_ ), .Y(\us31\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us31/_0916_ ( .A(\us31\/_0076_ ), .B(\us31\/_0088_ ), .C(\us31\/_0090_ ), .D(\us31\/_0095_ ), .X(\us31\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us31/_0917_ ( .A(\us31\/_0069_ ), .B(\us31\/_0026_ ), .X(\us31\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \us31/_0918_ ( .A(\us31\/_0098_ ), .X(\us31\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0919_ ( .A(\us31\/_0434_ ), .B(\us31\/_0099_ ), .X(\us31\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0920_ ( .A(\us31\/_0079_ ), .B(\us31\/_0098_ ), .X(\us31\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0921_ ( .A(\us31\/_0325_ ), .X(\us31\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_0922_ ( .A1(\us31\/_0102_ ), .A2(\us31\/_0734_ ), .B1(\us31\/_0038_ ), .C1(\us31\/_0099_ ), .Y(\us31\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us31/_0923_ ( .A(\us31\/_0100_ ), .B(\us31\/_0101_ ), .C_N(\us31\/_0103_ ), .Y(\us31\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_0924_ ( .A1(\us31\/_0554_ ), .A2(\us31\/_0586_ ), .B1(\us31\/_0099_ ), .Y(\us31\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_0925_ ( .A(\us31\/_0129_ ), .B(\us31\/_0099_ ), .Y(\us31\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0926_ ( .A(\us31\/_0105_ ), .B(\us31\/_0106_ ), .X(\us31\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0927_ ( .A(\us31\/_0423_ ), .X(\us31\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us31/_0928_ ( .A(\us31\/_0260_ ), .B(\sa31\[0\] ), .X(\us31\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0929_ ( .A(\us31\/_0069_ ), .B(\us31\/_0749_ ), .X(\us31\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0931_ ( .A(\us31\/_0111_ ), .X(\us31\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0932_ ( .A(\us31\/_0113_ ), .X(\us31\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_0933_ ( .A1(\us31\/_0109_ ), .A2(\us31\/_0110_ ), .B1(\us31\/_0114_ ), .Y(\us31\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us31/_0934_ ( .A(\us31\/_0022_ ), .Y(\us31\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us31/_0935_ ( .A(\us31\/_0554_ ), .Y(\us31\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us31/_0936_ ( .A1(\us31\/_0050_ ), .A2(\us31\/_0118_ ), .B1(\us31\/_0194_ ), .Y(\us31\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us31/_0937_ ( .A(\us31\/_0113_ ), .Y(\us31\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us31/_0938_ ( .A1(\us31\/_0116_ ), .A2(\us31\/_0117_ ), .A3(\us31\/_0119_ ), .B1(\us31\/_0120_ ), .X(\us31\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us31/_0939_ ( .A(\us31\/_0104_ ), .B(\us31\/_0108_ ), .C(\us31\/_0115_ ), .D(\us31\/_0121_ ), .X(\us31\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_0940_ ( .A(\sa31\[7\] ), .B(\sa31\[6\] ), .Y(\us31\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0941_ ( .A(\us31\/_0749_ ), .B(\us31\/_0123_ ), .X(\us31\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0943_ ( .A(\us31\/_0082_ ), .B(\us31\/_0124_ ), .X(\us31\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_0944_ ( .A(\us31\/_0271_ ), .B(\us31\/_0124_ ), .Y(\us31\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0945_ ( .A(\us31\/_0124_ ), .X(\us31\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0946_ ( .A(\us31\/_0260_ ), .B(\us31\/_0325_ ), .X(\us31\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_0948_ ( .A(\us31\/_0128_ ), .B(\us31\/_0130_ ), .Y(\us31\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_0949_ ( .A(\us31\/_0127_ ), .B(\us31\/_0132_ ), .Y(\us31\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us31/_0950_ ( .A(\us31\/_0434_ ), .X(\us31\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_0951_ ( .A(\us31\/_0134_ ), .B(\us31\/_0128_ ), .Y(\us31\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us31/_0952_ ( .A(\us31\/_0126_ ), .B(\us31\/_0133_ ), .C_N(\us31\/_0135_ ), .Y(\us31\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us31/_0953_ ( .A(\us31\/_0026_ ), .B(\us31\/_0123_ ), .X(\us31\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0955_ ( .A(\us31\/_0137_ ), .X(\us31\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_0956_ ( .A1(\us31\/_0110_ ), .A2(\us31\/_0293_ ), .A3(\us31\/_0084_ ), .B1(\us31\/_0139_ ), .Y(\us31\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0957_ ( .A(\us31\/_0096_ ), .B(\us31\/_0730_ ), .X(\us31\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0959_ ( .A(\us31\/_0142_ ), .X(\us31\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_0960_ ( .A1(\us31\/_0020_ ), .A2(\us31\/_0144_ ), .A3(\us31\/_0017_ ), .B1(\us31\/_0139_ ), .Y(\us31\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \us31/_0961_ ( .A(\sa31\[2\] ), .B(\us31\/_0050_ ), .C_N(\sa31\[3\] ), .Y(\us31\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0962_ ( .A(\us31\/_0128_ ), .X(\us31\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_0963_ ( .A1(\us31\/_0146_ ), .A2(\us31\/_0032_ ), .A3(\us31\/_0640_ ), .B1(\us31\/_0147_ ), .Y(\us31\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us31/_0964_ ( .A(\us31\/_0136_ ), .B(\us31\/_0141_ ), .C(\us31\/_0145_ ), .D(\us31\/_0148_ ), .X(\us31\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0965_ ( .A(\us31\/_0123_ ), .B(\us31\/_0151_ ), .X(\us31\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0967_ ( .A(\us31\/_0150_ ), .X(\us31\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \us31/_0968_ ( .A(\us31\/_0150_ ), .B(\us31\/_0062_ ), .X(\us31\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_0969_ ( .A(\us31\/_0079_ ), .B(\us31\/_0150_ ), .Y(\us31\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us31/_0970_ ( .A(\us31\/_0150_ ), .B(\us31\/_0423_ ), .C(\us31\/_0543_ ), .Y(\us31\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_0971_ ( .A(\us31\/_0155_ ), .B(\us31\/_0156_ ), .Y(\us31\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_0972_ ( .A1(\us31\/_0153_ ), .A2(\us31\/_0134_ ), .B1(\us31\/_0154_ ), .C1(\us31\/_0157_ ), .Y(\us31\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0973_ ( .A(\us31\/_0467_ ), .B(\us31\/_0123_ ), .X(\us31\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_0975_ ( .A(\us31\/_0159_ ), .X(\us31\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us31/_0976_ ( .A_N(\us31\/_0119_ ), .B(\us31\/_0161_ ), .X(\us31\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us31/_0977_ ( .A(\us31\/_0163_ ), .Y(\us31\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_0978_ ( .A1(\us31\/_0146_ ), .A2(\us31\/_0575_ ), .A3(\us31\/_0608_ ), .B1(\us31\/_0153_ ), .Y(\us31\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_0979_ ( .A1(\us31\/_0062_ ), .A2(\us31\/_0084_ ), .A3(\us31\/_0134_ ), .B1(\us31\/_0161_ ), .Y(\us31\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us31/_0980_ ( .A(\us31\/_0158_ ), .B(\us31\/_0164_ ), .C(\us31\/_0165_ ), .D(\us31\/_0166_ ), .X(\us31\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us31/_0981_ ( .A(\us31\/_0097_ ), .B(\us31\/_0122_ ), .C(\us31\/_0149_ ), .D(\us31\/_0167_ ), .X(\us31\/_0168_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0982_ ( .A(\us31\/_0662_ ), .B(\us31\/_0150_ ), .X(\us31\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_0983_ ( .A(\us31\/_0154_ ), .B(\us31\/_0169_ ), .Y(\us31\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us31/_0984_ ( .A(\us31\/_0123_ ), .B(\us31\/_0151_ ), .C(\us31\/_0038_ ), .X(\us31\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0985_ ( .A(\us31\/_0170_ ), .B(\us31\/_0171_ ), .X(\us31\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \us31/_0986_ ( .A(\us31\/_0172_ ), .Y(\us31\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \us31/_0987_ ( .A(\us31\/_0067_ ), .B(\us31\/_0168_ ), .C(\us31\/_0174_ ), .Y(\us31\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us31/_0988_ ( .A(\sa31\[1\] ), .B(\sa31\[0\] ), .Y(\us31\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us31/_0989_ ( .A(\us31\/_0175_ ), .B(\us31\/_0358_ ), .X(\us31\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0990_ ( .A(\us31\/_0176_ ), .B(\us31\/_0478_ ), .X(\us31\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_0991_ ( .A(\us31\/_0084_ ), .B(\us31\/_0113_ ), .Y(\us31\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0992_ ( .A(\us31\/_0111_ ), .B(\us31\/_0062_ ), .X(\us31\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0993_ ( .A(\us31\/_0111_ ), .B(\us31\/_0662_ ), .X(\us31\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_0994_ ( .A(\us31\/_0179_ ), .B(\us31\/_0180_ ), .Y(\us31\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0995_ ( .A(\us31\/_0054_ ), .B(\us31\/_0058_ ), .X(\us31\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us31/_0996_ ( .A(\us31\/_0182_ ), .Y(\us31\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us31/_0997_ ( .A_N(\us31\/_0177_ ), .B(\us31\/_0178_ ), .C(\us31\/_0181_ ), .D(\us31\/_0184_ ), .X(\us31\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0998_ ( .A(\us31\/_0098_ ), .B(\us31\/_0741_ ), .X(\us31\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us31/_0999_ ( .A(\us31\/_0047_ ), .B(\us31\/_0098_ ), .X(\us31\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us31/_1000_ ( .A(\us31\/_0186_ ), .B(\us31\/_0187_ ), .X(\us31\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1001_ ( .A(\us31\/_0188_ ), .Y(\us31\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1002_ ( .A(\us31\/_0738_ ), .B(\us31\/_0735_ ), .X(\us31\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1003_ ( .A(\us31\/_0271_ ), .B(\us31\/_0736_ ), .X(\us31\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_1004_ ( .A(\us31\/_0190_ ), .B(\us31\/_0191_ ), .Y(\us31\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us31/_1005_ ( .A(\us31\/_0096_ ), .B(\us31\/_0325_ ), .X(\us31\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1006_ ( .A1(\us31\/_0193_ ), .A2(\us31\/_0176_ ), .B1(\us31\/_0043_ ), .Y(\us31\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1007_ ( .A(\us31\/_0185_ ), .B(\us31\/_0189_ ), .C(\us31\/_0192_ ), .D(\us31\/_0195_ ), .X(\us31\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us31/_1008_ ( .A_N(\sa31\[3\] ), .B(\us31\/_0734_ ), .C(\sa31\[2\] ), .X(\us31\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1009_ ( .A(\us31\/_0137_ ), .B(\us31\/_0197_ ), .X(\us31\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_1010_ ( .A(\us31\/_0198_ ), .B(\us31\/_0040_ ), .Y(\us31\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1011_ ( .A(\us31\/_0293_ ), .B(\us31\/_0137_ ), .X(\us31\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1012_ ( .A(\us31\/_0200_ ), .Y(\us31\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1013_ ( .A(\us31\/_0137_ ), .B(\us31\/_0110_ ), .Y(\us31\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1014_ ( .A(\us31\/_0139_ ), .B(\us31\/_0020_ ), .Y(\us31\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1015_ ( .A(\us31\/_0199_ ), .B(\us31\/_0201_ ), .C(\us31\/_0202_ ), .D(\us31\/_0203_ ), .X(\us31\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us31/_1016_ ( .A1(\us31\/_0532_ ), .A2(\us31\/_0109_ ), .B1(\us31\/_0102_ ), .C1(\us31\/_0727_ ), .X(\us31\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1017_ ( .A(\us31\/_0022_ ), .B(\us31\/_0078_ ), .Y(\us31\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1018_ ( .A(\us31\/_0078_ ), .B(\us31\/_0142_ ), .Y(\us31\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1019_ ( .A(\us31\/_0207_ ), .B(\us31\/_0208_ ), .Y(\us31\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1020_ ( .A1(\us31\/_0094_ ), .A2(\us31\/_0176_ ), .B1(\us31\/_0206_ ), .C1(\us31\/_0209_ ), .Y(\us31\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1021_ ( .A(\us31\/_0662_ ), .B(\us31\/_0070_ ), .X(\us31\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us31/_1022_ ( .A(\us31\/_0731_ ), .B(\us31\/_0123_ ), .C(\us31\/_0749_ ), .Y(\us31\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us31/_1023_ ( .A(\us31\/_0731_ ), .B(\us31\/_0467_ ), .C(\us31\/_0069_ ), .Y(\us31\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us31/_1024_ ( .A_N(\us31\/_0211_ ), .B(\us31\/_0127_ ), .C(\us31\/_0212_ ), .D(\us31\/_0213_ ), .X(\us31\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1025_ ( .A(\us31\/_0137_ ), .Y(\us31\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1026_ ( .A(\us31\/_0128_ ), .B(\us31\/_0035_ ), .Y(\us31\/_0217_ ) );
sky130_fd_sc_hd__buf_2 \us31/_1027_ ( .A(\us31\/_0478_ ), .X(\us31\/_0218_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1028_ ( .A1(\us31\/_0159_ ), .A2(\us31\/_0746_ ), .B1(\us31\/_0434_ ), .B2(\us31\/_0218_ ), .Y(\us31\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us31/_1029_ ( .A1(\us31\/_0116_ ), .A2(\us31\/_0215_ ), .B1(\us31\/_0217_ ), .C1(\us31\/_0219_ ), .X(\us31\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1030_ ( .A(\us31\/_0113_ ), .B(\us31\/_0746_ ), .X(\us31\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us31/_1031_ ( .A1(\us31\/_0098_ ), .A2(\us31\/_0746_ ), .B1(\us31\/_0434_ ), .B2(\us31\/_0750_ ), .X(\us31\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1032_ ( .A1(\us31\/_0047_ ), .A2(\us31\/_0113_ ), .B1(\us31\/_0221_ ), .C1(\us31\/_0222_ ), .Y(\us31\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us31/_1033_ ( .A1(\us31\/_0129_ ), .A2(\us31\/_0162_ ), .B1(\us31\/_0271_ ), .B2(\us31\/_0705_ ), .X(\us31\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1034_ ( .A1(\us31\/_0093_ ), .A2(\us31\/_0738_ ), .B1(\us31\/_0081_ ), .C1(\us31\/_0224_ ), .Y(\us31\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1035_ ( .A(\us31\/_0214_ ), .B(\us31\/_0220_ ), .C(\us31\/_0223_ ), .D(\us31\/_0225_ ), .X(\us31\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1036_ ( .A(\us31\/_0196_ ), .B(\us31\/_0204_ ), .C(\us31\/_0210_ ), .D(\us31\/_0226_ ), .X(\us31\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1037_ ( .A(\us31\/_0111_ ), .B(\us31\/_0554_ ), .X(\us31\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1038_ ( .A(\us31\/_0229_ ), .Y(\us31\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1039_ ( .A(\us31\/_0111_ ), .B(\us31\/_0129_ ), .Y(\us31\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1040_ ( .A(\us31\/_0017_ ), .B(\us31\/_0738_ ), .Y(\us31\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1041_ ( .A(\us31\/_0030_ ), .B(\us31\/_0304_ ), .Y(\us31\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1042_ ( .A(\us31\/_0230_ ), .B(\us31\/_0231_ ), .C(\us31\/_0232_ ), .D(\us31\/_0233_ ), .X(\us31\/_0234_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1043_ ( .A(\us31\/_0047_ ), .B(\us31\/_0478_ ), .X(\us31\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1044_ ( .A1(\us31\/_0129_ ), .A2(\us31\/_0554_ ), .B1(\us31\/_0137_ ), .Y(\us31\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us31/_1045_ ( .A(\us31\/_0235_ ), .B(\us31\/_0049_ ), .C_N(\us31\/_0236_ ), .Y(\us31\/_0237_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1046_ ( .A(\us31\/_0047_ ), .B(\us31\/_0077_ ), .X(\us31\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1047_ ( .A(\us31\/_0070_ ), .B(\us31\/_0035_ ), .X(\us31\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us31/_1048_ ( .A1(\us31\/_0047_ ), .A2(\us31\/_0736_ ), .B1(\us31\/_0022_ ), .B2(\us31\/_0099_ ), .X(\us31\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us31/_1049_ ( .A(\us31\/_0239_ ), .B(\us31\/_0240_ ), .C(\us31\/_0241_ ), .Y(\us31\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1050_ ( .A(\us31\/_0554_ ), .B(\us31\/_0072_ ), .X(\us31\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us31/_1051_ ( .A1(\us31\/_0142_ ), .A2(\us31\/_0137_ ), .B1(\us31\/_0159_ ), .B2(\us31\/_0082_ ), .X(\us31\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1052_ ( .A1(\us31\/_0608_ ), .A2(\us31\/_0072_ ), .B1(\us31\/_0243_ ), .C1(\us31\/_0244_ ), .Y(\us31\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1053_ ( .A(\us31\/_0234_ ), .B(\us31\/_0237_ ), .C(\us31\/_0242_ ), .D(\us31\/_0245_ ), .X(\us31\/_0246_ ) );
sky130_fd_sc_hd__buf_2 \us31/_1054_ ( .A(\us31\/_0027_ ), .X(\us31\/_0247_ ) );
sky130_fd_sc_hd__o21a_1 \us31/_1055_ ( .A1(\us31\/_0554_ ), .A2(\us31\/_0586_ ), .B1(\us31\/_0247_ ), .X(\us31\/_0248_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1056_ ( .A(\us31\/_0082_ ), .B(\us31\/_0478_ ), .X(\us31\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_1057_ ( .A(\us31\/_0079_ ), .X(\us31\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1058_ ( .A(\us31\/_0251_ ), .B(\us31\/_0478_ ), .X(\us31\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_1059_ ( .A(\us31\/_0250_ ), .B(\us31\/_0252_ ), .Y(\us31\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1060_ ( .A(\us31\/_0016_ ), .B(\us31\/_0064_ ), .Y(\us31\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_1061_ ( .A(\us31\/_0304_ ), .X(\us31\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1062_ ( .A(\us31\/_0255_ ), .B(\us31\/_0640_ ), .Y(\us31\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us31/_1063_ ( .A_N(\us31\/_0248_ ), .B(\us31\/_0253_ ), .C(\us31\/_0254_ ), .D(\us31\/_0256_ ), .X(\us31\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1064_ ( .A(\us31\/_0099_ ), .B(\us31\/_0110_ ), .X(\us31\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us31/_1065_ ( .A1(\us31\/_0161_ ), .A2(\us31\/_0130_ ), .B1(\us31\/_0258_ ), .Y(\us31\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1066_ ( .A(\us31\/_0194_ ), .B(\sa31\[1\] ), .X(\us31\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1068_ ( .A(\us31\/_0261_ ), .B(\us31\/_0153_ ), .Y(\us31\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us31/_1069_ ( .A_N(\us31\/_0154_ ), .B(\us31\/_0259_ ), .C(\us31\/_0263_ ), .X(\us31\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1070_ ( .A(\us31\/_0246_ ), .B(\us31\/_0174_ ), .C(\us31\/_0257_ ), .D(\us31\/_0264_ ), .X(\us31\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us31/_1071_ ( .A1(\us31\/_0261_ ), .A2(\us31\/_0554_ ), .B1(\us31\/_0159_ ), .X(\us31\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1072_ ( .A(\us31\/_0746_ ), .B(\us31\/_0150_ ), .Y(\us31\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1073_ ( .A(\us31\/_0175_ ), .Y(\us31\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us31/_1074_ ( .A(\us31\/_0423_ ), .B(\us31\/_0123_ ), .C(\us31\/_0151_ ), .X(\us31\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1075_ ( .A(\us31\/_0268_ ), .B(\us31\/_0269_ ), .Y(\us31\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us31/_1076_ ( .A_N(\us31\/_0266_ ), .B(\us31\/_0267_ ), .C(\us31\/_0270_ ), .X(\us31\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1077_ ( .A(\us31\/_0554_ ), .B(\us31\/_0150_ ), .X(\us31\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1078_ ( .A(\us31\/_0273_ ), .Y(\us31\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1079_ ( .A1(\us31\/_0734_ ), .A2(\us31\/_0325_ ), .B1(\us31\/_0380_ ), .Y(\us31\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1080_ ( .A(\us31\/_0275_ ), .Y(\us31\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1081_ ( .A(\us31\/_0276_ ), .B(\us31\/_0153_ ), .Y(\us31\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us31/_1082_ ( .A(\us31\/_0272_ ), .B(\us31\/_0274_ ), .C(\us31\/_0277_ ), .X(\us31\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_1083_ ( .A(\us31\/_0035_ ), .X(\us31\/_0279_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1085_ ( .A1(\us31\/_0218_ ), .A2(\us31\/_0279_ ), .B1(\us31\/_0084_ ), .B2(\us31\/_0060_ ), .Y(\us31\/_0281_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1086_ ( .A1(\us31\/_0251_ ), .A2(\us31\/_0434_ ), .B1(\us31\/_0304_ ), .Y(\us31\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1087_ ( .A(\us31\/_0091_ ), .B(\us31\/_0292_ ), .Y(\us31\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1088_ ( .A1(\us31\/_0118_ ), .A2(\us31\/_0050_ ), .B1(\us31\/_0038_ ), .C1(\us31\/_0255_ ), .Y(\us31\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1089_ ( .A(\us31\/_0281_ ), .B(\us31\/_0283_ ), .C(\us31\/_0284_ ), .D(\us31\/_0285_ ), .X(\us31\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1090_ ( .A(\us31\/_0082_ ), .B(\us31\/_0027_ ), .X(\us31\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1091_ ( .A(\us31\/_0129_ ), .B(\us31\/_0027_ ), .X(\us31\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_1092_ ( .A(\us31\/_0287_ ), .B(\us31\/_0288_ ), .Y(\us31\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1093_ ( .A1(\us31\/_0752_ ), .A2(\us31\/_0683_ ), .B1(\us31\/_0093_ ), .B2(\us31\/_0247_ ), .Y(\us31\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1094_ ( .A1(\us31\/_0092_ ), .A2(\us31\/_0575_ ), .B1(\us31\/_0292_ ), .Y(\us31\/_0291_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_1095_ ( .A(\us31\/_0054_ ), .X(\us31\/_0292_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1096_ ( .A1(\us31\/_0218_ ), .A2(\us31\/_0662_ ), .B1(\us31\/_0084_ ), .B2(\us31\/_0292_ ), .Y(\us31\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1097_ ( .A(\us31\/_0289_ ), .B(\us31\/_0290_ ), .C(\us31\/_0291_ ), .D(\us31\/_0294_ ), .X(\us31\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1098_ ( .A(\us31\/_0750_ ), .B(\us31\/_0193_ ), .X(\us31\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1099_ ( .A(\us31\/_0705_ ), .B(\us31\/_0380_ ), .X(\us31\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1100_ ( .A(\us31\/_0752_ ), .B(\us31\/_0129_ ), .Y(\us31\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us31/_1101_ ( .A(\us31\/_0296_ ), .B(\us31\/_0297_ ), .C_N(\us31\/_0298_ ), .Y(\us31\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1102_ ( .A(\us31\/_0089_ ), .B(\us31\/_0532_ ), .Y(\us31\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1103_ ( .A(\sa31\[2\] ), .Y(\us31\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \us31/_1104_ ( .A(\us31\/_0301_ ), .B(\sa31\[3\] ), .C(\us31\/_0118_ ), .Y(\us31\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1105_ ( .A(\us31\/_0072_ ), .B(\us31\/_0302_ ), .X(\us31\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1106_ ( .A(\us31\/_0303_ ), .Y(\us31\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1107_ ( .A(\us31\/_0147_ ), .B(\us31\/_0302_ ), .Y(\us31\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1108_ ( .A(\us31\/_0299_ ), .B(\us31\/_0300_ ), .C(\us31\/_0305_ ), .D(\us31\/_0306_ ), .X(\us31\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1109_ ( .A(\us31\/_0278_ ), .B(\us31\/_0286_ ), .C(\us31\/_0295_ ), .D(\us31\/_0307_ ), .X(\us31\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us31/_1110_ ( .A(\us31\/_0228_ ), .B(\us31\/_0265_ ), .C(\us31\/_0308_ ), .Y(\us31\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1111_ ( .A(\us31\/_0235_ ), .Y(\us31\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1112_ ( .A(\us31\/_0478_ ), .B(\us31\/_0640_ ), .X(\us31\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1113_ ( .A(\us31\/_0310_ ), .Y(\us31\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1114_ ( .A(\us31\/_0022_ ), .B(\us31\/_0218_ ), .Y(\us31\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1115_ ( .A(\us31\/_0218_ ), .B(\us31\/_0032_ ), .Y(\us31\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1116_ ( .A(\us31\/_0309_ ), .B(\us31\/_0311_ ), .C(\us31\/_0312_ ), .D(\us31\/_0313_ ), .X(\us31\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1117_ ( .A(\us31\/_0218_ ), .B(\us31\/_0064_ ), .Y(\us31\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1118_ ( .A(\us31\/_0218_ ), .B(\us31\/_0683_ ), .Y(\us31\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1119_ ( .A(\us31\/_0315_ ), .B(\us31\/_0316_ ), .C(\us31\/_0317_ ), .D(\us31\/_0253_ ), .X(\us31\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1120_ ( .A(\us31\/_0047_ ), .B(\us31\/_0304_ ), .Y(\us31\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1121_ ( .A(\us31\/_0586_ ), .B(\us31\/_0162_ ), .Y(\us31\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1122_ ( .A(\us31\/_0319_ ), .B(\us31\/_0320_ ), .Y(\us31\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_1123_ ( .A(\us31\/_0321_ ), .B(\us31\/_0238_ ), .Y(\us31\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1124_ ( .A(\us31\/_0304_ ), .B(\us31\/_0062_ ), .Y(\us31\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_1125_ ( .A(\us31\/_0251_ ), .X(\us31\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1126_ ( .A1(\us31\/_0324_ ), .A2(\us31\/_0084_ ), .B1(\us31\/_0255_ ), .Y(\us31\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1127_ ( .A1(\us31\/_0050_ ), .A2(\us31\/_0205_ ), .B1(\us31\/_0109_ ), .C1(\us31\/_0255_ ), .Y(\us31\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1128_ ( .A(\us31\/_0322_ ), .B(\us31\/_0323_ ), .C(\us31\/_0326_ ), .D(\us31\/_0327_ ), .X(\us31\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1129_ ( .A1(\us31\/_0733_ ), .A2(\us31\/_0279_ ), .A3(\us31\/_0058_ ), .B1(\us31\/_0292_ ), .Y(\us31\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_1130_ ( .A(\us31\/_0047_ ), .X(\us31\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1131_ ( .A(\us31\/_0330_ ), .B(\us31\/_0292_ ), .Y(\us31\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1132_ ( .A(\us31\/_0054_ ), .B(\us31\/_0045_ ), .Y(\us31\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1133_ ( .A(\us31\/_0329_ ), .B(\us31\/_0331_ ), .C(\us31\/_0284_ ), .D(\us31\/_0332_ ), .X(\us31\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us31/_1134_ ( .A1(\us31\/_0543_ ), .A2(\us31\/_0205_ ), .B1(\us31\/_0532_ ), .C1(\us31\/_0060_ ), .X(\us31\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1135_ ( .A(\us31\/_0084_ ), .B(\us31\/_0060_ ), .Y(\us31\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1136_ ( .A(\us31\/_0324_ ), .B(\us31\/_0060_ ), .Y(\us31\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1137_ ( .A(\us31\/_0335_ ), .B(\us31\/_0337_ ), .Y(\us31\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1138_ ( .A1(\us31\/_0276_ ), .A2(\us31\/_0060_ ), .B1(\us31\/_0334_ ), .C1(\us31\/_0338_ ), .Y(\us31\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1139_ ( .A(\us31\/_0318_ ), .B(\us31\/_0328_ ), .C(\us31\/_0333_ ), .D(\us31\/_0339_ ), .X(\us31\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us31/_1140_ ( .A1(\us31\/_0746_ ), .A2(\us31\/_0134_ ), .B1(\us31\/_0128_ ), .X(\us31\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us31/_1141_ ( .A_N(\us31\/_0086_ ), .B(\us31\/_0128_ ), .X(\us31\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1142_ ( .A(\us31\/_0079_ ), .B(\us31\/_0124_ ), .X(\us31\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_1143_ ( .A(\us31\/_0126_ ), .B(\us31\/_0343_ ), .Y(\us31\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us31/_1144_ ( .A(\us31\/_0341_ ), .B(\us31\/_0342_ ), .C_N(\us31\/_0344_ ), .Y(\us31\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1146_ ( .A1(\us31\/_0193_ ), .A2(\us31\/_0092_ ), .A3(\us31\/_0330_ ), .B1(\us31\/_0147_ ), .Y(\us31\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1147_ ( .A1(\us31\/_0130_ ), .A2(\us31\/_0084_ ), .A3(\us31\/_0134_ ), .B1(\us31\/_0139_ ), .Y(\us31\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1148_ ( .A1(\us31\/_0144_ ), .A2(\us31\/_0608_ ), .A3(\us31\/_0092_ ), .B1(\us31\/_0139_ ), .Y(\us31\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1149_ ( .A(\us31\/_0345_ ), .B(\us31\/_0348_ ), .C(\us31\/_0349_ ), .D(\us31\/_0350_ ), .X(\us31\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us31/_1150_ ( .A(\us31\/_0150_ ), .B(\us31\/_0194_ ), .C(\us31\/_0543_ ), .X(\us31\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us31/_1151_ ( .A(\us31\/_0277_ ), .SLEEP(\us31\/_0352_ ), .X(\us31\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us31/_1152_ ( .A1(\us31\/_0268_ ), .A2(\us31\/_0171_ ), .B1(\us31\/_0157_ ), .Y(\us31\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us31/_1153_ ( .A(\us31\/_0161_ ), .X(\us31\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1154_ ( .A1(\us31\/_0279_ ), .A2(\us31\/_0084_ ), .B1(\us31\/_0355_ ), .Y(\us31\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1155_ ( .A1(\us31\/_0020_ ), .A2(\us31\/_0193_ ), .A3(\us31\/_0091_ ), .B1(\us31\/_0355_ ), .Y(\us31\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1156_ ( .A(\us31\/_0353_ ), .B(\us31\/_0354_ ), .C(\us31\/_0356_ ), .D(\us31\/_0357_ ), .X(\us31\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1157_ ( .A(\us31\/_0111_ ), .B(\us31\/_0586_ ), .X(\us31\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1158_ ( .A(\us31\/_0360_ ), .Y(\us31\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us31/_1159_ ( .A1(\us31\/_0119_ ), .A2(\us31\/_0120_ ), .B1(\us31\/_0230_ ), .C1(\us31\/_0361_ ), .X(\us31\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1160_ ( .A1(\us31\/_0662_ ), .A2(\us31\/_0251_ ), .A3(\us31\/_0134_ ), .B1(\us31\/_0114_ ), .Y(\us31\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1162_ ( .A1(\us31\/_0035_ ), .A2(\us31\/_0251_ ), .A3(\us31\/_0134_ ), .B1(\us31\/_0099_ ), .Y(\us31\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1163_ ( .A1(\us31\/_0193_ ), .A2(\us31\/_0608_ ), .B1(\us31\/_0099_ ), .Y(\us31\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1164_ ( .A(\us31\/_0362_ ), .B(\us31\/_0363_ ), .C(\us31\/_0365_ ), .D(\us31\/_0366_ ), .X(\us31\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1165_ ( .A1(\us31\/_0575_ ), .A2(\us31\/_0092_ ), .A3(\us31\/_0330_ ), .B1(\us31\/_0089_ ), .Y(\us31\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1166_ ( .A1(\us31\/_0586_ ), .A2(\us31\/_0017_ ), .A3(\us31\/_0330_ ), .B1(\us31\/_0094_ ), .Y(\us31\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \us31/_1167_ ( .A1(\us31\/_0293_ ), .A2(\us31\/_0134_ ), .B1(\us31\/_0089_ ), .Y(\us31\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1168_ ( .A1(\us31\/_0279_ ), .A2(\us31\/_0134_ ), .B1(\us31\/_0094_ ), .Y(\us31\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1169_ ( .A(\us31\/_0368_ ), .B(\us31\/_0370_ ), .C(\us31\/_0371_ ), .D(\us31\/_0372_ ), .X(\us31\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1170_ ( .A(\us31\/_0351_ ), .B(\us31\/_0359_ ), .C(\us31\/_0367_ ), .D(\us31\/_0373_ ), .X(\us31\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1171_ ( .A1(\us31\/_0102_ ), .A2(\us31\/_0347_ ), .B1(\us31\/_0109_ ), .C1(\us31\/_0247_ ), .Y(\us31\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1172_ ( .A1(\us31\/_0102_ ), .A2(\us31\/_0347_ ), .B1(\us31\/_0532_ ), .C1(\us31\/_0247_ ), .Y(\us31\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1173_ ( .A1(\us31\/_0050_ ), .A2(\us31\/_0543_ ), .B1(\us31\/_0380_ ), .C1(\us31\/_0247_ ), .Y(\us31\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1174_ ( .A(\us31\/_0041_ ), .B(\us31\/_0375_ ), .C(\us31\/_0376_ ), .D(\us31\/_0377_ ), .X(\us31\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1175_ ( .A(\us31\/_0047_ ), .B(\us31\/_0750_ ), .X(\us31\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1176_ ( .A(\us31\/_0379_ ), .Y(\us31\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1177_ ( .A(\us31\/_0016_ ), .B(\us31\/_0608_ ), .Y(\us31\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1178_ ( .A(\us31\/_0752_ ), .B(\us31\/_0554_ ), .Y(\us31\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1179_ ( .A1(\sa31\[1\] ), .A2(\us31\/_0734_ ), .B1(\us31\/_0109_ ), .C1(\us31\/_0016_ ), .Y(\us31\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1180_ ( .A(\us31\/_0381_ ), .B(\us31\/_0382_ ), .C(\us31\/_0383_ ), .D(\us31\/_0384_ ), .X(\us31\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us31/_1181_ ( .A(\us31\/_0086_ ), .B_N(\us31\/_0736_ ), .X(\us31\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1182_ ( .A1(\us31\/_0748_ ), .A2(\us31\/_0134_ ), .B1(\us31\/_0739_ ), .Y(\us31\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1183_ ( .A1(\us31\/_0118_ ), .A2(\us31\/_0543_ ), .B1(\us31\/_0109_ ), .C1(\us31\/_0739_ ), .Y(\us31\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1184_ ( .A1(\us31\/_0102_ ), .A2(\us31\/_0301_ ), .B1(\sa31\[3\] ), .C1(\us31\/_0739_ ), .Y(\us31\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1185_ ( .A(\us31\/_0386_ ), .B(\us31\/_0387_ ), .C(\us31\/_0388_ ), .D(\us31\/_0389_ ), .X(\us31\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1186_ ( .A(\us31\/_0020_ ), .Y(\us31\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1187_ ( .A(\us31\/_0727_ ), .Y(\us31\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1188_ ( .A(\us31\/_0727_ ), .B(\us31\/_0064_ ), .Y(\us31\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1189_ ( .A1(\us31\/_0102_ ), .A2(\us31\/_0734_ ), .B1(\us31\/_0532_ ), .C1(\us31\/_0727_ ), .Y(\us31\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us31/_1190_ ( .A1(\us31\/_0392_ ), .A2(\us31\/_0393_ ), .B1(\us31\/_0394_ ), .C1(\us31\/_0395_ ), .X(\us31\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1191_ ( .A(\us31\/_0378_ ), .B(\us31\/_0385_ ), .C(\us31\/_0390_ ), .D(\us31\/_0396_ ), .X(\us31\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us31/_1192_ ( .A(\us31\/_0340_ ), .B(\us31\/_0374_ ), .C(\us31\/_0397_ ), .Y(\us31\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1193_ ( .A(\us31\/_0077_ ), .B(\us31\/_0129_ ), .X(\us31\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_1194_ ( .A(\us31\/_0398_ ), .B(\us31\/_0239_ ), .Y(\us31\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1195_ ( .A(\us31\/_0022_ ), .B(\us31\/_0111_ ), .X(\us31\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us31/_1196_ ( .A_N(\us31\/_0400_ ), .B(\us31\/_0231_ ), .Y(\us31\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us31/_1197_ ( .A(\us31\/_0399_ ), .SLEEP(\us31\/_0402_ ), .X(\us31\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_1198_ ( .A(\us31\/_0746_ ), .B(\us31\/_0251_ ), .Y(\us31\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us31/_1199_ ( .A_N(\us31\/_0404_ ), .B(\us31\/_0752_ ), .Y(\us31\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us31/_1200_ ( .A(\us31\/_0467_ ), .B(\us31\/_0194_ ), .C(\us31\/_0694_ ), .X(\us31\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us31/_1201_ ( .A_N(\us31\/_0175_ ), .B(\us31\/_0406_ ), .X(\us31\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1202_ ( .A(\us31\/_0407_ ), .Y(\us31\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1203_ ( .A1(\us31\/_0094_ ), .A2(\us31\/_0197_ ), .B1(\us31\/_0114_ ), .B2(\us31\/_0640_ ), .Y(\us31\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1204_ ( .A(\us31\/_0403_ ), .B(\us31\/_0405_ ), .C(\us31\/_0408_ ), .D(\us31\/_0409_ ), .X(\us31\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1205_ ( .A(\us31\/_0030_ ), .B(\us31\/_0150_ ), .Y(\us31\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us31/_1206_ ( .A_N(\us31\/_0169_ ), .B(\us31\/_0289_ ), .C(\us31\/_0411_ ), .X(\us31\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us31/_1207_ ( .A1(\us31\/_0467_ ), .A2(\us31\/_0151_ ), .B1(\us31\/_0140_ ), .C1(\us31\/_0129_ ), .X(\us31\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1208_ ( .A1(\us31\/_0608_ ), .A2(\us31\/_0099_ ), .B1(\us31\/_0037_ ), .C1(\us31\/_0414_ ), .Y(\us31\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1209_ ( .A(\us31\/_0738_ ), .Y(\us31\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1210_ ( .A(\us31\/_0586_ ), .B(\us31\/_0736_ ), .Y(\us31\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1211_ ( .A1(\us31\/_0194_ ), .A2(\us31\/_0038_ ), .B1(\us31\/_0118_ ), .C1(\us31\/_0153_ ), .Y(\us31\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us31/_1212_ ( .A1(\us31\/_0416_ ), .A2(\us31\/_0117_ ), .B1(\us31\/_0417_ ), .C1(\us31\/_0418_ ), .X(\us31\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1213_ ( .A(\us31\/_0077_ ), .B(\us31\/_0035_ ), .X(\us31\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1214_ ( .A(\us31\/_0662_ ), .B(\us31\/_0124_ ), .Y(\us31\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1215_ ( .A(\us31\/_0030_ ), .B(\us31\/_0137_ ), .Y(\us31\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1216_ ( .A(\us31\/_0072_ ), .B(\us31\/_0731_ ), .Y(\us31\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us31/_1217_ ( .A_N(\us31\/_0420_ ), .B(\us31\/_0421_ ), .C(\us31\/_0422_ ), .D(\us31\/_0424_ ), .X(\us31\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1218_ ( .A(\us31\/_0413_ ), .B(\us31\/_0415_ ), .C(\us31\/_0419_ ), .D(\us31\/_0425_ ), .X(\us31\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us31/_1219_ ( .A(\us31\/_0355_ ), .B(\us31\/_0102_ ), .C(\us31\/_0109_ ), .Y(\us31\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1220_ ( .A(\us31\/_0077_ ), .B(\us31\/_0017_ ), .X(\us31\/_0428_ ) );
sky130_fd_sc_hd__and2_1 \us31/_1221_ ( .A(\us31\/_0077_ ), .B(\us31\/_0554_ ), .X(\us31\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us31/_1222_ ( .A1(\us31\/_0050_ ), .A2(\us31\/_0205_ ), .B1(\us31\/_0380_ ), .C1(\us31\/_0078_ ), .X(\us31\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us31/_1223_ ( .A(\us31\/_0428_ ), .B(\us31\/_0429_ ), .C(\us31\/_0430_ ), .Y(\us31\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us31/_1224_ ( .A_N(\us31\/_0209_ ), .B(\us31\/_0431_ ), .X(\us31\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us31/_1225_ ( .A1(\us31\/_0215_ ), .A2(\us31\/_0404_ ), .B1(\us31\/_0427_ ), .C1(\us31\/_0432_ ), .X(\us31\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1226_ ( .A(\us31\/_0043_ ), .B(\us31\/_0058_ ), .Y(\us31\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1227_ ( .A(\us31\/_0195_ ), .B(\us31\/_0233_ ), .C(\us31\/_0320_ ), .D(\us31\/_0435_ ), .X(\us31\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1228_ ( .A(\us31\/_0261_ ), .B(\us31\/_0738_ ), .Y(\us31\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1229_ ( .A1(\us31\/_0218_ ), .A2(\us31\/_0640_ ), .B1(\us31\/_0261_ ), .B2(\us31\/_0292_ ), .Y(\us31\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1230_ ( .A(\us31\/_0436_ ), .B(\us31\/_0394_ ), .C(\us31\/_0437_ ), .D(\us31\/_0438_ ), .X(\us31\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1231_ ( .A(\us31\/_0410_ ), .B(\us31\/_0426_ ), .C(\us31\/_0433_ ), .D(\us31\/_0439_ ), .X(\us31\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us31/_1232_ ( .A(\us31\/_0135_ ), .SLEEP(\us31\/_0273_ ), .X(\us31\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1233_ ( .A1(\us31\/_0279_ ), .A2(\us31\/_0134_ ), .B1(\us31\/_0099_ ), .Y(\us31\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1234_ ( .A(\us31\/_0441_ ), .B(\us31\/_0164_ ), .C(\us31\/_0270_ ), .D(\us31\/_0442_ ), .X(\us31\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1235_ ( .A(\us31\/_0051_ ), .B(\us31\/_0662_ ), .Y(\us31\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1236_ ( .A(\us31\/_0051_ ), .B(\us31\/_0271_ ), .Y(\us31\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1237_ ( .A(\us31\/_0444_ ), .B(\us31\/_0446_ ), .X(\us31\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1238_ ( .A(\us31\/_0193_ ), .B(\us31\/_0304_ ), .X(\us31\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1239_ ( .A(\us31\/_0448_ ), .Y(\us31\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1240_ ( .A(\us31\/_0162_ ), .B(\us31\/_0130_ ), .X(\us31\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1241_ ( .A(\us31\/_0450_ ), .Y(\us31\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1242_ ( .A1(\us31\/_0129_ ), .A2(\us31\/_0554_ ), .B1(\us31\/_0043_ ), .Y(\us31\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1243_ ( .A(\us31\/_0447_ ), .B(\us31\/_0449_ ), .C(\us31\/_0451_ ), .D(\us31\/_0452_ ), .X(\us31\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1244_ ( .A(\us31\/_0292_ ), .B(\us31\/_0064_ ), .Y(\us31\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us31/_1245_ ( .A_N(\us31\/_0248_ ), .B(\us31\/_0454_ ), .C(\us31\/_0254_ ), .D(\us31\/_0256_ ), .X(\us31\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1246_ ( .A1(\us31\/_0330_ ), .A2(\us31\/_0099_ ), .B1(\us31\/_0134_ ), .B2(\us31\/_0705_ ), .Y(\us31\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1247_ ( .A1(\us31\/_0748_ ), .A2(\us31\/_0738_ ), .B1(\us31\/_0092_ ), .B2(\us31\/_0752_ ), .Y(\us31\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1248_ ( .A1(\us31\/_0072_ ), .A2(\us31\/_0035_ ), .B1(\us31\/_0748_ ), .B2(\us31\/_0292_ ), .Y(\us31\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1249_ ( .A1(\us31\/_0748_ ), .A2(\us31\/_0251_ ), .B1(\us31\/_0247_ ), .Y(\us31\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1250_ ( .A(\us31\/_0457_ ), .B(\us31\/_0458_ ), .C(\us31\/_0459_ ), .D(\us31\/_0460_ ), .X(\us31\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1251_ ( .A(\us31\/_0443_ ), .B(\us31\/_0453_ ), .C(\us31\/_0455_ ), .D(\us31\/_0461_ ), .X(\us31\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1252_ ( .A(\us31\/_0705_ ), .B(\us31\/_0079_ ), .X(\us31\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1253_ ( .A(\us31\/_0586_ ), .B(\us31\/_0124_ ), .Y(\us31\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1254_ ( .A(\us31\/_0218_ ), .B(\us31\/_0746_ ), .Y(\us31\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us31/_1255_ ( .A_N(\us31\/_0463_ ), .B(\us31\/_0464_ ), .C(\us31\/_0465_ ), .X(\us31\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us31/_1256_ ( .A1(\us31\/_0271_ ), .A2(\us31\/_0072_ ), .B1(\us31\/_0142_ ), .B2(\us31\/_0027_ ), .X(\us31\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1257_ ( .A1(\us31\/_0144_ ), .A2(\us31\/_0099_ ), .B1(\us31\/_0360_ ), .C1(\us31\/_0468_ ), .Y(\us31\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us31/_1258_ ( .A1(\us31\/_0662_ ), .A2(\us31\/_0251_ ), .B1(\us31\/_0218_ ), .X(\us31\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1259_ ( .A1(\us31\/_0575_ ), .A2(\us31\/_0292_ ), .B1(\us31\/_0379_ ), .C1(\us31\/_0470_ ), .Y(\us31\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1260_ ( .A(\us31\/_0466_ ), .B(\us31\/_0469_ ), .C(\us31\/_0471_ ), .D(\us31\/_0305_ ), .X(\us31\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us31/_1261_ ( .A1(\us31\/_0247_ ), .A2(\us31\/_0683_ ), .B1(\us31\/_0324_ ), .B2(\us31\/_0292_ ), .X(\us31\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1262_ ( .A(\us31\/_0084_ ), .B(\us31\/_0099_ ), .X(\us31\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us31/_1263_ ( .A1(\us31\/_0092_ ), .A2(\us31\/_0247_ ), .B1(\us31\/_0474_ ), .X(\us31\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us31/_1264_ ( .A(\us31\/_0075_ ), .B(\us31\/_0473_ ), .C(\us31\/_0475_ ), .Y(\us31\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1265_ ( .A1(\us31\/_0279_ ), .A2(\us31\/_0255_ ), .B1(\us31\/_0084_ ), .B2(\us31\/_0060_ ), .Y(\us31\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1266_ ( .A1(\us31\/_0093_ ), .A2(\us31\/_0292_ ), .B1(\us31\/_0134_ ), .B2(\us31\/_0114_ ), .Y(\us31\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1267_ ( .A1(\us31\/_0161_ ), .A2(\us31\/_0032_ ), .B1(\us31\/_0324_ ), .B2(\us31\/_0147_ ), .Y(\us31\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1268_ ( .A1(\us31\/_0054_ ), .A2(\us31\/_0731_ ), .B1(\us31\/_0748_ ), .B2(\us31\/_0304_ ), .Y(\us31\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1269_ ( .A(\us31\/_0477_ ), .B(\us31\/_0479_ ), .C(\us31\/_0480_ ), .D(\us31\/_0481_ ), .X(\us31\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1270_ ( .A(\us31\/_0161_ ), .B(\us31\/_0064_ ), .Y(\us31\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us31/_1271_ ( .A(\us31\/_0731_ ), .B(\us31\/_0123_ ), .C(\us31\/_0467_ ), .Y(\us31\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1272_ ( .A(\us31\/_0483_ ), .B(\us31\/_0484_ ), .Y(\us31\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1273_ ( .A(\us31\/_0297_ ), .Y(\us31\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us31/_1274_ ( .A_N(\us31\/_0485_ ), .B(\us31\/_0181_ ), .C(\us31\/_0486_ ), .D(\us31\/_0386_ ), .X(\us31\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1275_ ( .A(\us31\/_0472_ ), .B(\us31\/_0476_ ), .C(\us31\/_0482_ ), .D(\us31\/_0487_ ), .X(\us31\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \us31/_1276_ ( .A(\us31\/_0440_ ), .B(\us31\/_0462_ ), .C(\us31\/_0488_ ), .Y(\us31\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1277_ ( .A(\us31\/_0403_ ), .B(\us31\/_0230_ ), .C(\us31\/_0451_ ), .D(\us31\/_0361_ ), .X(\us31\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1278_ ( .A1(\us31\/_0118_ ), .A2(\us31\/_0050_ ), .B1(\us31\/_0109_ ), .C1(\us31\/_0139_ ), .Y(\us31\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1279_ ( .A(\us31\/_0447_ ), .B(\us31\/_0437_ ), .C(\us31\/_0491_ ), .D(\us31\/_0427_ ), .X(\us31\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1280_ ( .A1(\us31\/_0084_ ), .A2(\us31\/_0255_ ), .B1(\us31\/_0608_ ), .B2(\us31\/_0247_ ), .Y(\us31\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1281_ ( .A1(\us31\/_0144_ ), .A2(\us31\/_0147_ ), .B1(\us31\/_0355_ ), .B2(\us31\/_0093_ ), .Y(\us31\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1282_ ( .A1(\us31\/_0705_ ), .A2(\us31\/_0279_ ), .B1(\us31\/_0330_ ), .B2(\us31\/_0247_ ), .Y(\us31\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1283_ ( .A1(\us31\/_0279_ ), .A2(\us31\/_0084_ ), .B1(\us31\/_0114_ ), .Y(\us31\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1284_ ( .A(\us31\/_0493_ ), .B(\us31\/_0494_ ), .C(\us31\/_0495_ ), .D(\us31\/_0496_ ), .X(\us31\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1285_ ( .A1(\us31\/_0134_ ), .A2(\us31\/_0137_ ), .B1(\us31\/_0355_ ), .B2(\us31\/_0575_ ), .Y(\us31\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1286_ ( .A1(\us31\/_0099_ ), .A2(\us31\/_0733_ ), .B1(\us31\/_0093_ ), .B2(\us31\/_0218_ ), .Y(\us31\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1287_ ( .A(\us31\/_0147_ ), .B(\us31\/_0640_ ), .Y(\us31\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1288_ ( .A1(\us31\/_0153_ ), .A2(\us31\/_0292_ ), .B1(\us31\/_0748_ ), .Y(\us31\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1289_ ( .A(\us31\/_0498_ ), .B(\us31\/_0500_ ), .C(\us31\/_0501_ ), .D(\us31\/_0502_ ), .X(\us31\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1290_ ( .A(\us31\/_0490_ ), .B(\us31\/_0492_ ), .C(\us31\/_0497_ ), .D(\us31\/_0503_ ), .X(\us31\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us31/_1291_ ( .A_N(\us31\/_0275_ ), .B(\us31\/_0705_ ), .X(\us31\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1292_ ( .A(\us31\/_0505_ ), .Y(\us31\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1293_ ( .A(\us31\/_0380_ ), .B(\us31\/_0347_ ), .X(\us31\/_0507_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1294_ ( .A1(\us31\/_0507_ ), .A2(\us31\/_0093_ ), .B1(\us31\/_0292_ ), .Y(\us31\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1295_ ( .A(\us31\/_0322_ ), .B(\us31\/_0277_ ), .C(\us31\/_0506_ ), .D(\us31\/_0508_ ), .X(\us31\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1296_ ( .A(\us31\/_0084_ ), .B(\us31\/_0705_ ), .X(\us31\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1297_ ( .A1(\us31\/_0733_ ), .A2(\us31\/_0114_ ), .B1(\us31\/_0429_ ), .C1(\us31\/_0511_ ), .Y(\us31\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_1298_ ( .A(\us31\/_0019_ ), .B(\us31\/_0024_ ), .Y(\us31\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1299_ ( .A(\us31\/_0512_ ), .B(\us31\/_0513_ ), .C(\us31\/_0742_ ), .D(\us31\/_0306_ ), .X(\us31\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1300_ ( .A1(\us31\/_0532_ ), .A2(\us31\/_0089_ ), .B1(\us31\/_0154_ ), .C1(\us31\/_0169_ ), .Y(\us31\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us31/_1301_ ( .A1(\us31\/_0749_ ), .A2(\us31\/_0026_ ), .B1(\us31\/_0069_ ), .C1(\us31\/_0032_ ), .X(\us31\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us31/_1302_ ( .A1(\us31\/_0324_ ), .A2(\us31\/_0355_ ), .B1(\us31\/_0330_ ), .B2(\us31\/_0727_ ), .X(\us31\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us31/_1303_ ( .A(\us31\/_0133_ ), .B(\us31\/_0516_ ), .C(\us31\/_0517_ ), .Y(\us31\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1304_ ( .A(\us31\/_0509_ ), .B(\us31\/_0514_ ), .C(\us31\/_0515_ ), .D(\us31\/_0518_ ), .X(\us31\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1305_ ( .A(\us31\/_0746_ ), .B(\us31\/_0072_ ), .Y(\us31\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1306_ ( .A1(\us31\/_0082_ ), .A2(\us31\/_0070_ ), .B1(\us31\/_0043_ ), .B2(\us31\/_0193_ ), .Y(\us31\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1307_ ( .A(\us31\/_0311_ ), .B(\us31\/_0520_ ), .C(\us31\/_0332_ ), .D(\us31\/_0522_ ), .X(\us31\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1308_ ( .A(\us31\/_0129_ ), .B(\us31\/_0218_ ), .X(\us31\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_1309_ ( .A(\us31\/_0235_ ), .B(\us31\/_0524_ ), .Y(\us31\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us31/_1310_ ( .A(\us31\/_0081_ ), .B(\us31\/_0085_ ), .Y(\us31\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1311_ ( .A1(\us31\/_0051_ ), .A2(\us31\/_0045_ ), .B1(\us31\/_0130_ ), .B2(\us31\/_0094_ ), .Y(\us31\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1312_ ( .A(\us31\/_0523_ ), .B(\us31\/_0525_ ), .C(\us31\/_0526_ ), .D(\us31\/_0527_ ), .X(\us31\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us31/_1313_ ( .A_N(\us31\/_0250_ ), .B(\us31\/_0521_ ), .Y(\us31\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1314_ ( .A(\us31\/_0128_ ), .B(\us31\/_0020_ ), .X(\us31\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1315_ ( .A(\us31\/_0530_ ), .Y(\us31\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1316_ ( .A(\us31\/_0099_ ), .B(\us31\/_0058_ ), .X(\us31\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1317_ ( .A(\us31\/_0533_ ), .Y(\us31\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us31/_1318_ ( .A_N(\us31\/_0529_ ), .B(\us31\/_0531_ ), .C(\us31\/_0534_ ), .D(\us31\/_0192_ ), .X(\us31\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1319_ ( .A(\us31\/_0434_ ), .B(\us31\/_0078_ ), .X(\us31\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us31/_1320_ ( .A1(\us31\/_0750_ ), .A2(\us31\/_0079_ ), .B1(\us31\/_0129_ ), .B2(\us31\/_0705_ ), .X(\us31\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1321_ ( .A1(\us31\/_0161_ ), .A2(\us31\/_0032_ ), .B1(\us31\/_0536_ ), .C1(\us31\/_0537_ ), .Y(\us31\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us31/_1322_ ( .A1(\us31\/_0746_ ), .A2(\us31\/_0162_ ), .B1(\us31\/_0079_ ), .B2(\us31\/_0043_ ), .X(\us31\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1323_ ( .A1(\us31\/_0093_ ), .A2(\us31\/_0247_ ), .B1(\us31\/_0240_ ), .C1(\us31\/_0539_ ), .Y(\us31\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1324_ ( .A(\us31\/_0434_ ), .B(\us31\/_0043_ ), .X(\us31\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us31/_1325_ ( .A1(\us31\/_0142_ ), .A2(\us31\/_0150_ ), .B1(\us31\/_0022_ ), .B2(\us31\/_0137_ ), .X(\us31\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1326_ ( .A1(\us31\/_0279_ ), .A2(\us31\/_0051_ ), .B1(\us31\/_0541_ ), .C1(\us31\/_0542_ ), .Y(\us31\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1327_ ( .A(\us31\/_0159_ ), .B(\us31\/_0035_ ), .X(\us31\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us31/_1328_ ( .A1(\us31\/_0271_ ), .A2(\us31\/_0434_ ), .B1(\us31\/_0027_ ), .X(\us31\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1329_ ( .A1(\us31\/_0091_ ), .A2(\us31\/_0128_ ), .B1(\us31\/_0545_ ), .C1(\us31\/_0546_ ), .Y(\us31\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1330_ ( .A(\us31\/_0538_ ), .B(\us31\/_0540_ ), .C(\us31\/_0544_ ), .D(\us31\/_0547_ ), .X(\us31\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1331_ ( .A(\us31\/_0099_ ), .B(\us31\/_0193_ ), .X(\us31\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us31/_1332_ ( .A(\us31\/_0549_ ), .B(\us31\/_0186_ ), .C(\us31\/_0187_ ), .Y(\us31\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1333_ ( .A(\us31\/_0062_ ), .B(\us31\/_0347_ ), .C(\us31\/_0749_ ), .D(\us31\/_0694_ ), .X(\us31\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1334_ ( .A1(\us31\/_0130_ ), .A2(\us31\/_0218_ ), .B1(\us31\/_0551_ ), .C1(\us31\/_0101_ ), .Y(\us31\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1335_ ( .A(\us31\/_0139_ ), .B(\us31\/_0640_ ), .Y(\us31\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1336_ ( .A1(\us31\/_0752_ ), .A2(\us31\/_0662_ ), .B1(\us31\/_0084_ ), .B2(\us31\/_0099_ ), .Y(\us31\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1337_ ( .A(\us31\/_0550_ ), .B(\us31\/_0552_ ), .C(\us31\/_0553_ ), .D(\us31\/_0555_ ), .X(\us31\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1338_ ( .A(\us31\/_0528_ ), .B(\us31\/_0535_ ), .C(\us31\/_0548_ ), .D(\us31\/_0556_ ), .X(\us31\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us31/_1339_ ( .A(\us31\/_0504_ ), .B(\us31\/_0519_ ), .C(\us31\/_0557_ ), .Y(\us31\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1340_ ( .A(\us31\/_0054_ ), .B(\us31\/_0507_ ), .X(\us31\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us31/_1341_ ( .A_N(\us31\/_0558_ ), .B(\us31\/_0408_ ), .C(\us31\/_0451_ ), .D(\us31\/_0452_ ), .X(\us31\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1342_ ( .A(\us31\/_0549_ ), .Y(\us31\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1343_ ( .A(\us31\/_0559_ ), .B(\us31\/_0403_ ), .C(\us31\/_0560_ ), .D(\us31\/_0371_ ), .X(\us31\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1344_ ( .A(\us31\/_0181_ ), .B(\us31\/_0178_ ), .X(\us31\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1345_ ( .A(\us31\/_0562_ ), .B(\us31\/_0552_ ), .C(\us31\/_0553_ ), .D(\us31\/_0555_ ), .X(\us31\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1346_ ( .A(\us31\/_0247_ ), .B(\us31\/_0020_ ), .Y(\us31\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1347_ ( .A(\us31\/_0051_ ), .B(\us31\/_0130_ ), .X(\us31\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1348_ ( .A(\us31\/_0566_ ), .Y(\us31\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1349_ ( .A(\us31\/_0159_ ), .B(\us31\/_0423_ ), .X(\us31\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1350_ ( .A1(\us31\/_0752_ ), .A2(\us31\/_0640_ ), .B1(\us31\/_0568_ ), .B2(\us31\/_0175_ ), .Y(\us31\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1351_ ( .A(\us31\/_0076_ ), .B(\us31\/_0565_ ), .C(\us31\/_0567_ ), .D(\us31\/_0569_ ), .X(\us31\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us31/_1352_ ( .A1(\us31\/_0035_ ), .A2(\us31\/_0142_ ), .B1(\us31\/_0161_ ), .X(\us31\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1353_ ( .A(\us31\/_0099_ ), .B(\us31\/_0662_ ), .Y(\us31\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us31/_1354_ ( .A(\us31\/_0420_ ), .B(\us31\/_0571_ ), .C_N(\us31\/_0572_ ), .Y(\us31\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1355_ ( .A(\us31\/_0051_ ), .B(\us31\/_0746_ ), .Y(\us31\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1356_ ( .A(\us31\/_0574_ ), .B(\us31\/_0319_ ), .C(\us31\/_0320_ ), .D(\us31\/_0411_ ), .X(\us31\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1357_ ( .A(\us31\/_0736_ ), .B(\us31\/_0035_ ), .Y(\us31\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1358_ ( .A(\us31\/_0736_ ), .B(\us31\/_0030_ ), .Y(\us31\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1359_ ( .A(\us31\/_0298_ ), .B(\us31\/_0208_ ), .C(\us31\/_0577_ ), .D(\us31\/_0578_ ), .X(\us31\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1360_ ( .A1(\us31\/_0020_ ), .A2(\us31\/_0137_ ), .B1(\us31\/_0261_ ), .B2(\us31\/_0128_ ), .Y(\us31\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1361_ ( .A(\us31\/_0573_ ), .B(\us31\/_0576_ ), .C(\us31\/_0579_ ), .D(\us31\/_0580_ ), .X(\us31\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1362_ ( .A(\us31\/_0561_ ), .B(\us31\/_0563_ ), .C(\us31\/_0570_ ), .D(\us31\/_0581_ ), .X(\us31\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1363_ ( .A(\us31\/_0128_ ), .B(\us31\/_0193_ ), .X(\us31\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1364_ ( .A(\us31\/_0082_ ), .B(\us31\/_0162_ ), .X(\us31\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us31/_1365_ ( .A(\us31\/_0583_ ), .B(\us31\/_0584_ ), .C_N(\us31\/_0437_ ), .Y(\us31\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us31/_1366_ ( .A(\us31\/_0150_ ), .B(\us31\/_0118_ ), .C(\us31\/_0380_ ), .Y(\us31\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us31/_1367_ ( .A_N(\us31\/_0182_ ), .B(\us31\/_0587_ ), .C(\us31\/_0323_ ), .X(\us31\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1368_ ( .A1(\us31\/_0575_ ), .A2(\us31\/_0153_ ), .B1(\us31\/_0727_ ), .B2(\us31\/_0058_ ), .Y(\us31\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1369_ ( .A1(\us31\/_0218_ ), .A2(\us31\/_0064_ ), .B1(\us31\/_0134_ ), .B2(\us31\/_0255_ ), .Y(\us31\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1370_ ( .A(\us31\/_0585_ ), .B(\us31\/_0588_ ), .C(\us31\/_0589_ ), .D(\us31\/_0590_ ), .X(\us31\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us31/_1371_ ( .A1(\us31\/_0091_ ), .A2(\us31\/_0139_ ), .B1(\us31\/_0250_ ), .Y(\us31\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1372_ ( .A1(\us31\/_0092_ ), .A2(\us31\/_0739_ ), .B1(\us31\/_0324_ ), .B2(\us31\/_0247_ ), .Y(\us31\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1373_ ( .A1(\us31\/_0144_ ), .A2(\us31\/_0153_ ), .B1(\us31\/_0683_ ), .B2(\us31\/_0292_ ), .Y(\us31\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1374_ ( .A1(\us31\/_0091_ ), .A2(\us31\/_0218_ ), .B1(\us31\/_0330_ ), .B2(\us31\/_0292_ ), .Y(\us31\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1375_ ( .A(\us31\/_0592_ ), .B(\us31\/_0593_ ), .C(\us31\/_0594_ ), .D(\us31\/_0595_ ), .X(\us31\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1376_ ( .A(\us31\/_0218_ ), .B(\us31\/_0144_ ), .Y(\us31\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1377_ ( .A(\us31\/_0312_ ), .B(\us31\/_0598_ ), .Y(\us31\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1378_ ( .A(\us31\/_0575_ ), .B(\us31\/_0147_ ), .Y(\us31\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1379_ ( .A1(\us31\/_0293_ ), .A2(\us31\/_0137_ ), .B1(\us31\/_0093_ ), .B2(\us31\/_0739_ ), .Y(\us31\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1380_ ( .A1(\us31\/_0734_ ), .A2(\us31\/_0531_ ), .B1(\us31\/_0600_ ), .C1(\us31\/_0601_ ), .Y(\us31\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1381_ ( .A1(\us31\/_0153_ ), .A2(\us31\/_0261_ ), .B1(\us31\/_0599_ ), .C1(\us31\/_0602_ ), .Y(\us31\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1382_ ( .A(\us31\/_0591_ ), .B(\us31\/_0596_ ), .C(\us31\/_0174_ ), .D(\us31\/_0603_ ), .X(\us31\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1383_ ( .A(\us31\/_0247_ ), .B(\us31\/_0144_ ), .Y(\us31\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1384_ ( .A(\us31\/_0113_ ), .B(\us31\/_0017_ ), .Y(\us31\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1385_ ( .A(\us31\/_0381_ ), .B(\us31\/_0605_ ), .C(\us31\/_0361_ ), .D(\us31\/_0606_ ), .X(\us31\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1386_ ( .A1(\us31\/_0016_ ), .A2(\us31\/_0727_ ), .B1(\us31\/_0733_ ), .Y(\us31\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1387_ ( .A1(\us31\/_0586_ ), .A2(\us31\/_0159_ ), .B1(\us31\/_0082_ ), .B2(\us31\/_0750_ ), .Y(\us31\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1388_ ( .A1(\us31\/_0142_ ), .A2(\us31\/_0162_ ), .B1(\us31\/_0079_ ), .B2(\us31\/_0054_ ), .Y(\us31\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1389_ ( .A(\us31\/_0610_ ), .B(\us31\/_0611_ ), .C(\us31\/_0105_ ), .D(\us31\/_0106_ ), .X(\us31\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1390_ ( .A1(\us31\/_0094_ ), .A2(\us31\/_0302_ ), .B1(\us31\/_0324_ ), .B2(\us31\/_0089_ ), .Y(\us31\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1391_ ( .A(\us31\/_0607_ ), .B(\us31\/_0609_ ), .C(\us31\/_0612_ ), .D(\us31\/_0613_ ), .X(\us31\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1392_ ( .A(\us31\/_0041_ ), .B(\us31\/_0170_ ), .X(\us31\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1393_ ( .A(\us31\/_0554_ ), .B(\us31\/_0027_ ), .X(\us31\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1394_ ( .A(\us31\/_0027_ ), .B(\us31\/_0261_ ), .Y(\us31\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us31/_1395_ ( .A_N(\us31\/_0616_ ), .B(\us31\/_0617_ ), .Y(\us31\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1396_ ( .A1(\us31\/_0147_ ), .A2(\us31\/_0302_ ), .B1(\us31\/_0342_ ), .C1(\us31\/_0618_ ), .Y(\us31\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1397_ ( .A(\us31\/_0614_ ), .B(\us31\/_0272_ ), .C(\us31\/_0615_ ), .D(\us31\/_0620_ ), .X(\us31\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us31/_1398_ ( .A(\us31\/_0582_ ), .B(\us31\/_0604_ ), .C(\us31\/_0621_ ), .Y(\us31\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1399_ ( .A1(\us31\/_0084_ ), .A2(\us31\/_0134_ ), .B1(\us31\/_0089_ ), .Y(\us31\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1400_ ( .A1(\us31\/_0144_ ), .A2(\us31\/_0608_ ), .A3(\us31\/_0330_ ), .B1(\us31\/_0089_ ), .Y(\us31\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1401_ ( .A1(\us31\/_0197_ ), .A2(\us31\/_0130_ ), .A3(\us31\/_0110_ ), .B1(\us31\/_0094_ ), .Y(\us31\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1402_ ( .A(\us31\/_0432_ ), .B(\us31\/_0622_ ), .C(\us31\/_0623_ ), .D(\us31\/_0624_ ), .X(\us31\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us31/_1403_ ( .A1(\us31\/_0554_ ), .A2(\us31\/_0017_ ), .A3(\us31\/_0022_ ), .B1(\us31\/_0161_ ), .X(\us31\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us31/_1404_ ( .A_N(\us31\/_0269_ ), .B(\us31\/_0170_ ), .X(\us31\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1405_ ( .A1(\us31\/_0109_ ), .A2(\us31\/_0064_ ), .A3(\us31\/_0733_ ), .B1(\us31\/_0355_ ), .Y(\us31\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us31/_1406_ ( .A_N(\us31\/_0626_ ), .B(\us31\/_0627_ ), .C(\us31\/_0353_ ), .D(\us31\/_0628_ ), .X(\us31\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1407_ ( .A1(\us31\/_0091_ ), .A2(\us31\/_0110_ ), .A3(\us31\/_0176_ ), .B1(\us31\/_0139_ ), .Y(\us31\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1408_ ( .A1(\us31\/_0020_ ), .A2(\us31\/_0261_ ), .B1(\us31\/_0147_ ), .Y(\us31\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1409_ ( .A(\us31\/_0631_ ), .B(\us31\/_0344_ ), .C(\us31\/_0421_ ), .D(\us31\/_0632_ ), .X(\us31\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us31/_1410_ ( .A1(\us31\/_0325_ ), .A2(\us31\/_0734_ ), .B1(\us31\/_0038_ ), .C1(\us31\/_0113_ ), .X(\us31\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1411_ ( .A1(\us31\/_0134_ ), .A2(\us31\/_0114_ ), .B1(\us31\/_0221_ ), .C1(\us31\/_0634_ ), .Y(\us31\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us31/_1412_ ( .A(\us31\/_0119_ ), .B_N(\us31\/_0111_ ), .Y(\us31\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1413_ ( .A1(\us31\/_0032_ ), .A2(\us31\/_0113_ ), .B1(\us31\/_0636_ ), .C1(\us31\/_0400_ ), .Y(\us31\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1414_ ( .A1(\us31\/_0731_ ), .A2(\us31\/_0293_ ), .A3(\us31\/_0251_ ), .B1(\us31\/_0099_ ), .Y(\us31\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1415_ ( .A(\us31\/_0189_ ), .B(\us31\/_0635_ ), .C(\us31\/_0637_ ), .D(\us31\/_0638_ ), .X(\us31\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1416_ ( .A(\us31\/_0625_ ), .B(\us31\/_0630_ ), .C(\us31\/_0633_ ), .D(\us31\/_0639_ ), .X(\us31\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1417_ ( .A(\us31\/_0746_ ), .B(\us31\/_0738_ ), .X(\us31\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1418_ ( .A(\us31\/_0736_ ), .B(\us31\/_0731_ ), .X(\us31\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us31/_1419_ ( .A_N(\us31\/_0643_ ), .B(\us31\/_0577_ ), .Y(\us31\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1420_ ( .A1(\us31\/_0084_ ), .A2(\us31\/_0739_ ), .B1(\us31\/_0642_ ), .C1(\us31\/_0644_ ), .Y(\us31\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1421_ ( .A1(\us31\/_0050_ ), .A2(\us31\/_0543_ ), .B1(\us31\/_0194_ ), .C1(\us31\/_0738_ ), .Y(\us31\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1422_ ( .A(\us31\/_0646_ ), .B(\us31\/_0232_ ), .C(\us31\/_0417_ ), .D(\us31\/_0578_ ), .X(\us31\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1423_ ( .A1(\us31\/_0064_ ), .A2(\us31\/_0733_ ), .B1(\us31\/_0727_ ), .Y(\us31\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1424_ ( .A1(\us31\/_0193_ ), .A2(\us31\/_0276_ ), .B1(\us31\/_0727_ ), .Y(\us31\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1425_ ( .A(\us31\/_0645_ ), .B(\us31\/_0647_ ), .C(\us31\/_0648_ ), .D(\us31\/_0649_ ), .X(\us31\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1426_ ( .A1(\us31\/_0325_ ), .A2(\us31\/_0734_ ), .B1(\us31\/_0038_ ), .C1(\us31\/_0247_ ), .Y(\us31\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1427_ ( .A1(\us31\/_0543_ ), .A2(\us31\/_0205_ ), .B1(\us31\/_0423_ ), .C1(\us31\/_0247_ ), .Y(\us31\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1428_ ( .A(\us31\/_0652_ ), .B(\us31\/_0653_ ), .X(\us31\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1429_ ( .A1(\us31\/_0733_ ), .A2(\us31\/_0748_ ), .A3(\us31\/_0324_ ), .B1(\us31\/_0016_ ), .Y(\us31\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1430_ ( .A1(\us31\/_0640_ ), .A2(\us31\/_0193_ ), .A3(\us31\/_0091_ ), .B1(\us31\/_0016_ ), .Y(\us31\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1431_ ( .A1(\us31\/_0102_ ), .A2(\us31\/_0301_ ), .B1(\sa31\[3\] ), .C1(\us31\/_0247_ ), .Y(\us31\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1432_ ( .A(\us31\/_0654_ ), .B(\us31\/_0655_ ), .C(\us31\/_0656_ ), .D(\us31\/_0657_ ), .X(\us31\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1433_ ( .A1(\us31\/_0118_ ), .A2(\us31\/_0050_ ), .B1(\us31\/_0038_ ), .C1(\us31\/_0478_ ), .Y(\us31\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us31/_1434_ ( .A_N(\us31\/_0250_ ), .B(\us31\/_0465_ ), .C(\us31\/_0659_ ), .X(\us31\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1435_ ( .A1(\us31\/_0683_ ), .A2(\us31\/_0324_ ), .B1(\us31\/_0255_ ), .Y(\us31\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1436_ ( .A1(\us31\/_0032_ ), .A2(\us31\/_0193_ ), .A3(\us31\/_0047_ ), .B1(\us31\/_0255_ ), .Y(\us31\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1437_ ( .A1(\us31\/_0144_ ), .A2(\us31\/_0586_ ), .A3(\us31\/_0047_ ), .B1(\us31\/_0218_ ), .Y(\us31\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1438_ ( .A(\us31\/_0660_ ), .B(\us31\/_0661_ ), .C(\us31\/_0663_ ), .D(\us31\/_0664_ ), .X(\us31\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1439_ ( .A1(\us31\/_0091_ ), .A2(\us31\/_0276_ ), .B1(\us31\/_0060_ ), .Y(\us31\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1440_ ( .A1(\us31\/_0144_ ), .A2(\us31\/_0608_ ), .B1(\us31\/_0292_ ), .Y(\us31\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1441_ ( .A1(\us31\/_0423_ ), .A2(\us31\/_0038_ ), .B1(\us31\/_0102_ ), .C1(\us31\/_0060_ ), .Y(\us31\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1442_ ( .A1(\sa31\[1\] ), .A2(\us31\/_0734_ ), .B1(\us31\/_0109_ ), .C1(\us31\/_0292_ ), .Y(\us31\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1443_ ( .A(\us31\/_0666_ ), .B(\us31\/_0667_ ), .C(\us31\/_0668_ ), .D(\us31\/_0669_ ), .X(\us31\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1444_ ( .A(\us31\/_0650_ ), .B(\us31\/_0658_ ), .C(\us31\/_0665_ ), .D(\us31\/_0670_ ), .X(\us31\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us31/_1445_ ( .A(\us31\/_0641_ ), .B(\us31\/_0174_ ), .C(\us31\/_0671_ ), .Y(\us31\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us31/_1446_ ( .A(\us31\/_0049_ ), .B(\us31\/_0618_ ), .C_N(\us31\/_0052_ ), .Y(\us31\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us31/_1447_ ( .A(\us31\/_0239_ ), .Y(\us31\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1448_ ( .A(\us31\/_0705_ ), .B(\us31\/_0032_ ), .Y(\us31\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1449_ ( .A1(\us31\/_0054_ ), .A2(\us31\/_0731_ ), .B1(\us31\/_0035_ ), .B2(\us31\/_0705_ ), .Y(\us31\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1450_ ( .A1(\us31\/_0304_ ), .A2(\us31\/_0731_ ), .B1(\us31\/_0047_ ), .B2(\us31\/_0750_ ), .Y(\us31\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1451_ ( .A(\us31\/_0674_ ), .B(\us31\/_0675_ ), .C(\us31\/_0676_ ), .D(\us31\/_0677_ ), .X(\us31\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us31/_1452_ ( .A_N(\us31\/_0584_ ), .B(\us31\/_0283_ ), .X(\us31\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1453_ ( .A(\us31\/_0673_ ), .B(\us31\/_0678_ ), .C(\us31\/_0679_ ), .D(\us31\/_0508_ ), .X(\us31\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1454_ ( .A1(\us31\/_0016_ ), .A2(\us31\/_0733_ ), .B1(\us31\/_0355_ ), .B2(\us31\/_0092_ ), .Y(\us31\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1455_ ( .A(\us31\/_0681_ ), .B(\us31\/_0034_ ), .X(\us31\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us31/_1456_ ( .A1(\us31\/_0330_ ), .A2(\us31\/_0139_ ), .B1(\us31\/_0324_ ), .B2(\us31\/_0089_ ), .X(\us31\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1457_ ( .A1(\us31\/_0146_ ), .A2(\us31\/_0147_ ), .B1(\us31\/_0133_ ), .C1(\us31\/_0684_ ), .Y(\us31\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1458_ ( .A(\us31\/_0113_ ), .B(\us31\/_0251_ ), .Y(\us31\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us31/_1459_ ( .A_N(\us31\/_0463_ ), .B(\us31\/_0686_ ), .C(\us31\/_0383_ ), .D(\us31\/_0464_ ), .X(\us31\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1460_ ( .A1(\us31\/_0051_ ), .A2(\us31\/_0293_ ), .B1(\us31\/_0084_ ), .B2(\us31\/_0705_ ), .Y(\us31\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1461_ ( .A1(\us31\/_0017_ ), .A2(\us31\/_0072_ ), .B1(\us31\/_0134_ ), .B2(\us31\/_0078_ ), .Y(\us31\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1462_ ( .A(\us31\/_0687_ ), .B(\us31\/_0236_ ), .C(\us31\/_0688_ ), .D(\us31\/_0689_ ), .X(\us31\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1463_ ( .A(\us31\/_0680_ ), .B(\us31\/_0682_ ), .C(\us31\/_0685_ ), .D(\us31\/_0690_ ), .X(\us31\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us31/_1464_ ( .A1(\us31\/_0532_ ), .A2(\us31\/_0380_ ), .B1(\us31\/_0102_ ), .C1(\us31\/_0355_ ), .X(\us31\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us31/_1465_ ( .A(\us31\/_0692_ ), .B(\us31\/_0338_ ), .C(\us31\/_0644_ ), .Y(\us31\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1466_ ( .A(\us31\/_0016_ ), .B(\us31\/_0020_ ), .Y(\us31\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1467_ ( .A1(\us31\/_0032_ ), .A2(\us31\/_0137_ ), .B1(\us31\/_0279_ ), .B2(\us31\/_0094_ ), .Y(\us31\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1468_ ( .A1(\us31\/_0575_ ), .A2(\us31\/_0153_ ), .B1(\us31\/_0161_ ), .B2(\us31\/_0293_ ), .Y(\us31\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1469_ ( .A(\us31\/_0259_ ), .B(\us31\/_0695_ ), .C(\us31\/_0696_ ), .D(\us31\/_0697_ ), .X(\us31\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us31/_1470_ ( .A1(\us31\/_0255_ ), .A2(\us31\/_0640_ ), .B1(\us31\/_0016_ ), .B2(\us31\/_0193_ ), .X(\us31\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1471_ ( .A1(\us31\/_0060_ ), .A2(\us31\/_0176_ ), .B1(\us31\/_0699_ ), .C1(\us31\/_0177_ ), .Y(\us31\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1472_ ( .A1(\us31\/_0091_ ), .A2(\us31\/_0218_ ), .B1(\us31\/_0092_ ), .B2(\us31\/_0705_ ), .Y(\us31\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us31/_1473_ ( .A1(\us31\/_0705_ ), .A2(\us31\/_0683_ ), .B1(\us31\/_0093_ ), .B2(\us31\/_0114_ ), .Y(\us31\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us31/_1474_ ( .A1(\us31\/_0683_ ), .A2(\us31\/_0084_ ), .B1(\us31\/_0094_ ), .Y(\us31\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us31/_1475_ ( .A1(\us31\/_0543_ ), .A2(\us31\/_0205_ ), .B1(\us31\/_0038_ ), .C1(\us31\/_0292_ ), .Y(\us31\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1476_ ( .A(\us31\/_0701_ ), .B(\us31\/_0702_ ), .C(\us31\/_0703_ ), .D(\us31\/_0704_ ), .X(\us31\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1477_ ( .A(\us31\/_0693_ ), .B(\us31\/_0698_ ), .C(\us31\/_0700_ ), .D(\us31\/_0706_ ), .X(\us31\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us31/_1478_ ( .A1(\us31\/_0113_ ), .A2(\us31\/_0640_ ), .B1(\us31\/_0099_ ), .B2(\us31\/_0058_ ), .X(\us31\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us31/_1479_ ( .A(\us31\/_0407_ ), .B(\us31\/_0708_ ), .C(\us31\/_0529_ ), .Y(\us31\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1480_ ( .A(\us31\/_0568_ ), .B(\us31\/_0175_ ), .Y(\us31\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us31/_1481_ ( .A1(\us31\/_0247_ ), .A2(\us31\/_0114_ ), .A3(\us31\/_0051_ ), .B1(\us31\/_0130_ ), .Y(\us31\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1482_ ( .A(\us31\/_0709_ ), .B(\us31\/_0550_ ), .C(\us31\/_0710_ ), .D(\us31\/_0711_ ), .X(\us31\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us31/_1483_ ( .A1(\us31\/_0114_ ), .A2(\us31\/_0064_ ), .B1(\us31\/_0261_ ), .B2(\us31\/_0089_ ), .X(\us31\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1484_ ( .A1(\us31\/_0355_ ), .A2(\us31\/_0261_ ), .B1(\us31\/_0198_ ), .C1(\us31\/_0713_ ), .Y(\us31\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1485_ ( .A(\us31\/_0586_ ), .B(\us31\/_0478_ ), .Y(\us31\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us31/_1486_ ( .A_N(\us31\/_0541_ ), .B(\us31\/_0267_ ), .C(\us31\/_0715_ ), .D(\us31\/_0320_ ), .X(\us31\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1487_ ( .A(\us31\/_0586_ ), .B(\us31\/_0070_ ), .Y(\us31\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us31/_1488_ ( .A_N(\us31\/_0211_ ), .B(\us31\/_0155_ ), .C(\us31\/_0202_ ), .D(\us31\/_0718_ ), .X(\us31\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us31/_1489_ ( .A(\us31\/_0150_ ), .B(\us31\/_0205_ ), .C(\us31\/_0380_ ), .Y(\us31\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us31/_1490_ ( .A(\us31\/_0411_ ), .B(\us31\/_0720_ ), .X(\us31\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us31/_1491_ ( .A1(\us31\/_0017_ ), .A2(\us31\/_0022_ ), .B1(\us31\/_0078_ ), .X(\us31\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us31/_1492_ ( .A1(\us31\/_0134_ ), .A2(\us31\/_0738_ ), .B1(\us31\/_0101_ ), .C1(\us31\/_0722_ ), .Y(\us31\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1493_ ( .A(\us31\/_0717_ ), .B(\us31\/_0719_ ), .C(\us31\/_0721_ ), .D(\us31\/_0723_ ), .X(\us31\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us31/_1494_ ( .A(\us31\/_0739_ ), .B(\us31\/_0193_ ), .Y(\us31\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1495_ ( .A(\us31\/_0344_ ), .B(\us31\/_0184_ ), .C(\us31\/_0449_ ), .D(\us31\/_0725_ ), .X(\us31\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us31/_1496_ ( .A(\us31\/_0712_ ), .B(\us31\/_0714_ ), .C(\us31\/_0724_ ), .D(\us31\/_0726_ ), .X(\us31\/_0728_ ) );
sky130_fd_sc_hd__nand3_2 \us31/_1497_ ( .A(\us31\/_0691_ ), .B(\us31\/_0707_ ), .C(\us31\/_0728_ ), .Y(\us31\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \us32/_0753_ ( .A(\sa32\[2\] ), .B_N(\sa32\[3\] ), .Y(\us32\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \us32/_0755_ ( .A(\sa32\[1\] ), .B(\sa32\[0\] ), .X(\us32\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us32/_0756_ ( .A(\us32\/_0096_ ), .B(\us32\/_0118_ ), .X(\us32\/_0129_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0757_ ( .A(\sa32\[7\] ), .B(\sa32\[6\] ), .X(\us32\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_0758_ ( .A(\sa32\[4\] ), .B(\sa32\[5\] ), .Y(\us32\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0759_ ( .A(\us32\/_0140_ ), .B(\us32\/_0151_ ), .X(\us32\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0761_ ( .A(\us32\/_0129_ ), .B(\us32\/_0162_ ), .X(\us32\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0762_ ( .A(\us32\/_0096_ ), .X(\us32\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \us32/_0763_ ( .A(\sa32\[1\] ), .B_N(\sa32\[0\] ), .Y(\us32\/_0205_ ) );
sky130_fd_sc_hd__and3_1 \us32/_0765_ ( .A(\us32\/_0162_ ), .B(\us32\/_0194_ ), .C(\us32\/_0205_ ), .X(\us32\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us32/_0766_ ( .A(\us32\/_0183_ ), .SLEEP(\us32\/_0227_ ), .X(\us32\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \us32/_0767_ ( .A(\sa32\[0\] ), .B_N(\sa32\[1\] ), .Y(\us32\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_0768_ ( .A(\sa32\[2\] ), .B(\sa32\[3\] ), .Y(\us32\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0769_ ( .A(\us32\/_0249_ ), .B(\us32\/_0260_ ), .X(\us32\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0771_ ( .A(\us32\/_0271_ ), .X(\us32\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0772_ ( .A(\us32\/_0162_ ), .X(\us32\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_0773_ ( .A(\us32\/_0293_ ), .B(\us32\/_0304_ ), .Y(\us32\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us32/_0774_ ( .A(\sa32\[1\] ), .Y(\us32\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us32/_0776_ ( .A(\sa32\[0\] ), .Y(\us32\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0777_ ( .A(\sa32\[2\] ), .B(\sa32\[3\] ), .X(\us32\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0779_ ( .A(\us32\/_0358_ ), .X(\us32\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_0780_ ( .A1(\us32\/_0325_ ), .A2(\us32\/_0347_ ), .B1(\us32\/_0380_ ), .C1(\us32\/_0304_ ), .Y(\us32\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us32/_0781_ ( .A_N(\us32\/_0238_ ), .B(\us32\/_0314_ ), .C(\us32\/_0391_ ), .X(\us32\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us32/_0782_ ( .A(\sa32\[3\] ), .B_N(\sa32\[2\] ), .Y(\us32\/_0412_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0784_ ( .A(\us32\/_0412_ ), .B(\us32\/_0205_ ), .X(\us32\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \us32/_0787_ ( .A(\sa32\[5\] ), .B_N(\sa32\[4\] ), .Y(\us32\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0788_ ( .A(\us32\/_0467_ ), .B(\us32\/_0140_ ), .X(\us32\/_0478_ ) );
sky130_fd_sc_hd__buf_2 \us32/_0790_ ( .A(\us32\/_0478_ ), .X(\us32\/_0499_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_0791_ ( .A(\us32\/_0134_ ), .B(\us32\/_0499_ ), .Y(\us32\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_0792_ ( .A(\us32\/_0478_ ), .B(\us32\/_0271_ ), .Y(\us32\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0793_ ( .A(\us32\/_0194_ ), .X(\us32\/_0532_ ) );
sky130_fd_sc_hd__and2_1 \us32/_0795_ ( .A(\us32\/_0249_ ), .B(\us32\/_0358_ ), .X(\us32\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0797_ ( .A(\us32\/_0554_ ), .X(\us32\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us32/_0798_ ( .A(\us32\/_0205_ ), .B(\us32\/_0358_ ), .X(\us32\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0800_ ( .A(\us32\/_0586_ ), .X(\us32\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_0801_ ( .A1(\us32\/_0532_ ), .A2(\us32\/_0575_ ), .A3(\us32\/_0608_ ), .B1(\us32\/_0499_ ), .Y(\us32\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us32/_0802_ ( .A(\us32\/_0401_ ), .B(\us32\/_0510_ ), .C(\us32\/_0521_ ), .D(\us32\/_0619_ ), .X(\us32\/_0629_ ) );
sky130_fd_sc_hd__and2_1 \us32/_0803_ ( .A(\us32\/_0358_ ), .B(\sa32\[1\] ), .X(\us32\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0805_ ( .A(\us32\/_0205_ ), .B(\us32\/_0260_ ), .X(\us32\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0807_ ( .A(\us32\/_0662_ ), .X(\us32\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us32/_0808_ ( .A(\sa32\[6\] ), .B_N(\sa32\[7\] ), .Y(\us32\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \us32/_0809_ ( .A(\us32\/_0467_ ), .B(\us32\/_0694_ ), .X(\us32\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0811_ ( .A(\us32\/_0705_ ), .X(\us32\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_0812_ ( .A1(\us32\/_0640_ ), .A2(\us32\/_0293_ ), .A3(\us32\/_0683_ ), .B1(\us32\/_0727_ ), .Y(\us32\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_0813_ ( .A(\sa32\[1\] ), .B(\sa32\[0\] ), .Y(\us32\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0814_ ( .A(\us32\/_0730_ ), .B(\us32\/_0260_ ), .X(\us32\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0816_ ( .A(\us32\/_0731_ ), .X(\us32\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0817_ ( .A(\sa32\[0\] ), .X(\us32\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us32/_0818_ ( .A1(\us32\/_0325_ ), .A2(\us32\/_0734_ ), .B1(\us32\/_0412_ ), .X(\us32\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0819_ ( .A(\us32\/_0694_ ), .B(\us32\/_0151_ ), .X(\us32\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0821_ ( .A(\us32\/_0736_ ), .X(\us32\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0822_ ( .A(\us32\/_0738_ ), .X(\us32\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_0823_ ( .A1(\us32\/_0733_ ), .A2(\us32\/_0735_ ), .A3(\us32\/_0293_ ), .B1(\us32\/_0739_ ), .Y(\us32\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us32/_0824_ ( .A(\us32\/_0730_ ), .B_N(\us32\/_0358_ ), .Y(\us32\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_0825_ ( .A(\us32\/_0741_ ), .B(\us32\/_0739_ ), .Y(\us32\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_0827_ ( .A1(\us32\/_0118_ ), .A2(\us32\/_0205_ ), .B1(\us32\/_0532_ ), .C1(\us32\/_0739_ ), .Y(\us32\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us32/_0828_ ( .A(\us32\/_0729_ ), .B(\us32\/_0740_ ), .C(\us32\/_0742_ ), .D(\us32\/_0744_ ), .X(\us32\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0829_ ( .A(\us32\/_0412_ ), .B(\us32\/_0730_ ), .X(\us32\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0831_ ( .A(\us32\/_0746_ ), .X(\us32\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us32/_0832_ ( .A(\sa32\[4\] ), .B_N(\sa32\[5\] ), .Y(\us32\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0833_ ( .A(\us32\/_0749_ ), .B(\us32\/_0694_ ), .X(\us32\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0835_ ( .A(\us32\/_0750_ ), .X(\us32\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0836_ ( .A(\us32\/_0752_ ), .X(\us32\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0837_ ( .A(\us32\/_0118_ ), .B(\us32\/_0358_ ), .X(\us32\/_0017_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0839_ ( .A(\us32\/_0752_ ), .B(\us32\/_0017_ ), .X(\us32\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0840_ ( .A(\us32\/_0358_ ), .B(\us32\/_0325_ ), .X(\us32\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0842_ ( .A(\us32\/_0096_ ), .B(\us32\/_0205_ ), .X(\us32\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \us32/_0844_ ( .A1(\us32\/_0020_ ), .A2(\us32\/_0022_ ), .B1(\us32\/_0752_ ), .X(\us32\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_0845_ ( .A1(\us32\/_0748_ ), .A2(\us32\/_0016_ ), .B1(\us32\/_0019_ ), .C1(\us32\/_0024_ ), .Y(\us32\/_0025_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0846_ ( .A(\sa32\[4\] ), .B(\sa32\[5\] ), .X(\us32\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0847_ ( .A(\us32\/_0694_ ), .B(\us32\/_0026_ ), .X(\us32\/_0027_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0850_ ( .A(\us32\/_0358_ ), .B(\us32\/_0730_ ), .X(\us32\/_0030_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0852_ ( .A(\us32\/_0030_ ), .X(\us32\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_0853_ ( .A(\us32\/_0247_ ), .B(\us32\/_0032_ ), .Y(\us32\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_0854_ ( .A(\us32\/_0247_ ), .B(\us32\/_0735_ ), .Y(\us32\/_0034_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0855_ ( .A(\us32\/_0118_ ), .B(\us32\/_0260_ ), .X(\us32\/_0035_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0857_ ( .A(\us32\/_0027_ ), .B(\us32\/_0035_ ), .X(\us32\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0858_ ( .A(\us32\/_0260_ ), .X(\us32\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_0859_ ( .A(\us32\/_0038_ ), .B(\us32\/_0347_ ), .Y(\us32\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us32/_0860_ ( .A_N(\us32\/_0039_ ), .B(\us32\/_0027_ ), .X(\us32\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_0861_ ( .A(\us32\/_0037_ ), .B(\us32\/_0040_ ), .Y(\us32\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us32/_0862_ ( .A(\us32\/_0025_ ), .B(\us32\/_0033_ ), .C(\us32\/_0034_ ), .D(\us32\/_0041_ ), .X(\us32\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0863_ ( .A(\us32\/_0749_ ), .B(\us32\/_0140_ ), .X(\us32\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us32/_0865_ ( .A(\sa32\[0\] ), .B(\sa32\[2\] ), .C(\sa32\[3\] ), .X(\us32\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0866_ ( .A(\us32\/_0043_ ), .B(\us32\/_0045_ ), .X(\us32\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0867_ ( .A(\us32\/_0096_ ), .B(\us32\/_0249_ ), .X(\us32\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0869_ ( .A(\us32\/_0047_ ), .B(\us32\/_0043_ ), .X(\us32\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0870_ ( .A(\us32\/_0730_ ), .X(\us32\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0871_ ( .A(\us32\/_0043_ ), .X(\us32\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_0872_ ( .A1(\us32\/_0118_ ), .A2(\us32\/_0050_ ), .B1(\us32\/_0194_ ), .C1(\us32\/_0051_ ), .Y(\us32\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us32/_0873_ ( .A(\us32\/_0046_ ), .B(\us32\/_0049_ ), .C_N(\us32\/_0052_ ), .Y(\us32\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0874_ ( .A(\us32\/_0026_ ), .B(\us32\/_0140_ ), .X(\us32\/_0054_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0876_ ( .A(\us32\/_0054_ ), .X(\us32\/_0056_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_0877_ ( .A1(\us32\/_0532_ ), .A2(\us32\/_0575_ ), .B1(\us32\/_0056_ ), .Y(\us32\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0878_ ( .A(\us32\/_0412_ ), .B(\us32\/_0325_ ), .X(\us32\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0880_ ( .A(\us32\/_0051_ ), .X(\us32\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_0881_ ( .A1(\us32\/_0731_ ), .A2(\us32\/_0035_ ), .A3(\us32\/_0058_ ), .B1(\us32\/_0060_ ), .Y(\us32\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0882_ ( .A(\us32\/_0260_ ), .B(\sa32\[1\] ), .X(\us32\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0884_ ( .A(\us32\/_0062_ ), .X(\us32\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_0885_ ( .A1(\us32\/_0064_ ), .A2(\us32\/_0748_ ), .A3(\us32\/_0683_ ), .B1(\us32\/_0056_ ), .Y(\us32\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us32/_0886_ ( .A(\us32\/_0053_ ), .B(\us32\/_0057_ ), .C(\us32\/_0061_ ), .D(\us32\/_0065_ ), .X(\us32\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us32/_0887_ ( .A(\us32\/_0629_ ), .B(\us32\/_0745_ ), .C(\us32\/_0042_ ), .D(\us32\/_0066_ ), .X(\us32\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us32/_0889_ ( .A(\sa32\[7\] ), .B_N(\sa32\[6\] ), .Y(\us32\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0890_ ( .A(\us32\/_0069_ ), .B(\us32\/_0151_ ), .X(\us32\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0892_ ( .A(\us32\/_0070_ ), .X(\us32\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_0893_ ( .A1(\us32\/_0129_ ), .A2(\us32\/_0586_ ), .B1(\us32\/_0072_ ), .Y(\us32\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_0894_ ( .A1(\us32\/_0380_ ), .A2(\us32\/_0347_ ), .B1(\us32\/_0194_ ), .B2(\us32\/_0205_ ), .Y(\us32\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us32/_0895_ ( .A(\us32\/_0074_ ), .B_N(\us32\/_0070_ ), .Y(\us32\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us32/_0896_ ( .A(\us32\/_0073_ ), .SLEEP(\us32\/_0075_ ), .X(\us32\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us32/_0897_ ( .A(\us32\/_0467_ ), .B(\us32\/_0069_ ), .X(\us32\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0898_ ( .A(\us32\/_0077_ ), .X(\us32\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0899_ ( .A(\us32\/_0412_ ), .B(\us32\/_0118_ ), .X(\us32\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0901_ ( .A(\us32\/_0078_ ), .B(\us32\/_0079_ ), .X(\us32\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0902_ ( .A(\us32\/_0412_ ), .B(\us32\/_0249_ ), .X(\us32\/_0082_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0905_ ( .A(\us32\/_0280_ ), .B(\us32\/_0078_ ), .X(\us32\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us32/_0906_ ( .A1(\sa32\[0\] ), .A2(\us32\/_0325_ ), .B1(\us32\/_0260_ ), .Y(\us32\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us32/_0907_ ( .A_N(\us32\/_0086_ ), .B(\us32\/_0078_ ), .X(\us32\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us32/_0908_ ( .A(\us32\/_0081_ ), .B(\us32\/_0085_ ), .C(\us32\/_0087_ ), .Y(\us32\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0909_ ( .A(\us32\/_0072_ ), .X(\us32\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_0910_ ( .A1(\us32\/_0733_ ), .A2(\us32\/_0748_ ), .A3(\us32\/_0683_ ), .B1(\us32\/_0089_ ), .Y(\us32\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0911_ ( .A(\us32\/_0129_ ), .X(\us32\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0912_ ( .A(\us32\/_0017_ ), .X(\us32\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0913_ ( .A(\us32\/_0022_ ), .X(\us32\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0914_ ( .A(\us32\/_0078_ ), .X(\us32\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_0915_ ( .A1(\us32\/_0091_ ), .A2(\us32\/_0092_ ), .A3(\us32\/_0093_ ), .B1(\us32\/_0094_ ), .Y(\us32\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us32/_0916_ ( .A(\us32\/_0076_ ), .B(\us32\/_0088_ ), .C(\us32\/_0090_ ), .D(\us32\/_0095_ ), .X(\us32\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us32/_0917_ ( .A(\us32\/_0069_ ), .B(\us32\/_0026_ ), .X(\us32\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \us32/_0918_ ( .A(\us32\/_0098_ ), .X(\us32\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0919_ ( .A(\us32\/_0434_ ), .B(\us32\/_0099_ ), .X(\us32\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0920_ ( .A(\us32\/_0079_ ), .B(\us32\/_0098_ ), .X(\us32\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0921_ ( .A(\us32\/_0325_ ), .X(\us32\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_0922_ ( .A1(\us32\/_0102_ ), .A2(\us32\/_0734_ ), .B1(\us32\/_0038_ ), .C1(\us32\/_0099_ ), .Y(\us32\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us32/_0923_ ( .A(\us32\/_0100_ ), .B(\us32\/_0101_ ), .C_N(\us32\/_0103_ ), .Y(\us32\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_0924_ ( .A1(\us32\/_0554_ ), .A2(\us32\/_0586_ ), .B1(\us32\/_0099_ ), .Y(\us32\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_0925_ ( .A(\us32\/_0129_ ), .B(\us32\/_0099_ ), .Y(\us32\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0926_ ( .A(\us32\/_0105_ ), .B(\us32\/_0106_ ), .X(\us32\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0927_ ( .A(\us32\/_0412_ ), .X(\us32\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us32/_0928_ ( .A(\us32\/_0260_ ), .B(\sa32\[0\] ), .X(\us32\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0929_ ( .A(\us32\/_0069_ ), .B(\us32\/_0749_ ), .X(\us32\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0931_ ( .A(\us32\/_0111_ ), .X(\us32\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0932_ ( .A(\us32\/_0113_ ), .X(\us32\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_0933_ ( .A1(\us32\/_0109_ ), .A2(\us32\/_0110_ ), .B1(\us32\/_0114_ ), .Y(\us32\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us32/_0934_ ( .A(\us32\/_0022_ ), .Y(\us32\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us32/_0935_ ( .A(\us32\/_0554_ ), .Y(\us32\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us32/_0936_ ( .A1(\us32\/_0050_ ), .A2(\us32\/_0118_ ), .B1(\us32\/_0194_ ), .Y(\us32\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us32/_0937_ ( .A(\us32\/_0113_ ), .Y(\us32\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us32/_0938_ ( .A1(\us32\/_0116_ ), .A2(\us32\/_0117_ ), .A3(\us32\/_0119_ ), .B1(\us32\/_0120_ ), .X(\us32\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us32/_0939_ ( .A(\us32\/_0104_ ), .B(\us32\/_0108_ ), .C(\us32\/_0115_ ), .D(\us32\/_0121_ ), .X(\us32\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_0940_ ( .A(\sa32\[7\] ), .B(\sa32\[6\] ), .Y(\us32\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0941_ ( .A(\us32\/_0749_ ), .B(\us32\/_0123_ ), .X(\us32\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0943_ ( .A(\us32\/_0082_ ), .B(\us32\/_0124_ ), .X(\us32\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_0944_ ( .A(\us32\/_0271_ ), .B(\us32\/_0124_ ), .Y(\us32\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0945_ ( .A(\us32\/_0124_ ), .X(\us32\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0946_ ( .A(\us32\/_0260_ ), .B(\us32\/_0325_ ), .X(\us32\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_0948_ ( .A(\us32\/_0128_ ), .B(\us32\/_0130_ ), .Y(\us32\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_0949_ ( .A(\us32\/_0127_ ), .B(\us32\/_0132_ ), .Y(\us32\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us32/_0950_ ( .A(\us32\/_0434_ ), .X(\us32\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_0951_ ( .A(\us32\/_0134_ ), .B(\us32\/_0128_ ), .Y(\us32\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us32/_0952_ ( .A(\us32\/_0126_ ), .B(\us32\/_0133_ ), .C_N(\us32\/_0135_ ), .Y(\us32\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us32/_0953_ ( .A(\us32\/_0026_ ), .B(\us32\/_0123_ ), .X(\us32\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0955_ ( .A(\us32\/_0137_ ), .X(\us32\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_0956_ ( .A1(\us32\/_0110_ ), .A2(\us32\/_0293_ ), .A3(\us32\/_0280_ ), .B1(\us32\/_0139_ ), .Y(\us32\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0957_ ( .A(\us32\/_0096_ ), .B(\us32\/_0730_ ), .X(\us32\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0959_ ( .A(\us32\/_0142_ ), .X(\us32\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_0960_ ( .A1(\us32\/_0020_ ), .A2(\us32\/_0144_ ), .A3(\us32\/_0017_ ), .B1(\us32\/_0139_ ), .Y(\us32\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \us32/_0961_ ( .A(\sa32\[2\] ), .B(\us32\/_0050_ ), .C_N(\sa32\[3\] ), .Y(\us32\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0962_ ( .A(\us32\/_0128_ ), .X(\us32\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_0963_ ( .A1(\us32\/_0146_ ), .A2(\us32\/_0032_ ), .A3(\us32\/_0640_ ), .B1(\us32\/_0147_ ), .Y(\us32\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us32/_0964_ ( .A(\us32\/_0136_ ), .B(\us32\/_0141_ ), .C(\us32\/_0145_ ), .D(\us32\/_0148_ ), .X(\us32\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0965_ ( .A(\us32\/_0123_ ), .B(\us32\/_0151_ ), .X(\us32\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0967_ ( .A(\us32\/_0150_ ), .X(\us32\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \us32/_0968_ ( .A(\us32\/_0150_ ), .B(\us32\/_0062_ ), .X(\us32\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_0969_ ( .A(\us32\/_0079_ ), .B(\us32\/_0150_ ), .Y(\us32\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us32/_0970_ ( .A(\us32\/_0150_ ), .B(\us32\/_0412_ ), .C(\us32\/_0249_ ), .Y(\us32\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_0971_ ( .A(\us32\/_0155_ ), .B(\us32\/_0156_ ), .Y(\us32\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_0972_ ( .A1(\us32\/_0153_ ), .A2(\us32\/_0134_ ), .B1(\us32\/_0154_ ), .C1(\us32\/_0157_ ), .Y(\us32\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0973_ ( .A(\us32\/_0467_ ), .B(\us32\/_0123_ ), .X(\us32\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_0975_ ( .A(\us32\/_0159_ ), .X(\us32\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us32/_0976_ ( .A_N(\us32\/_0119_ ), .B(\us32\/_0161_ ), .X(\us32\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us32/_0977_ ( .A(\us32\/_0163_ ), .Y(\us32\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_0978_ ( .A1(\us32\/_0146_ ), .A2(\us32\/_0575_ ), .A3(\us32\/_0608_ ), .B1(\us32\/_0153_ ), .Y(\us32\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_0979_ ( .A1(\us32\/_0062_ ), .A2(\us32\/_0280_ ), .A3(\us32\/_0134_ ), .B1(\us32\/_0161_ ), .Y(\us32\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us32/_0980_ ( .A(\us32\/_0158_ ), .B(\us32\/_0164_ ), .C(\us32\/_0165_ ), .D(\us32\/_0166_ ), .X(\us32\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us32/_0981_ ( .A(\us32\/_0097_ ), .B(\us32\/_0122_ ), .C(\us32\/_0149_ ), .D(\us32\/_0167_ ), .X(\us32\/_0168_ ) );
sky130_fd_sc_hd__and2_1 \us32/_0982_ ( .A(\us32\/_0662_ ), .B(\us32\/_0150_ ), .X(\us32\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_0983_ ( .A(\us32\/_0154_ ), .B(\us32\/_0169_ ), .Y(\us32\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us32/_0984_ ( .A(\us32\/_0123_ ), .B(\us32\/_0151_ ), .C(\us32\/_0038_ ), .X(\us32\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0985_ ( .A(\us32\/_0170_ ), .B(\us32\/_0171_ ), .X(\us32\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \us32/_0986_ ( .A(\us32\/_0172_ ), .Y(\us32\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \us32/_0987_ ( .A(\us32\/_0067_ ), .B(\us32\/_0168_ ), .C(\us32\/_0174_ ), .Y(\us32\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us32/_0988_ ( .A(\sa32\[1\] ), .B(\sa32\[0\] ), .Y(\us32\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us32/_0989_ ( .A(\us32\/_0175_ ), .B(\us32\/_0358_ ), .X(\us32\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0990_ ( .A(\us32\/_0176_ ), .B(\us32\/_0478_ ), .X(\us32\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_0991_ ( .A(\us32\/_0280_ ), .B(\us32\/_0113_ ), .Y(\us32\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0992_ ( .A(\us32\/_0111_ ), .B(\us32\/_0062_ ), .X(\us32\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0993_ ( .A(\us32\/_0111_ ), .B(\us32\/_0662_ ), .X(\us32\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_0994_ ( .A(\us32\/_0179_ ), .B(\us32\/_0180_ ), .Y(\us32\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0995_ ( .A(\us32\/_0054_ ), .B(\us32\/_0058_ ), .X(\us32\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us32/_0996_ ( .A(\us32\/_0182_ ), .Y(\us32\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us32/_0997_ ( .A_N(\us32\/_0177_ ), .B(\us32\/_0178_ ), .C(\us32\/_0181_ ), .D(\us32\/_0184_ ), .X(\us32\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0998_ ( .A(\us32\/_0098_ ), .B(\us32\/_0741_ ), .X(\us32\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us32/_0999_ ( .A(\us32\/_0047_ ), .B(\us32\/_0098_ ), .X(\us32\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us32/_1000_ ( .A(\us32\/_0186_ ), .B(\us32\/_0187_ ), .X(\us32\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1001_ ( .A(\us32\/_0188_ ), .Y(\us32\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1002_ ( .A(\us32\/_0738_ ), .B(\us32\/_0735_ ), .X(\us32\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1003_ ( .A(\us32\/_0271_ ), .B(\us32\/_0736_ ), .X(\us32\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_1004_ ( .A(\us32\/_0190_ ), .B(\us32\/_0191_ ), .Y(\us32\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us32/_1005_ ( .A(\us32\/_0096_ ), .B(\us32\/_0325_ ), .X(\us32\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1006_ ( .A1(\us32\/_0193_ ), .A2(\us32\/_0176_ ), .B1(\us32\/_0043_ ), .Y(\us32\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1007_ ( .A(\us32\/_0185_ ), .B(\us32\/_0189_ ), .C(\us32\/_0192_ ), .D(\us32\/_0195_ ), .X(\us32\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us32/_1008_ ( .A_N(\sa32\[3\] ), .B(\us32\/_0734_ ), .C(\sa32\[2\] ), .X(\us32\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1009_ ( .A(\us32\/_0137_ ), .B(\us32\/_0197_ ), .X(\us32\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_1010_ ( .A(\us32\/_0198_ ), .B(\us32\/_0040_ ), .Y(\us32\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1011_ ( .A(\us32\/_0293_ ), .B(\us32\/_0137_ ), .X(\us32\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1012_ ( .A(\us32\/_0200_ ), .Y(\us32\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1013_ ( .A(\us32\/_0137_ ), .B(\us32\/_0110_ ), .Y(\us32\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1014_ ( .A(\us32\/_0139_ ), .B(\us32\/_0020_ ), .Y(\us32\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1015_ ( .A(\us32\/_0199_ ), .B(\us32\/_0201_ ), .C(\us32\/_0202_ ), .D(\us32\/_0203_ ), .X(\us32\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us32/_1016_ ( .A1(\us32\/_0532_ ), .A2(\us32\/_0109_ ), .B1(\us32\/_0102_ ), .C1(\us32\/_0727_ ), .X(\us32\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1017_ ( .A(\us32\/_0022_ ), .B(\us32\/_0078_ ), .Y(\us32\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1018_ ( .A(\us32\/_0078_ ), .B(\us32\/_0142_ ), .Y(\us32\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1019_ ( .A(\us32\/_0207_ ), .B(\us32\/_0208_ ), .Y(\us32\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1020_ ( .A1(\us32\/_0094_ ), .A2(\us32\/_0176_ ), .B1(\us32\/_0206_ ), .C1(\us32\/_0209_ ), .Y(\us32\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1021_ ( .A(\us32\/_0662_ ), .B(\us32\/_0070_ ), .X(\us32\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us32/_1022_ ( .A(\us32\/_0731_ ), .B(\us32\/_0123_ ), .C(\us32\/_0749_ ), .Y(\us32\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us32/_1023_ ( .A(\us32\/_0731_ ), .B(\us32\/_0467_ ), .C(\us32\/_0069_ ), .Y(\us32\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us32/_1024_ ( .A_N(\us32\/_0211_ ), .B(\us32\/_0127_ ), .C(\us32\/_0212_ ), .D(\us32\/_0213_ ), .X(\us32\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1025_ ( .A(\us32\/_0137_ ), .Y(\us32\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1026_ ( .A(\us32\/_0128_ ), .B(\us32\/_0035_ ), .Y(\us32\/_0217_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1028_ ( .A1(\us32\/_0159_ ), .A2(\us32\/_0746_ ), .B1(\us32\/_0434_ ), .B2(\us32\/_0499_ ), .Y(\us32\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us32/_1029_ ( .A1(\us32\/_0116_ ), .A2(\us32\/_0215_ ), .B1(\us32\/_0217_ ), .C1(\us32\/_0219_ ), .X(\us32\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1030_ ( .A(\us32\/_0113_ ), .B(\us32\/_0746_ ), .X(\us32\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us32/_1031_ ( .A1(\us32\/_0098_ ), .A2(\us32\/_0746_ ), .B1(\us32\/_0434_ ), .B2(\us32\/_0750_ ), .X(\us32\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1032_ ( .A1(\us32\/_0047_ ), .A2(\us32\/_0113_ ), .B1(\us32\/_0221_ ), .C1(\us32\/_0222_ ), .Y(\us32\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us32/_1033_ ( .A1(\us32\/_0129_ ), .A2(\us32\/_0162_ ), .B1(\us32\/_0271_ ), .B2(\us32\/_0705_ ), .X(\us32\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1034_ ( .A1(\us32\/_0093_ ), .A2(\us32\/_0738_ ), .B1(\us32\/_0081_ ), .C1(\us32\/_0224_ ), .Y(\us32\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1035_ ( .A(\us32\/_0214_ ), .B(\us32\/_0220_ ), .C(\us32\/_0223_ ), .D(\us32\/_0225_ ), .X(\us32\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1036_ ( .A(\us32\/_0196_ ), .B(\us32\/_0204_ ), .C(\us32\/_0210_ ), .D(\us32\/_0226_ ), .X(\us32\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1037_ ( .A(\us32\/_0111_ ), .B(\us32\/_0554_ ), .X(\us32\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1038_ ( .A(\us32\/_0229_ ), .Y(\us32\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1039_ ( .A(\us32\/_0111_ ), .B(\us32\/_0129_ ), .Y(\us32\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1040_ ( .A(\us32\/_0017_ ), .B(\us32\/_0738_ ), .Y(\us32\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1041_ ( .A(\us32\/_0030_ ), .B(\us32\/_0304_ ), .Y(\us32\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1042_ ( .A(\us32\/_0230_ ), .B(\us32\/_0231_ ), .C(\us32\/_0232_ ), .D(\us32\/_0233_ ), .X(\us32\/_0234_ ) );
sky130_fd_sc_hd__and2_1 \us32/_1043_ ( .A(\us32\/_0047_ ), .B(\us32\/_0478_ ), .X(\us32\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1044_ ( .A1(\us32\/_0129_ ), .A2(\us32\/_0554_ ), .B1(\us32\/_0137_ ), .Y(\us32\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us32/_1045_ ( .A(\us32\/_0235_ ), .B(\us32\/_0049_ ), .C_N(\us32\/_0236_ ), .Y(\us32\/_0237_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1046_ ( .A(\us32\/_0047_ ), .B(\us32\/_0077_ ), .X(\us32\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1047_ ( .A(\us32\/_0070_ ), .B(\us32\/_0035_ ), .X(\us32\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us32/_1048_ ( .A1(\us32\/_0047_ ), .A2(\us32\/_0736_ ), .B1(\us32\/_0022_ ), .B2(\us32\/_0099_ ), .X(\us32\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us32/_1049_ ( .A(\us32\/_0239_ ), .B(\us32\/_0240_ ), .C(\us32\/_0241_ ), .Y(\us32\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1050_ ( .A(\us32\/_0554_ ), .B(\us32\/_0072_ ), .X(\us32\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us32/_1051_ ( .A1(\us32\/_0142_ ), .A2(\us32\/_0137_ ), .B1(\us32\/_0159_ ), .B2(\us32\/_0082_ ), .X(\us32\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1052_ ( .A1(\us32\/_0608_ ), .A2(\us32\/_0072_ ), .B1(\us32\/_0243_ ), .C1(\us32\/_0244_ ), .Y(\us32\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1053_ ( .A(\us32\/_0234_ ), .B(\us32\/_0237_ ), .C(\us32\/_0242_ ), .D(\us32\/_0245_ ), .X(\us32\/_0246_ ) );
sky130_fd_sc_hd__buf_2 \us32/_1054_ ( .A(\us32\/_0027_ ), .X(\us32\/_0247_ ) );
sky130_fd_sc_hd__o21a_1 \us32/_1055_ ( .A1(\us32\/_0554_ ), .A2(\us32\/_0586_ ), .B1(\us32\/_0247_ ), .X(\us32\/_0248_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1056_ ( .A(\us32\/_0082_ ), .B(\us32\/_0478_ ), .X(\us32\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_1057_ ( .A(\us32\/_0079_ ), .X(\us32\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1058_ ( .A(\us32\/_0251_ ), .B(\us32\/_0478_ ), .X(\us32\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_1059_ ( .A(\us32\/_0250_ ), .B(\us32\/_0252_ ), .Y(\us32\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1060_ ( .A(\us32\/_0016_ ), .B(\us32\/_0064_ ), .Y(\us32\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_1061_ ( .A(\us32\/_0304_ ), .X(\us32\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1062_ ( .A(\us32\/_0255_ ), .B(\us32\/_0640_ ), .Y(\us32\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us32/_1063_ ( .A_N(\us32\/_0248_ ), .B(\us32\/_0253_ ), .C(\us32\/_0254_ ), .D(\us32\/_0256_ ), .X(\us32\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1064_ ( .A(\us32\/_0099_ ), .B(\us32\/_0110_ ), .X(\us32\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us32/_1065_ ( .A1(\us32\/_0161_ ), .A2(\us32\/_0130_ ), .B1(\us32\/_0258_ ), .Y(\us32\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1066_ ( .A(\us32\/_0194_ ), .B(\sa32\[1\] ), .X(\us32\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1068_ ( .A(\us32\/_0261_ ), .B(\us32\/_0153_ ), .Y(\us32\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us32/_1069_ ( .A_N(\us32\/_0154_ ), .B(\us32\/_0259_ ), .C(\us32\/_0263_ ), .X(\us32\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1070_ ( .A(\us32\/_0246_ ), .B(\us32\/_0174_ ), .C(\us32\/_0257_ ), .D(\us32\/_0264_ ), .X(\us32\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us32/_1071_ ( .A1(\us32\/_0261_ ), .A2(\us32\/_0554_ ), .B1(\us32\/_0159_ ), .X(\us32\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1072_ ( .A(\us32\/_0746_ ), .B(\us32\/_0150_ ), .Y(\us32\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1073_ ( .A(\us32\/_0175_ ), .Y(\us32\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us32/_1074_ ( .A(\us32\/_0412_ ), .B(\us32\/_0123_ ), .C(\us32\/_0151_ ), .X(\us32\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1075_ ( .A(\us32\/_0268_ ), .B(\us32\/_0269_ ), .Y(\us32\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us32/_1076_ ( .A_N(\us32\/_0266_ ), .B(\us32\/_0267_ ), .C(\us32\/_0270_ ), .X(\us32\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1077_ ( .A(\us32\/_0554_ ), .B(\us32\/_0150_ ), .X(\us32\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1078_ ( .A(\us32\/_0273_ ), .Y(\us32\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1079_ ( .A1(\us32\/_0734_ ), .A2(\us32\/_0325_ ), .B1(\us32\/_0380_ ), .Y(\us32\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1080_ ( .A(\us32\/_0275_ ), .Y(\us32\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1081_ ( .A(\us32\/_0276_ ), .B(\us32\/_0153_ ), .Y(\us32\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us32/_1082_ ( .A(\us32\/_0272_ ), .B(\us32\/_0274_ ), .C(\us32\/_0277_ ), .X(\us32\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_1083_ ( .A(\us32\/_0035_ ), .X(\us32\/_0279_ ) );
sky130_fd_sc_hd__buf_2 \us32/_1084_ ( .A(\us32\/_0082_ ), .X(\us32\/_0280_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1085_ ( .A1(\us32\/_0499_ ), .A2(\us32\/_0279_ ), .B1(\us32\/_0280_ ), .B2(\us32\/_0060_ ), .Y(\us32\/_0281_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1086_ ( .A1(\us32\/_0251_ ), .A2(\us32\/_0434_ ), .B1(\us32\/_0304_ ), .Y(\us32\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1087_ ( .A(\us32\/_0091_ ), .B(\us32\/_0056_ ), .Y(\us32\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1088_ ( .A1(\us32\/_0118_ ), .A2(\us32\/_0050_ ), .B1(\us32\/_0038_ ), .C1(\us32\/_0255_ ), .Y(\us32\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1089_ ( .A(\us32\/_0281_ ), .B(\us32\/_0283_ ), .C(\us32\/_0284_ ), .D(\us32\/_0285_ ), .X(\us32\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1090_ ( .A(\us32\/_0082_ ), .B(\us32\/_0027_ ), .X(\us32\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1091_ ( .A(\us32\/_0129_ ), .B(\us32\/_0027_ ), .X(\us32\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_1092_ ( .A(\us32\/_0287_ ), .B(\us32\/_0288_ ), .Y(\us32\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1093_ ( .A1(\us32\/_0752_ ), .A2(\us32\/_0683_ ), .B1(\us32\/_0093_ ), .B2(\us32\/_0247_ ), .Y(\us32\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1094_ ( .A1(\us32\/_0092_ ), .A2(\us32\/_0575_ ), .B1(\us32\/_0056_ ), .Y(\us32\/_0291_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1096_ ( .A1(\us32\/_0499_ ), .A2(\us32\/_0662_ ), .B1(\us32\/_0280_ ), .B2(\us32\/_0056_ ), .Y(\us32\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1097_ ( .A(\us32\/_0289_ ), .B(\us32\/_0290_ ), .C(\us32\/_0291_ ), .D(\us32\/_0294_ ), .X(\us32\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1098_ ( .A(\us32\/_0750_ ), .B(\us32\/_0193_ ), .X(\us32\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1099_ ( .A(\us32\/_0705_ ), .B(\us32\/_0380_ ), .X(\us32\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1100_ ( .A(\us32\/_0752_ ), .B(\us32\/_0129_ ), .Y(\us32\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us32/_1101_ ( .A(\us32\/_0296_ ), .B(\us32\/_0297_ ), .C_N(\us32\/_0298_ ), .Y(\us32\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1102_ ( .A(\us32\/_0089_ ), .B(\us32\/_0532_ ), .Y(\us32\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1103_ ( .A(\sa32\[2\] ), .Y(\us32\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \us32/_1104_ ( .A(\us32\/_0301_ ), .B(\sa32\[3\] ), .C(\us32\/_0118_ ), .Y(\us32\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1105_ ( .A(\us32\/_0072_ ), .B(\us32\/_0302_ ), .X(\us32\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1106_ ( .A(\us32\/_0303_ ), .Y(\us32\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1107_ ( .A(\us32\/_0147_ ), .B(\us32\/_0302_ ), .Y(\us32\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1108_ ( .A(\us32\/_0299_ ), .B(\us32\/_0300_ ), .C(\us32\/_0305_ ), .D(\us32\/_0306_ ), .X(\us32\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1109_ ( .A(\us32\/_0278_ ), .B(\us32\/_0286_ ), .C(\us32\/_0295_ ), .D(\us32\/_0307_ ), .X(\us32\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us32/_1110_ ( .A(\us32\/_0228_ ), .B(\us32\/_0265_ ), .C(\us32\/_0308_ ), .Y(\us32\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1111_ ( .A(\us32\/_0235_ ), .Y(\us32\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1112_ ( .A(\us32\/_0478_ ), .B(\us32\/_0640_ ), .X(\us32\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1113_ ( .A(\us32\/_0310_ ), .Y(\us32\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1114_ ( .A(\us32\/_0022_ ), .B(\us32\/_0499_ ), .Y(\us32\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1115_ ( .A(\us32\/_0499_ ), .B(\us32\/_0032_ ), .Y(\us32\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1116_ ( .A(\us32\/_0309_ ), .B(\us32\/_0311_ ), .C(\us32\/_0312_ ), .D(\us32\/_0313_ ), .X(\us32\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1117_ ( .A(\us32\/_0499_ ), .B(\us32\/_0064_ ), .Y(\us32\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1118_ ( .A(\us32\/_0499_ ), .B(\us32\/_0683_ ), .Y(\us32\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1119_ ( .A(\us32\/_0315_ ), .B(\us32\/_0316_ ), .C(\us32\/_0317_ ), .D(\us32\/_0253_ ), .X(\us32\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1120_ ( .A(\us32\/_0047_ ), .B(\us32\/_0304_ ), .Y(\us32\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1121_ ( .A(\us32\/_0586_ ), .B(\us32\/_0162_ ), .Y(\us32\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1122_ ( .A(\us32\/_0319_ ), .B(\us32\/_0320_ ), .Y(\us32\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_1123_ ( .A(\us32\/_0321_ ), .B(\us32\/_0238_ ), .Y(\us32\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1124_ ( .A(\us32\/_0304_ ), .B(\us32\/_0062_ ), .Y(\us32\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_1125_ ( .A(\us32\/_0251_ ), .X(\us32\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1126_ ( .A1(\us32\/_0324_ ), .A2(\us32\/_0280_ ), .B1(\us32\/_0255_ ), .Y(\us32\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1127_ ( .A1(\us32\/_0050_ ), .A2(\us32\/_0205_ ), .B1(\us32\/_0109_ ), .C1(\us32\/_0255_ ), .Y(\us32\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1128_ ( .A(\us32\/_0322_ ), .B(\us32\/_0323_ ), .C(\us32\/_0326_ ), .D(\us32\/_0327_ ), .X(\us32\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1129_ ( .A1(\us32\/_0733_ ), .A2(\us32\/_0279_ ), .A3(\us32\/_0058_ ), .B1(\us32\/_0056_ ), .Y(\us32\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_1130_ ( .A(\us32\/_0047_ ), .X(\us32\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1131_ ( .A(\us32\/_0330_ ), .B(\us32\/_0056_ ), .Y(\us32\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1132_ ( .A(\us32\/_0054_ ), .B(\us32\/_0045_ ), .Y(\us32\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1133_ ( .A(\us32\/_0329_ ), .B(\us32\/_0331_ ), .C(\us32\/_0284_ ), .D(\us32\/_0332_ ), .X(\us32\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us32/_1134_ ( .A1(\us32\/_0249_ ), .A2(\us32\/_0205_ ), .B1(\us32\/_0532_ ), .C1(\us32\/_0060_ ), .X(\us32\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1135_ ( .A(\us32\/_0280_ ), .B(\us32\/_0060_ ), .Y(\us32\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1136_ ( .A(\us32\/_0324_ ), .B(\us32\/_0060_ ), .Y(\us32\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1137_ ( .A(\us32\/_0335_ ), .B(\us32\/_0337_ ), .Y(\us32\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1138_ ( .A1(\us32\/_0276_ ), .A2(\us32\/_0060_ ), .B1(\us32\/_0334_ ), .C1(\us32\/_0338_ ), .Y(\us32\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1139_ ( .A(\us32\/_0318_ ), .B(\us32\/_0328_ ), .C(\us32\/_0333_ ), .D(\us32\/_0339_ ), .X(\us32\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us32/_1140_ ( .A1(\us32\/_0746_ ), .A2(\us32\/_0134_ ), .B1(\us32\/_0128_ ), .X(\us32\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us32/_1141_ ( .A_N(\us32\/_0086_ ), .B(\us32\/_0128_ ), .X(\us32\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1142_ ( .A(\us32\/_0079_ ), .B(\us32\/_0124_ ), .X(\us32\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_1143_ ( .A(\us32\/_0126_ ), .B(\us32\/_0343_ ), .Y(\us32\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us32/_1144_ ( .A(\us32\/_0341_ ), .B(\us32\/_0342_ ), .C_N(\us32\/_0344_ ), .Y(\us32\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1146_ ( .A1(\us32\/_0193_ ), .A2(\us32\/_0092_ ), .A3(\us32\/_0330_ ), .B1(\us32\/_0147_ ), .Y(\us32\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1147_ ( .A1(\us32\/_0130_ ), .A2(\us32\/_0280_ ), .A3(\us32\/_0134_ ), .B1(\us32\/_0139_ ), .Y(\us32\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1148_ ( .A1(\us32\/_0144_ ), .A2(\us32\/_0608_ ), .A3(\us32\/_0092_ ), .B1(\us32\/_0139_ ), .Y(\us32\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1149_ ( .A(\us32\/_0345_ ), .B(\us32\/_0348_ ), .C(\us32\/_0349_ ), .D(\us32\/_0350_ ), .X(\us32\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us32/_1150_ ( .A(\us32\/_0150_ ), .B(\us32\/_0194_ ), .C(\us32\/_0249_ ), .X(\us32\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us32/_1151_ ( .A(\us32\/_0277_ ), .SLEEP(\us32\/_0352_ ), .X(\us32\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us32/_1152_ ( .A1(\us32\/_0268_ ), .A2(\us32\/_0171_ ), .B1(\us32\/_0157_ ), .Y(\us32\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us32/_1153_ ( .A(\us32\/_0161_ ), .X(\us32\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1154_ ( .A1(\us32\/_0279_ ), .A2(\us32\/_0280_ ), .B1(\us32\/_0355_ ), .Y(\us32\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1155_ ( .A1(\us32\/_0020_ ), .A2(\us32\/_0193_ ), .A3(\us32\/_0091_ ), .B1(\us32\/_0355_ ), .Y(\us32\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1156_ ( .A(\us32\/_0353_ ), .B(\us32\/_0354_ ), .C(\us32\/_0356_ ), .D(\us32\/_0357_ ), .X(\us32\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1157_ ( .A(\us32\/_0111_ ), .B(\us32\/_0586_ ), .X(\us32\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1158_ ( .A(\us32\/_0360_ ), .Y(\us32\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us32/_1159_ ( .A1(\us32\/_0119_ ), .A2(\us32\/_0120_ ), .B1(\us32\/_0230_ ), .C1(\us32\/_0361_ ), .X(\us32\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1160_ ( .A1(\us32\/_0662_ ), .A2(\us32\/_0251_ ), .A3(\us32\/_0134_ ), .B1(\us32\/_0114_ ), .Y(\us32\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1162_ ( .A1(\us32\/_0035_ ), .A2(\us32\/_0251_ ), .A3(\us32\/_0134_ ), .B1(\us32\/_0099_ ), .Y(\us32\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1163_ ( .A1(\us32\/_0193_ ), .A2(\us32\/_0608_ ), .B1(\us32\/_0099_ ), .Y(\us32\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1164_ ( .A(\us32\/_0362_ ), .B(\us32\/_0363_ ), .C(\us32\/_0365_ ), .D(\us32\/_0366_ ), .X(\us32\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1165_ ( .A1(\us32\/_0575_ ), .A2(\us32\/_0092_ ), .A3(\us32\/_0330_ ), .B1(\us32\/_0089_ ), .Y(\us32\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1166_ ( .A1(\us32\/_0586_ ), .A2(\us32\/_0017_ ), .A3(\us32\/_0330_ ), .B1(\us32\/_0094_ ), .Y(\us32\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \us32/_1167_ ( .A1(\us32\/_0293_ ), .A2(\us32\/_0134_ ), .B1(\us32\/_0089_ ), .Y(\us32\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1168_ ( .A1(\us32\/_0279_ ), .A2(\us32\/_0134_ ), .B1(\us32\/_0094_ ), .Y(\us32\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1169_ ( .A(\us32\/_0368_ ), .B(\us32\/_0370_ ), .C(\us32\/_0371_ ), .D(\us32\/_0372_ ), .X(\us32\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1170_ ( .A(\us32\/_0351_ ), .B(\us32\/_0359_ ), .C(\us32\/_0367_ ), .D(\us32\/_0373_ ), .X(\us32\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1171_ ( .A1(\us32\/_0102_ ), .A2(\us32\/_0347_ ), .B1(\us32\/_0109_ ), .C1(\us32\/_0247_ ), .Y(\us32\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1172_ ( .A1(\us32\/_0102_ ), .A2(\us32\/_0347_ ), .B1(\us32\/_0532_ ), .C1(\us32\/_0247_ ), .Y(\us32\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1173_ ( .A1(\us32\/_0050_ ), .A2(\us32\/_0249_ ), .B1(\us32\/_0380_ ), .C1(\us32\/_0247_ ), .Y(\us32\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1174_ ( .A(\us32\/_0041_ ), .B(\us32\/_0375_ ), .C(\us32\/_0376_ ), .D(\us32\/_0377_ ), .X(\us32\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1175_ ( .A(\us32\/_0047_ ), .B(\us32\/_0750_ ), .X(\us32\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1176_ ( .A(\us32\/_0379_ ), .Y(\us32\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1177_ ( .A(\us32\/_0016_ ), .B(\us32\/_0608_ ), .Y(\us32\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1178_ ( .A(\us32\/_0752_ ), .B(\us32\/_0554_ ), .Y(\us32\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1179_ ( .A1(\sa32\[1\] ), .A2(\us32\/_0734_ ), .B1(\us32\/_0109_ ), .C1(\us32\/_0016_ ), .Y(\us32\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1180_ ( .A(\us32\/_0381_ ), .B(\us32\/_0382_ ), .C(\us32\/_0383_ ), .D(\us32\/_0384_ ), .X(\us32\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us32/_1181_ ( .A(\us32\/_0086_ ), .B_N(\us32\/_0736_ ), .X(\us32\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1182_ ( .A1(\us32\/_0748_ ), .A2(\us32\/_0134_ ), .B1(\us32\/_0739_ ), .Y(\us32\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1183_ ( .A1(\us32\/_0118_ ), .A2(\us32\/_0249_ ), .B1(\us32\/_0109_ ), .C1(\us32\/_0739_ ), .Y(\us32\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1184_ ( .A1(\us32\/_0102_ ), .A2(\us32\/_0301_ ), .B1(\sa32\[3\] ), .C1(\us32\/_0739_ ), .Y(\us32\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1185_ ( .A(\us32\/_0386_ ), .B(\us32\/_0387_ ), .C(\us32\/_0388_ ), .D(\us32\/_0389_ ), .X(\us32\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1186_ ( .A(\us32\/_0020_ ), .Y(\us32\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1187_ ( .A(\us32\/_0727_ ), .Y(\us32\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1188_ ( .A(\us32\/_0727_ ), .B(\us32\/_0064_ ), .Y(\us32\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1189_ ( .A1(\us32\/_0102_ ), .A2(\us32\/_0734_ ), .B1(\us32\/_0532_ ), .C1(\us32\/_0727_ ), .Y(\us32\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us32/_1190_ ( .A1(\us32\/_0392_ ), .A2(\us32\/_0393_ ), .B1(\us32\/_0394_ ), .C1(\us32\/_0395_ ), .X(\us32\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1191_ ( .A(\us32\/_0378_ ), .B(\us32\/_0385_ ), .C(\us32\/_0390_ ), .D(\us32\/_0396_ ), .X(\us32\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us32/_1192_ ( .A(\us32\/_0340_ ), .B(\us32\/_0374_ ), .C(\us32\/_0397_ ), .Y(\us32\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1193_ ( .A(\us32\/_0077_ ), .B(\us32\/_0129_ ), .X(\us32\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_1194_ ( .A(\us32\/_0398_ ), .B(\us32\/_0239_ ), .Y(\us32\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1195_ ( .A(\us32\/_0022_ ), .B(\us32\/_0111_ ), .X(\us32\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us32/_1196_ ( .A_N(\us32\/_0400_ ), .B(\us32\/_0231_ ), .Y(\us32\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us32/_1197_ ( .A(\us32\/_0399_ ), .SLEEP(\us32\/_0402_ ), .X(\us32\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_1198_ ( .A(\us32\/_0746_ ), .B(\us32\/_0251_ ), .Y(\us32\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us32/_1199_ ( .A_N(\us32\/_0404_ ), .B(\us32\/_0752_ ), .Y(\us32\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us32/_1200_ ( .A(\us32\/_0467_ ), .B(\us32\/_0194_ ), .C(\us32\/_0694_ ), .X(\us32\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us32/_1201_ ( .A_N(\us32\/_0175_ ), .B(\us32\/_0406_ ), .X(\us32\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1202_ ( .A(\us32\/_0407_ ), .Y(\us32\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1203_ ( .A1(\us32\/_0094_ ), .A2(\us32\/_0197_ ), .B1(\us32\/_0114_ ), .B2(\us32\/_0640_ ), .Y(\us32\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1204_ ( .A(\us32\/_0403_ ), .B(\us32\/_0405_ ), .C(\us32\/_0408_ ), .D(\us32\/_0409_ ), .X(\us32\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1205_ ( .A(\us32\/_0030_ ), .B(\us32\/_0150_ ), .Y(\us32\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us32/_1206_ ( .A_N(\us32\/_0169_ ), .B(\us32\/_0289_ ), .C(\us32\/_0411_ ), .X(\us32\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us32/_1207_ ( .A1(\us32\/_0467_ ), .A2(\us32\/_0151_ ), .B1(\us32\/_0140_ ), .C1(\us32\/_0129_ ), .X(\us32\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1208_ ( .A1(\us32\/_0608_ ), .A2(\us32\/_0099_ ), .B1(\us32\/_0037_ ), .C1(\us32\/_0414_ ), .Y(\us32\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1209_ ( .A(\us32\/_0738_ ), .Y(\us32\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1210_ ( .A(\us32\/_0586_ ), .B(\us32\/_0736_ ), .Y(\us32\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1211_ ( .A1(\us32\/_0194_ ), .A2(\us32\/_0038_ ), .B1(\us32\/_0118_ ), .C1(\us32\/_0153_ ), .Y(\us32\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us32/_1212_ ( .A1(\us32\/_0416_ ), .A2(\us32\/_0117_ ), .B1(\us32\/_0417_ ), .C1(\us32\/_0418_ ), .X(\us32\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1213_ ( .A(\us32\/_0077_ ), .B(\us32\/_0035_ ), .X(\us32\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1214_ ( .A(\us32\/_0662_ ), .B(\us32\/_0124_ ), .Y(\us32\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1215_ ( .A(\us32\/_0030_ ), .B(\us32\/_0137_ ), .Y(\us32\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1216_ ( .A(\us32\/_0072_ ), .B(\us32\/_0731_ ), .Y(\us32\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us32/_1217_ ( .A_N(\us32\/_0420_ ), .B(\us32\/_0421_ ), .C(\us32\/_0422_ ), .D(\us32\/_0424_ ), .X(\us32\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1218_ ( .A(\us32\/_0413_ ), .B(\us32\/_0415_ ), .C(\us32\/_0419_ ), .D(\us32\/_0425_ ), .X(\us32\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us32/_1219_ ( .A(\us32\/_0355_ ), .B(\us32\/_0102_ ), .C(\us32\/_0109_ ), .Y(\us32\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1220_ ( .A(\us32\/_0077_ ), .B(\us32\/_0017_ ), .X(\us32\/_0428_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1221_ ( .A(\us32\/_0077_ ), .B(\us32\/_0554_ ), .X(\us32\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us32/_1222_ ( .A1(\us32\/_0050_ ), .A2(\us32\/_0205_ ), .B1(\us32\/_0380_ ), .C1(\us32\/_0078_ ), .X(\us32\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us32/_1223_ ( .A(\us32\/_0428_ ), .B(\us32\/_0429_ ), .C(\us32\/_0430_ ), .Y(\us32\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us32/_1224_ ( .A_N(\us32\/_0209_ ), .B(\us32\/_0431_ ), .X(\us32\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us32/_1225_ ( .A1(\us32\/_0215_ ), .A2(\us32\/_0404_ ), .B1(\us32\/_0427_ ), .C1(\us32\/_0432_ ), .X(\us32\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1226_ ( .A(\us32\/_0043_ ), .B(\us32\/_0058_ ), .Y(\us32\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1227_ ( .A(\us32\/_0195_ ), .B(\us32\/_0233_ ), .C(\us32\/_0320_ ), .D(\us32\/_0435_ ), .X(\us32\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1228_ ( .A(\us32\/_0261_ ), .B(\us32\/_0738_ ), .Y(\us32\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1229_ ( .A1(\us32\/_0499_ ), .A2(\us32\/_0640_ ), .B1(\us32\/_0261_ ), .B2(\us32\/_0056_ ), .Y(\us32\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1230_ ( .A(\us32\/_0436_ ), .B(\us32\/_0394_ ), .C(\us32\/_0437_ ), .D(\us32\/_0438_ ), .X(\us32\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1231_ ( .A(\us32\/_0410_ ), .B(\us32\/_0426_ ), .C(\us32\/_0433_ ), .D(\us32\/_0439_ ), .X(\us32\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us32/_1232_ ( .A(\us32\/_0135_ ), .SLEEP(\us32\/_0273_ ), .X(\us32\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1233_ ( .A1(\us32\/_0279_ ), .A2(\us32\/_0134_ ), .B1(\us32\/_0099_ ), .Y(\us32\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1234_ ( .A(\us32\/_0441_ ), .B(\us32\/_0164_ ), .C(\us32\/_0270_ ), .D(\us32\/_0442_ ), .X(\us32\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1235_ ( .A(\us32\/_0051_ ), .B(\us32\/_0662_ ), .Y(\us32\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1236_ ( .A(\us32\/_0051_ ), .B(\us32\/_0271_ ), .Y(\us32\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1237_ ( .A(\us32\/_0444_ ), .B(\us32\/_0446_ ), .X(\us32\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1238_ ( .A(\us32\/_0193_ ), .B(\us32\/_0304_ ), .X(\us32\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1239_ ( .A(\us32\/_0448_ ), .Y(\us32\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1240_ ( .A(\us32\/_0162_ ), .B(\us32\/_0130_ ), .X(\us32\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1241_ ( .A(\us32\/_0450_ ), .Y(\us32\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1242_ ( .A1(\us32\/_0129_ ), .A2(\us32\/_0554_ ), .B1(\us32\/_0043_ ), .Y(\us32\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1243_ ( .A(\us32\/_0447_ ), .B(\us32\/_0449_ ), .C(\us32\/_0451_ ), .D(\us32\/_0452_ ), .X(\us32\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1244_ ( .A(\us32\/_0056_ ), .B(\us32\/_0064_ ), .Y(\us32\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us32/_1245_ ( .A_N(\us32\/_0248_ ), .B(\us32\/_0454_ ), .C(\us32\/_0254_ ), .D(\us32\/_0256_ ), .X(\us32\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1246_ ( .A1(\us32\/_0330_ ), .A2(\us32\/_0099_ ), .B1(\us32\/_0134_ ), .B2(\us32\/_0705_ ), .Y(\us32\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1247_ ( .A1(\us32\/_0748_ ), .A2(\us32\/_0738_ ), .B1(\us32\/_0092_ ), .B2(\us32\/_0752_ ), .Y(\us32\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1248_ ( .A1(\us32\/_0072_ ), .A2(\us32\/_0035_ ), .B1(\us32\/_0748_ ), .B2(\us32\/_0056_ ), .Y(\us32\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1249_ ( .A1(\us32\/_0748_ ), .A2(\us32\/_0251_ ), .B1(\us32\/_0247_ ), .Y(\us32\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1250_ ( .A(\us32\/_0457_ ), .B(\us32\/_0458_ ), .C(\us32\/_0459_ ), .D(\us32\/_0460_ ), .X(\us32\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1251_ ( .A(\us32\/_0443_ ), .B(\us32\/_0453_ ), .C(\us32\/_0455_ ), .D(\us32\/_0461_ ), .X(\us32\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1252_ ( .A(\us32\/_0705_ ), .B(\us32\/_0079_ ), .X(\us32\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1253_ ( .A(\us32\/_0586_ ), .B(\us32\/_0124_ ), .Y(\us32\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1254_ ( .A(\us32\/_0499_ ), .B(\us32\/_0746_ ), .Y(\us32\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us32/_1255_ ( .A_N(\us32\/_0463_ ), .B(\us32\/_0464_ ), .C(\us32\/_0465_ ), .X(\us32\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us32/_1256_ ( .A1(\us32\/_0271_ ), .A2(\us32\/_0072_ ), .B1(\us32\/_0142_ ), .B2(\us32\/_0027_ ), .X(\us32\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1257_ ( .A1(\us32\/_0144_ ), .A2(\us32\/_0099_ ), .B1(\us32\/_0360_ ), .C1(\us32\/_0468_ ), .Y(\us32\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us32/_1258_ ( .A1(\us32\/_0662_ ), .A2(\us32\/_0251_ ), .B1(\us32\/_0499_ ), .X(\us32\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1259_ ( .A1(\us32\/_0575_ ), .A2(\us32\/_0056_ ), .B1(\us32\/_0379_ ), .C1(\us32\/_0470_ ), .Y(\us32\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1260_ ( .A(\us32\/_0466_ ), .B(\us32\/_0469_ ), .C(\us32\/_0471_ ), .D(\us32\/_0305_ ), .X(\us32\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us32/_1261_ ( .A1(\us32\/_0247_ ), .A2(\us32\/_0683_ ), .B1(\us32\/_0324_ ), .B2(\us32\/_0056_ ), .X(\us32\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1262_ ( .A(\us32\/_0280_ ), .B(\us32\/_0099_ ), .X(\us32\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us32/_1263_ ( .A1(\us32\/_0092_ ), .A2(\us32\/_0247_ ), .B1(\us32\/_0474_ ), .X(\us32\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us32/_1264_ ( .A(\us32\/_0075_ ), .B(\us32\/_0473_ ), .C(\us32\/_0475_ ), .Y(\us32\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1265_ ( .A1(\us32\/_0279_ ), .A2(\us32\/_0255_ ), .B1(\us32\/_0280_ ), .B2(\us32\/_0060_ ), .Y(\us32\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1266_ ( .A1(\us32\/_0093_ ), .A2(\us32\/_0056_ ), .B1(\us32\/_0134_ ), .B2(\us32\/_0114_ ), .Y(\us32\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1267_ ( .A1(\us32\/_0161_ ), .A2(\us32\/_0032_ ), .B1(\us32\/_0324_ ), .B2(\us32\/_0147_ ), .Y(\us32\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1268_ ( .A1(\us32\/_0054_ ), .A2(\us32\/_0731_ ), .B1(\us32\/_0748_ ), .B2(\us32\/_0304_ ), .Y(\us32\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1269_ ( .A(\us32\/_0477_ ), .B(\us32\/_0479_ ), .C(\us32\/_0480_ ), .D(\us32\/_0481_ ), .X(\us32\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1270_ ( .A(\us32\/_0161_ ), .B(\us32\/_0064_ ), .Y(\us32\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us32/_1271_ ( .A(\us32\/_0731_ ), .B(\us32\/_0123_ ), .C(\us32\/_0467_ ), .Y(\us32\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1272_ ( .A(\us32\/_0483_ ), .B(\us32\/_0484_ ), .Y(\us32\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1273_ ( .A(\us32\/_0297_ ), .Y(\us32\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us32/_1274_ ( .A_N(\us32\/_0485_ ), .B(\us32\/_0181_ ), .C(\us32\/_0486_ ), .D(\us32\/_0386_ ), .X(\us32\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1275_ ( .A(\us32\/_0472_ ), .B(\us32\/_0476_ ), .C(\us32\/_0482_ ), .D(\us32\/_0487_ ), .X(\us32\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \us32/_1276_ ( .A(\us32\/_0440_ ), .B(\us32\/_0462_ ), .C(\us32\/_0488_ ), .Y(\us32\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1277_ ( .A(\us32\/_0403_ ), .B(\us32\/_0230_ ), .C(\us32\/_0451_ ), .D(\us32\/_0361_ ), .X(\us32\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1278_ ( .A1(\us32\/_0118_ ), .A2(\us32\/_0050_ ), .B1(\us32\/_0109_ ), .C1(\us32\/_0139_ ), .Y(\us32\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1279_ ( .A(\us32\/_0447_ ), .B(\us32\/_0437_ ), .C(\us32\/_0491_ ), .D(\us32\/_0427_ ), .X(\us32\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1280_ ( .A1(\us32\/_0280_ ), .A2(\us32\/_0255_ ), .B1(\us32\/_0608_ ), .B2(\us32\/_0247_ ), .Y(\us32\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1281_ ( .A1(\us32\/_0144_ ), .A2(\us32\/_0147_ ), .B1(\us32\/_0355_ ), .B2(\us32\/_0093_ ), .Y(\us32\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1282_ ( .A1(\us32\/_0705_ ), .A2(\us32\/_0279_ ), .B1(\us32\/_0330_ ), .B2(\us32\/_0247_ ), .Y(\us32\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1283_ ( .A1(\us32\/_0279_ ), .A2(\us32\/_0280_ ), .B1(\us32\/_0114_ ), .Y(\us32\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1284_ ( .A(\us32\/_0493_ ), .B(\us32\/_0494_ ), .C(\us32\/_0495_ ), .D(\us32\/_0496_ ), .X(\us32\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1285_ ( .A1(\us32\/_0134_ ), .A2(\us32\/_0137_ ), .B1(\us32\/_0355_ ), .B2(\us32\/_0575_ ), .Y(\us32\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1286_ ( .A1(\us32\/_0099_ ), .A2(\us32\/_0733_ ), .B1(\us32\/_0093_ ), .B2(\us32\/_0499_ ), .Y(\us32\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1287_ ( .A(\us32\/_0147_ ), .B(\us32\/_0640_ ), .Y(\us32\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1288_ ( .A1(\us32\/_0153_ ), .A2(\us32\/_0056_ ), .B1(\us32\/_0748_ ), .Y(\us32\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1289_ ( .A(\us32\/_0498_ ), .B(\us32\/_0500_ ), .C(\us32\/_0501_ ), .D(\us32\/_0502_ ), .X(\us32\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1290_ ( .A(\us32\/_0490_ ), .B(\us32\/_0492_ ), .C(\us32\/_0497_ ), .D(\us32\/_0503_ ), .X(\us32\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us32/_1291_ ( .A_N(\us32\/_0275_ ), .B(\us32\/_0705_ ), .X(\us32\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1292_ ( .A(\us32\/_0505_ ), .Y(\us32\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1293_ ( .A(\us32\/_0380_ ), .B(\us32\/_0347_ ), .X(\us32\/_0507_ ) );
sky130_fd_sc_hd__o21ai_1 \us32/_1294_ ( .A1(\us32\/_0507_ ), .A2(\us32\/_0093_ ), .B1(\us32\/_0056_ ), .Y(\us32\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1295_ ( .A(\us32\/_0322_ ), .B(\us32\/_0277_ ), .C(\us32\/_0506_ ), .D(\us32\/_0508_ ), .X(\us32\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1296_ ( .A(\us32\/_0280_ ), .B(\us32\/_0705_ ), .X(\us32\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1297_ ( .A1(\us32\/_0733_ ), .A2(\us32\/_0114_ ), .B1(\us32\/_0429_ ), .C1(\us32\/_0511_ ), .Y(\us32\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_1298_ ( .A(\us32\/_0019_ ), .B(\us32\/_0024_ ), .Y(\us32\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1299_ ( .A(\us32\/_0512_ ), .B(\us32\/_0513_ ), .C(\us32\/_0742_ ), .D(\us32\/_0306_ ), .X(\us32\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1300_ ( .A1(\us32\/_0532_ ), .A2(\us32\/_0089_ ), .B1(\us32\/_0154_ ), .C1(\us32\/_0169_ ), .Y(\us32\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us32/_1301_ ( .A1(\us32\/_0749_ ), .A2(\us32\/_0026_ ), .B1(\us32\/_0069_ ), .C1(\us32\/_0032_ ), .X(\us32\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us32/_1302_ ( .A1(\us32\/_0324_ ), .A2(\us32\/_0355_ ), .B1(\us32\/_0330_ ), .B2(\us32\/_0727_ ), .X(\us32\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us32/_1303_ ( .A(\us32\/_0133_ ), .B(\us32\/_0516_ ), .C(\us32\/_0517_ ), .Y(\us32\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1304_ ( .A(\us32\/_0509_ ), .B(\us32\/_0514_ ), .C(\us32\/_0515_ ), .D(\us32\/_0518_ ), .X(\us32\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1305_ ( .A(\us32\/_0746_ ), .B(\us32\/_0072_ ), .Y(\us32\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1306_ ( .A1(\us32\/_0082_ ), .A2(\us32\/_0070_ ), .B1(\us32\/_0043_ ), .B2(\us32\/_0193_ ), .Y(\us32\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1307_ ( .A(\us32\/_0311_ ), .B(\us32\/_0520_ ), .C(\us32\/_0332_ ), .D(\us32\/_0522_ ), .X(\us32\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1308_ ( .A(\us32\/_0129_ ), .B(\us32\/_0499_ ), .X(\us32\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_1309_ ( .A(\us32\/_0235_ ), .B(\us32\/_0524_ ), .Y(\us32\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us32/_1310_ ( .A(\us32\/_0081_ ), .B(\us32\/_0085_ ), .Y(\us32\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1311_ ( .A1(\us32\/_0051_ ), .A2(\us32\/_0045_ ), .B1(\us32\/_0130_ ), .B2(\us32\/_0094_ ), .Y(\us32\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1312_ ( .A(\us32\/_0523_ ), .B(\us32\/_0525_ ), .C(\us32\/_0526_ ), .D(\us32\/_0527_ ), .X(\us32\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us32/_1313_ ( .A_N(\us32\/_0250_ ), .B(\us32\/_0521_ ), .Y(\us32\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1314_ ( .A(\us32\/_0128_ ), .B(\us32\/_0020_ ), .X(\us32\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1315_ ( .A(\us32\/_0530_ ), .Y(\us32\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1316_ ( .A(\us32\/_0099_ ), .B(\us32\/_0058_ ), .X(\us32\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1317_ ( .A(\us32\/_0533_ ), .Y(\us32\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us32/_1318_ ( .A_N(\us32\/_0529_ ), .B(\us32\/_0531_ ), .C(\us32\/_0534_ ), .D(\us32\/_0192_ ), .X(\us32\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1319_ ( .A(\us32\/_0434_ ), .B(\us32\/_0078_ ), .X(\us32\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us32/_1320_ ( .A1(\us32\/_0750_ ), .A2(\us32\/_0079_ ), .B1(\us32\/_0129_ ), .B2(\us32\/_0705_ ), .X(\us32\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1321_ ( .A1(\us32\/_0161_ ), .A2(\us32\/_0032_ ), .B1(\us32\/_0536_ ), .C1(\us32\/_0537_ ), .Y(\us32\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us32/_1322_ ( .A1(\us32\/_0746_ ), .A2(\us32\/_0162_ ), .B1(\us32\/_0079_ ), .B2(\us32\/_0043_ ), .X(\us32\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1323_ ( .A1(\us32\/_0093_ ), .A2(\us32\/_0247_ ), .B1(\us32\/_0240_ ), .C1(\us32\/_0539_ ), .Y(\us32\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1324_ ( .A(\us32\/_0434_ ), .B(\us32\/_0043_ ), .X(\us32\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us32/_1325_ ( .A1(\us32\/_0142_ ), .A2(\us32\/_0150_ ), .B1(\us32\/_0022_ ), .B2(\us32\/_0137_ ), .X(\us32\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1326_ ( .A1(\us32\/_0279_ ), .A2(\us32\/_0051_ ), .B1(\us32\/_0541_ ), .C1(\us32\/_0542_ ), .Y(\us32\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1327_ ( .A(\us32\/_0159_ ), .B(\us32\/_0035_ ), .X(\us32\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us32/_1328_ ( .A1(\us32\/_0271_ ), .A2(\us32\/_0434_ ), .B1(\us32\/_0027_ ), .X(\us32\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1329_ ( .A1(\us32\/_0091_ ), .A2(\us32\/_0128_ ), .B1(\us32\/_0545_ ), .C1(\us32\/_0546_ ), .Y(\us32\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1330_ ( .A(\us32\/_0538_ ), .B(\us32\/_0540_ ), .C(\us32\/_0544_ ), .D(\us32\/_0547_ ), .X(\us32\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1331_ ( .A(\us32\/_0099_ ), .B(\us32\/_0193_ ), .X(\us32\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us32/_1332_ ( .A(\us32\/_0549_ ), .B(\us32\/_0186_ ), .C(\us32\/_0187_ ), .Y(\us32\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1333_ ( .A(\us32\/_0062_ ), .B(\us32\/_0347_ ), .C(\us32\/_0749_ ), .D(\us32\/_0694_ ), .X(\us32\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1334_ ( .A1(\us32\/_0130_ ), .A2(\us32\/_0499_ ), .B1(\us32\/_0551_ ), .C1(\us32\/_0101_ ), .Y(\us32\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1335_ ( .A(\us32\/_0139_ ), .B(\us32\/_0640_ ), .Y(\us32\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1336_ ( .A1(\us32\/_0752_ ), .A2(\us32\/_0662_ ), .B1(\us32\/_0280_ ), .B2(\us32\/_0099_ ), .Y(\us32\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1337_ ( .A(\us32\/_0550_ ), .B(\us32\/_0552_ ), .C(\us32\/_0553_ ), .D(\us32\/_0555_ ), .X(\us32\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1338_ ( .A(\us32\/_0528_ ), .B(\us32\/_0535_ ), .C(\us32\/_0548_ ), .D(\us32\/_0556_ ), .X(\us32\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us32/_1339_ ( .A(\us32\/_0504_ ), .B(\us32\/_0519_ ), .C(\us32\/_0557_ ), .Y(\us32\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1340_ ( .A(\us32\/_0054_ ), .B(\us32\/_0507_ ), .X(\us32\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us32/_1341_ ( .A_N(\us32\/_0558_ ), .B(\us32\/_0408_ ), .C(\us32\/_0451_ ), .D(\us32\/_0452_ ), .X(\us32\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1342_ ( .A(\us32\/_0549_ ), .Y(\us32\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1343_ ( .A(\us32\/_0559_ ), .B(\us32\/_0403_ ), .C(\us32\/_0560_ ), .D(\us32\/_0371_ ), .X(\us32\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1344_ ( .A(\us32\/_0181_ ), .B(\us32\/_0178_ ), .X(\us32\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1345_ ( .A(\us32\/_0562_ ), .B(\us32\/_0552_ ), .C(\us32\/_0553_ ), .D(\us32\/_0555_ ), .X(\us32\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1346_ ( .A(\us32\/_0247_ ), .B(\us32\/_0020_ ), .Y(\us32\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1347_ ( .A(\us32\/_0051_ ), .B(\us32\/_0130_ ), .X(\us32\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1348_ ( .A(\us32\/_0566_ ), .Y(\us32\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1349_ ( .A(\us32\/_0159_ ), .B(\us32\/_0412_ ), .X(\us32\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1350_ ( .A1(\us32\/_0752_ ), .A2(\us32\/_0640_ ), .B1(\us32\/_0568_ ), .B2(\us32\/_0175_ ), .Y(\us32\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1351_ ( .A(\us32\/_0076_ ), .B(\us32\/_0565_ ), .C(\us32\/_0567_ ), .D(\us32\/_0569_ ), .X(\us32\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us32/_1352_ ( .A1(\us32\/_0035_ ), .A2(\us32\/_0142_ ), .B1(\us32\/_0161_ ), .X(\us32\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1353_ ( .A(\us32\/_0099_ ), .B(\us32\/_0662_ ), .Y(\us32\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us32/_1354_ ( .A(\us32\/_0420_ ), .B(\us32\/_0571_ ), .C_N(\us32\/_0572_ ), .Y(\us32\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1355_ ( .A(\us32\/_0051_ ), .B(\us32\/_0746_ ), .Y(\us32\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1356_ ( .A(\us32\/_0574_ ), .B(\us32\/_0319_ ), .C(\us32\/_0320_ ), .D(\us32\/_0411_ ), .X(\us32\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1357_ ( .A(\us32\/_0736_ ), .B(\us32\/_0035_ ), .Y(\us32\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1358_ ( .A(\us32\/_0736_ ), .B(\us32\/_0030_ ), .Y(\us32\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1359_ ( .A(\us32\/_0298_ ), .B(\us32\/_0208_ ), .C(\us32\/_0577_ ), .D(\us32\/_0578_ ), .X(\us32\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1360_ ( .A1(\us32\/_0020_ ), .A2(\us32\/_0137_ ), .B1(\us32\/_0261_ ), .B2(\us32\/_0128_ ), .Y(\us32\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1361_ ( .A(\us32\/_0573_ ), .B(\us32\/_0576_ ), .C(\us32\/_0579_ ), .D(\us32\/_0580_ ), .X(\us32\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1362_ ( .A(\us32\/_0561_ ), .B(\us32\/_0563_ ), .C(\us32\/_0570_ ), .D(\us32\/_0581_ ), .X(\us32\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1363_ ( .A(\us32\/_0128_ ), .B(\us32\/_0193_ ), .X(\us32\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1364_ ( .A(\us32\/_0082_ ), .B(\us32\/_0162_ ), .X(\us32\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us32/_1365_ ( .A(\us32\/_0583_ ), .B(\us32\/_0584_ ), .C_N(\us32\/_0437_ ), .Y(\us32\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us32/_1366_ ( .A(\us32\/_0150_ ), .B(\us32\/_0118_ ), .C(\us32\/_0380_ ), .Y(\us32\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us32/_1367_ ( .A_N(\us32\/_0182_ ), .B(\us32\/_0587_ ), .C(\us32\/_0323_ ), .X(\us32\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1368_ ( .A1(\us32\/_0575_ ), .A2(\us32\/_0153_ ), .B1(\us32\/_0727_ ), .B2(\us32\/_0058_ ), .Y(\us32\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1369_ ( .A1(\us32\/_0499_ ), .A2(\us32\/_0064_ ), .B1(\us32\/_0134_ ), .B2(\us32\/_0255_ ), .Y(\us32\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1370_ ( .A(\us32\/_0585_ ), .B(\us32\/_0588_ ), .C(\us32\/_0589_ ), .D(\us32\/_0590_ ), .X(\us32\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us32/_1371_ ( .A1(\us32\/_0091_ ), .A2(\us32\/_0139_ ), .B1(\us32\/_0250_ ), .Y(\us32\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1372_ ( .A1(\us32\/_0092_ ), .A2(\us32\/_0739_ ), .B1(\us32\/_0324_ ), .B2(\us32\/_0247_ ), .Y(\us32\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1373_ ( .A1(\us32\/_0144_ ), .A2(\us32\/_0153_ ), .B1(\us32\/_0683_ ), .B2(\us32\/_0056_ ), .Y(\us32\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1374_ ( .A1(\us32\/_0091_ ), .A2(\us32\/_0499_ ), .B1(\us32\/_0330_ ), .B2(\us32\/_0056_ ), .Y(\us32\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1375_ ( .A(\us32\/_0592_ ), .B(\us32\/_0593_ ), .C(\us32\/_0594_ ), .D(\us32\/_0595_ ), .X(\us32\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1376_ ( .A(\us32\/_0499_ ), .B(\us32\/_0144_ ), .Y(\us32\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1377_ ( .A(\us32\/_0312_ ), .B(\us32\/_0598_ ), .Y(\us32\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1378_ ( .A(\us32\/_0575_ ), .B(\us32\/_0147_ ), .Y(\us32\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1379_ ( .A1(\us32\/_0293_ ), .A2(\us32\/_0137_ ), .B1(\us32\/_0093_ ), .B2(\us32\/_0739_ ), .Y(\us32\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1380_ ( .A1(\us32\/_0734_ ), .A2(\us32\/_0531_ ), .B1(\us32\/_0600_ ), .C1(\us32\/_0601_ ), .Y(\us32\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1381_ ( .A1(\us32\/_0153_ ), .A2(\us32\/_0261_ ), .B1(\us32\/_0599_ ), .C1(\us32\/_0602_ ), .Y(\us32\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1382_ ( .A(\us32\/_0591_ ), .B(\us32\/_0596_ ), .C(\us32\/_0174_ ), .D(\us32\/_0603_ ), .X(\us32\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1383_ ( .A(\us32\/_0247_ ), .B(\us32\/_0144_ ), .Y(\us32\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1384_ ( .A(\us32\/_0113_ ), .B(\us32\/_0017_ ), .Y(\us32\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1385_ ( .A(\us32\/_0381_ ), .B(\us32\/_0605_ ), .C(\us32\/_0361_ ), .D(\us32\/_0606_ ), .X(\us32\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1386_ ( .A1(\us32\/_0016_ ), .A2(\us32\/_0727_ ), .B1(\us32\/_0733_ ), .Y(\us32\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1387_ ( .A1(\us32\/_0586_ ), .A2(\us32\/_0159_ ), .B1(\us32\/_0082_ ), .B2(\us32\/_0750_ ), .Y(\us32\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1388_ ( .A1(\us32\/_0142_ ), .A2(\us32\/_0162_ ), .B1(\us32\/_0079_ ), .B2(\us32\/_0054_ ), .Y(\us32\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1389_ ( .A(\us32\/_0610_ ), .B(\us32\/_0611_ ), .C(\us32\/_0105_ ), .D(\us32\/_0106_ ), .X(\us32\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1390_ ( .A1(\us32\/_0094_ ), .A2(\us32\/_0302_ ), .B1(\us32\/_0324_ ), .B2(\us32\/_0089_ ), .Y(\us32\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1391_ ( .A(\us32\/_0607_ ), .B(\us32\/_0609_ ), .C(\us32\/_0612_ ), .D(\us32\/_0613_ ), .X(\us32\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1392_ ( .A(\us32\/_0041_ ), .B(\us32\/_0170_ ), .X(\us32\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1393_ ( .A(\us32\/_0554_ ), .B(\us32\/_0027_ ), .X(\us32\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1394_ ( .A(\us32\/_0027_ ), .B(\us32\/_0261_ ), .Y(\us32\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us32/_1395_ ( .A_N(\us32\/_0616_ ), .B(\us32\/_0617_ ), .Y(\us32\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1396_ ( .A1(\us32\/_0147_ ), .A2(\us32\/_0302_ ), .B1(\us32\/_0342_ ), .C1(\us32\/_0618_ ), .Y(\us32\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1397_ ( .A(\us32\/_0614_ ), .B(\us32\/_0272_ ), .C(\us32\/_0615_ ), .D(\us32\/_0620_ ), .X(\us32\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us32/_1398_ ( .A(\us32\/_0582_ ), .B(\us32\/_0604_ ), .C(\us32\/_0621_ ), .Y(\us32\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1399_ ( .A1(\us32\/_0280_ ), .A2(\us32\/_0134_ ), .B1(\us32\/_0089_ ), .Y(\us32\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1400_ ( .A1(\us32\/_0144_ ), .A2(\us32\/_0608_ ), .A3(\us32\/_0330_ ), .B1(\us32\/_0089_ ), .Y(\us32\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1401_ ( .A1(\us32\/_0197_ ), .A2(\us32\/_0130_ ), .A3(\us32\/_0110_ ), .B1(\us32\/_0094_ ), .Y(\us32\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1402_ ( .A(\us32\/_0432_ ), .B(\us32\/_0622_ ), .C(\us32\/_0623_ ), .D(\us32\/_0624_ ), .X(\us32\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us32/_1403_ ( .A1(\us32\/_0554_ ), .A2(\us32\/_0017_ ), .A3(\us32\/_0022_ ), .B1(\us32\/_0161_ ), .X(\us32\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us32/_1404_ ( .A_N(\us32\/_0269_ ), .B(\us32\/_0170_ ), .X(\us32\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1405_ ( .A1(\us32\/_0109_ ), .A2(\us32\/_0064_ ), .A3(\us32\/_0733_ ), .B1(\us32\/_0355_ ), .Y(\us32\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us32/_1406_ ( .A_N(\us32\/_0626_ ), .B(\us32\/_0627_ ), .C(\us32\/_0353_ ), .D(\us32\/_0628_ ), .X(\us32\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1407_ ( .A1(\us32\/_0091_ ), .A2(\us32\/_0110_ ), .A3(\us32\/_0176_ ), .B1(\us32\/_0139_ ), .Y(\us32\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1408_ ( .A1(\us32\/_0020_ ), .A2(\us32\/_0261_ ), .B1(\us32\/_0147_ ), .Y(\us32\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1409_ ( .A(\us32\/_0631_ ), .B(\us32\/_0344_ ), .C(\us32\/_0421_ ), .D(\us32\/_0632_ ), .X(\us32\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us32/_1410_ ( .A1(\us32\/_0325_ ), .A2(\us32\/_0734_ ), .B1(\us32\/_0038_ ), .C1(\us32\/_0113_ ), .X(\us32\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1411_ ( .A1(\us32\/_0134_ ), .A2(\us32\/_0114_ ), .B1(\us32\/_0221_ ), .C1(\us32\/_0634_ ), .Y(\us32\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us32/_1412_ ( .A(\us32\/_0119_ ), .B_N(\us32\/_0111_ ), .Y(\us32\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1413_ ( .A1(\us32\/_0032_ ), .A2(\us32\/_0113_ ), .B1(\us32\/_0636_ ), .C1(\us32\/_0400_ ), .Y(\us32\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1414_ ( .A1(\us32\/_0731_ ), .A2(\us32\/_0293_ ), .A3(\us32\/_0251_ ), .B1(\us32\/_0099_ ), .Y(\us32\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1415_ ( .A(\us32\/_0189_ ), .B(\us32\/_0635_ ), .C(\us32\/_0637_ ), .D(\us32\/_0638_ ), .X(\us32\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1416_ ( .A(\us32\/_0625_ ), .B(\us32\/_0630_ ), .C(\us32\/_0633_ ), .D(\us32\/_0639_ ), .X(\us32\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1417_ ( .A(\us32\/_0746_ ), .B(\us32\/_0738_ ), .X(\us32\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1418_ ( .A(\us32\/_0736_ ), .B(\us32\/_0731_ ), .X(\us32\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us32/_1419_ ( .A_N(\us32\/_0643_ ), .B(\us32\/_0577_ ), .Y(\us32\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1420_ ( .A1(\us32\/_0280_ ), .A2(\us32\/_0739_ ), .B1(\us32\/_0642_ ), .C1(\us32\/_0644_ ), .Y(\us32\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1421_ ( .A1(\us32\/_0050_ ), .A2(\us32\/_0249_ ), .B1(\us32\/_0194_ ), .C1(\us32\/_0738_ ), .Y(\us32\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1422_ ( .A(\us32\/_0646_ ), .B(\us32\/_0232_ ), .C(\us32\/_0417_ ), .D(\us32\/_0578_ ), .X(\us32\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1423_ ( .A1(\us32\/_0064_ ), .A2(\us32\/_0733_ ), .B1(\us32\/_0727_ ), .Y(\us32\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1424_ ( .A1(\us32\/_0193_ ), .A2(\us32\/_0276_ ), .B1(\us32\/_0727_ ), .Y(\us32\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1425_ ( .A(\us32\/_0645_ ), .B(\us32\/_0647_ ), .C(\us32\/_0648_ ), .D(\us32\/_0649_ ), .X(\us32\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1426_ ( .A1(\us32\/_0325_ ), .A2(\us32\/_0734_ ), .B1(\us32\/_0038_ ), .C1(\us32\/_0247_ ), .Y(\us32\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1427_ ( .A1(\us32\/_0249_ ), .A2(\us32\/_0205_ ), .B1(\us32\/_0412_ ), .C1(\us32\/_0247_ ), .Y(\us32\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1428_ ( .A(\us32\/_0652_ ), .B(\us32\/_0653_ ), .X(\us32\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1429_ ( .A1(\us32\/_0733_ ), .A2(\us32\/_0748_ ), .A3(\us32\/_0324_ ), .B1(\us32\/_0016_ ), .Y(\us32\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1430_ ( .A1(\us32\/_0640_ ), .A2(\us32\/_0193_ ), .A3(\us32\/_0091_ ), .B1(\us32\/_0016_ ), .Y(\us32\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1431_ ( .A1(\us32\/_0102_ ), .A2(\us32\/_0301_ ), .B1(\sa32\[3\] ), .C1(\us32\/_0247_ ), .Y(\us32\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1432_ ( .A(\us32\/_0654_ ), .B(\us32\/_0655_ ), .C(\us32\/_0656_ ), .D(\us32\/_0657_ ), .X(\us32\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1433_ ( .A1(\us32\/_0118_ ), .A2(\us32\/_0050_ ), .B1(\us32\/_0038_ ), .C1(\us32\/_0478_ ), .Y(\us32\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us32/_1434_ ( .A_N(\us32\/_0250_ ), .B(\us32\/_0465_ ), .C(\us32\/_0659_ ), .X(\us32\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1435_ ( .A1(\us32\/_0683_ ), .A2(\us32\/_0324_ ), .B1(\us32\/_0255_ ), .Y(\us32\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1436_ ( .A1(\us32\/_0032_ ), .A2(\us32\/_0193_ ), .A3(\us32\/_0047_ ), .B1(\us32\/_0255_ ), .Y(\us32\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1437_ ( .A1(\us32\/_0144_ ), .A2(\us32\/_0586_ ), .A3(\us32\/_0047_ ), .B1(\us32\/_0499_ ), .Y(\us32\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1438_ ( .A(\us32\/_0660_ ), .B(\us32\/_0661_ ), .C(\us32\/_0663_ ), .D(\us32\/_0664_ ), .X(\us32\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1439_ ( .A1(\us32\/_0091_ ), .A2(\us32\/_0276_ ), .B1(\us32\/_0060_ ), .Y(\us32\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1440_ ( .A1(\us32\/_0144_ ), .A2(\us32\/_0608_ ), .B1(\us32\/_0056_ ), .Y(\us32\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1441_ ( .A1(\us32\/_0412_ ), .A2(\us32\/_0038_ ), .B1(\us32\/_0102_ ), .C1(\us32\/_0060_ ), .Y(\us32\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1442_ ( .A1(\sa32\[1\] ), .A2(\us32\/_0734_ ), .B1(\us32\/_0109_ ), .C1(\us32\/_0056_ ), .Y(\us32\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1443_ ( .A(\us32\/_0666_ ), .B(\us32\/_0667_ ), .C(\us32\/_0668_ ), .D(\us32\/_0669_ ), .X(\us32\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1444_ ( .A(\us32\/_0650_ ), .B(\us32\/_0658_ ), .C(\us32\/_0665_ ), .D(\us32\/_0670_ ), .X(\us32\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us32/_1445_ ( .A(\us32\/_0641_ ), .B(\us32\/_0174_ ), .C(\us32\/_0671_ ), .Y(\us32\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us32/_1446_ ( .A(\us32\/_0049_ ), .B(\us32\/_0618_ ), .C_N(\us32\/_0052_ ), .Y(\us32\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us32/_1447_ ( .A(\us32\/_0239_ ), .Y(\us32\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1448_ ( .A(\us32\/_0705_ ), .B(\us32\/_0032_ ), .Y(\us32\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1449_ ( .A1(\us32\/_0054_ ), .A2(\us32\/_0731_ ), .B1(\us32\/_0035_ ), .B2(\us32\/_0705_ ), .Y(\us32\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1450_ ( .A1(\us32\/_0304_ ), .A2(\us32\/_0731_ ), .B1(\us32\/_0047_ ), .B2(\us32\/_0750_ ), .Y(\us32\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1451_ ( .A(\us32\/_0674_ ), .B(\us32\/_0675_ ), .C(\us32\/_0676_ ), .D(\us32\/_0677_ ), .X(\us32\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us32/_1452_ ( .A_N(\us32\/_0584_ ), .B(\us32\/_0283_ ), .X(\us32\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1453_ ( .A(\us32\/_0673_ ), .B(\us32\/_0678_ ), .C(\us32\/_0679_ ), .D(\us32\/_0508_ ), .X(\us32\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1454_ ( .A1(\us32\/_0016_ ), .A2(\us32\/_0733_ ), .B1(\us32\/_0355_ ), .B2(\us32\/_0092_ ), .Y(\us32\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1455_ ( .A(\us32\/_0681_ ), .B(\us32\/_0034_ ), .X(\us32\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us32/_1456_ ( .A1(\us32\/_0330_ ), .A2(\us32\/_0139_ ), .B1(\us32\/_0324_ ), .B2(\us32\/_0089_ ), .X(\us32\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1457_ ( .A1(\us32\/_0146_ ), .A2(\us32\/_0147_ ), .B1(\us32\/_0133_ ), .C1(\us32\/_0684_ ), .Y(\us32\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1458_ ( .A(\us32\/_0113_ ), .B(\us32\/_0251_ ), .Y(\us32\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us32/_1459_ ( .A_N(\us32\/_0463_ ), .B(\us32\/_0686_ ), .C(\us32\/_0383_ ), .D(\us32\/_0464_ ), .X(\us32\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1460_ ( .A1(\us32\/_0051_ ), .A2(\us32\/_0293_ ), .B1(\us32\/_0280_ ), .B2(\us32\/_0705_ ), .Y(\us32\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1461_ ( .A1(\us32\/_0017_ ), .A2(\us32\/_0072_ ), .B1(\us32\/_0134_ ), .B2(\us32\/_0078_ ), .Y(\us32\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1462_ ( .A(\us32\/_0687_ ), .B(\us32\/_0236_ ), .C(\us32\/_0688_ ), .D(\us32\/_0689_ ), .X(\us32\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1463_ ( .A(\us32\/_0680_ ), .B(\us32\/_0682_ ), .C(\us32\/_0685_ ), .D(\us32\/_0690_ ), .X(\us32\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us32/_1464_ ( .A1(\us32\/_0532_ ), .A2(\us32\/_0380_ ), .B1(\us32\/_0102_ ), .C1(\us32\/_0355_ ), .X(\us32\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us32/_1465_ ( .A(\us32\/_0692_ ), .B(\us32\/_0338_ ), .C(\us32\/_0644_ ), .Y(\us32\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1466_ ( .A(\us32\/_0016_ ), .B(\us32\/_0020_ ), .Y(\us32\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1467_ ( .A1(\us32\/_0032_ ), .A2(\us32\/_0137_ ), .B1(\us32\/_0279_ ), .B2(\us32\/_0094_ ), .Y(\us32\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1468_ ( .A1(\us32\/_0575_ ), .A2(\us32\/_0153_ ), .B1(\us32\/_0161_ ), .B2(\us32\/_0293_ ), .Y(\us32\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1469_ ( .A(\us32\/_0259_ ), .B(\us32\/_0695_ ), .C(\us32\/_0696_ ), .D(\us32\/_0697_ ), .X(\us32\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us32/_1470_ ( .A1(\us32\/_0255_ ), .A2(\us32\/_0640_ ), .B1(\us32\/_0016_ ), .B2(\us32\/_0193_ ), .X(\us32\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1471_ ( .A1(\us32\/_0060_ ), .A2(\us32\/_0176_ ), .B1(\us32\/_0699_ ), .C1(\us32\/_0177_ ), .Y(\us32\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1472_ ( .A1(\us32\/_0091_ ), .A2(\us32\/_0499_ ), .B1(\us32\/_0092_ ), .B2(\us32\/_0705_ ), .Y(\us32\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us32/_1473_ ( .A1(\us32\/_0705_ ), .A2(\us32\/_0683_ ), .B1(\us32\/_0093_ ), .B2(\us32\/_0114_ ), .Y(\us32\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us32/_1474_ ( .A1(\us32\/_0683_ ), .A2(\us32\/_0280_ ), .B1(\us32\/_0094_ ), .Y(\us32\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us32/_1475_ ( .A1(\us32\/_0249_ ), .A2(\us32\/_0205_ ), .B1(\us32\/_0038_ ), .C1(\us32\/_0056_ ), .Y(\us32\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1476_ ( .A(\us32\/_0701_ ), .B(\us32\/_0702_ ), .C(\us32\/_0703_ ), .D(\us32\/_0704_ ), .X(\us32\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1477_ ( .A(\us32\/_0693_ ), .B(\us32\/_0698_ ), .C(\us32\/_0700_ ), .D(\us32\/_0706_ ), .X(\us32\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us32/_1478_ ( .A1(\us32\/_0113_ ), .A2(\us32\/_0640_ ), .B1(\us32\/_0099_ ), .B2(\us32\/_0058_ ), .X(\us32\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us32/_1479_ ( .A(\us32\/_0407_ ), .B(\us32\/_0708_ ), .C(\us32\/_0529_ ), .Y(\us32\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1480_ ( .A(\us32\/_0568_ ), .B(\us32\/_0175_ ), .Y(\us32\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us32/_1481_ ( .A1(\us32\/_0247_ ), .A2(\us32\/_0114_ ), .A3(\us32\/_0051_ ), .B1(\us32\/_0130_ ), .Y(\us32\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1482_ ( .A(\us32\/_0709_ ), .B(\us32\/_0550_ ), .C(\us32\/_0710_ ), .D(\us32\/_0711_ ), .X(\us32\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us32/_1483_ ( .A1(\us32\/_0114_ ), .A2(\us32\/_0064_ ), .B1(\us32\/_0261_ ), .B2(\us32\/_0089_ ), .X(\us32\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1484_ ( .A1(\us32\/_0355_ ), .A2(\us32\/_0261_ ), .B1(\us32\/_0198_ ), .C1(\us32\/_0713_ ), .Y(\us32\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1485_ ( .A(\us32\/_0586_ ), .B(\us32\/_0478_ ), .Y(\us32\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us32/_1486_ ( .A_N(\us32\/_0541_ ), .B(\us32\/_0267_ ), .C(\us32\/_0715_ ), .D(\us32\/_0320_ ), .X(\us32\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1487_ ( .A(\us32\/_0586_ ), .B(\us32\/_0070_ ), .Y(\us32\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us32/_1488_ ( .A_N(\us32\/_0211_ ), .B(\us32\/_0155_ ), .C(\us32\/_0202_ ), .D(\us32\/_0718_ ), .X(\us32\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us32/_1489_ ( .A(\us32\/_0150_ ), .B(\us32\/_0205_ ), .C(\us32\/_0380_ ), .Y(\us32\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us32/_1490_ ( .A(\us32\/_0411_ ), .B(\us32\/_0720_ ), .X(\us32\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us32/_1491_ ( .A1(\us32\/_0017_ ), .A2(\us32\/_0022_ ), .B1(\us32\/_0078_ ), .X(\us32\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us32/_1492_ ( .A1(\us32\/_0134_ ), .A2(\us32\/_0738_ ), .B1(\us32\/_0101_ ), .C1(\us32\/_0722_ ), .Y(\us32\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1493_ ( .A(\us32\/_0717_ ), .B(\us32\/_0719_ ), .C(\us32\/_0721_ ), .D(\us32\/_0723_ ), .X(\us32\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us32/_1494_ ( .A(\us32\/_0739_ ), .B(\us32\/_0193_ ), .Y(\us32\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1495_ ( .A(\us32\/_0344_ ), .B(\us32\/_0184_ ), .C(\us32\/_0449_ ), .D(\us32\/_0725_ ), .X(\us32\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us32/_1496_ ( .A(\us32\/_0712_ ), .B(\us32\/_0714_ ), .C(\us32\/_0724_ ), .D(\us32\/_0726_ ), .X(\us32\/_0728_ ) );
sky130_fd_sc_hd__nand3_1 \us32/_1497_ ( .A(\us32\/_0691_ ), .B(\us32\/_0707_ ), .C(\us32\/_0728_ ), .Y(\us32\/_0015_ ) );
sky130_fd_sc_hd__nor2b_1 \us33/_0753_ ( .A(\sa33\[2\] ), .B_N(\sa33\[3\] ), .Y(\us33\/_0096_ ) );
sky130_fd_sc_hd__and2_1 \us33/_0755_ ( .A(\sa33\[1\] ), .B(\sa33\[0\] ), .X(\us33\/_0118_ ) );
sky130_fd_sc_hd__and2_1 \us33/_0756_ ( .A(\us33\/_0096_ ), .B(\us33\/_0118_ ), .X(\us33\/_0129_ ) );
sky130_fd_sc_hd__and2_1 \us33/_0757_ ( .A(\sa33\[7\] ), .B(\sa33\[6\] ), .X(\us33\/_0140_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_0758_ ( .A(\sa33\[4\] ), .B(\sa33\[5\] ), .Y(\us33\/_0151_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0759_ ( .A(\us33\/_0140_ ), .B(\us33\/_0151_ ), .X(\us33\/_0162_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0761_ ( .A(\us33\/_0129_ ), .B(\us33\/_0162_ ), .X(\us33\/_0183_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0762_ ( .A(\us33\/_0096_ ), .X(\us33\/_0194_ ) );
sky130_fd_sc_hd__nor2b_1 \us33/_0763_ ( .A(\sa33\[1\] ), .B_N(\sa33\[0\] ), .Y(\us33\/_0205_ ) );
sky130_fd_sc_hd__and3_1 \us33/_0765_ ( .A(\us33\/_0162_ ), .B(\us33\/_0194_ ), .C(\us33\/_0205_ ), .X(\us33\/_0227_ ) );
sky130_fd_sc_hd__lpflow_inputiso1p_1 \us33/_0766_ ( .A(\us33\/_0183_ ), .SLEEP(\us33\/_0227_ ), .X(\us33\/_0238_ ) );
sky130_fd_sc_hd__nor2b_1 \us33/_0767_ ( .A(\sa33\[0\] ), .B_N(\sa33\[1\] ), .Y(\us33\/_0249_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_0768_ ( .A(\sa33\[2\] ), .B(\sa33\[3\] ), .Y(\us33\/_0260_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0769_ ( .A(\us33\/_0249_ ), .B(\us33\/_0260_ ), .X(\us33\/_0271_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0771_ ( .A(\us33\/_0271_ ), .X(\us33\/_0293_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0772_ ( .A(\us33\/_0162_ ), .X(\us33\/_0304_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_0773_ ( .A(\us33\/_0293_ ), .B(\us33\/_0304_ ), .Y(\us33\/_0314_ ) );
sky130_fd_sc_hd__inv_2 \us33/_0774_ ( .A(\sa33\[1\] ), .Y(\us33\/_0325_ ) );
sky130_fd_sc_hd__inv_2 \us33/_0776_ ( .A(\sa33\[0\] ), .Y(\us33\/_0347_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0777_ ( .A(\sa33\[2\] ), .B(\sa33\[3\] ), .X(\us33\/_0358_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0779_ ( .A(\us33\/_0358_ ), .X(\us33\/_0380_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_0780_ ( .A1(\us33\/_0325_ ), .A2(\us33\/_0347_ ), .B1(\us33\/_0380_ ), .C1(\us33\/_0304_ ), .Y(\us33\/_0391_ ) );
sky130_fd_sc_hd__and3b_1 \us33/_0781_ ( .A_N(\us33\/_0238_ ), .B(\us33\/_0314_ ), .C(\us33\/_0391_ ), .X(\us33\/_0401_ ) );
sky130_fd_sc_hd__nor2b_1 \us33/_0782_ ( .A(\sa33\[3\] ), .B_N(\sa33\[2\] ), .Y(\us33\/_0412_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0784_ ( .A(\us33\/_0412_ ), .B(\us33\/_0205_ ), .X(\us33\/_0434_ ) );
sky130_fd_sc_hd__nor2b_1 \us33/_0787_ ( .A(\sa33\[5\] ), .B_N(\sa33\[4\] ), .Y(\us33\/_0467_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0788_ ( .A(\us33\/_0467_ ), .B(\us33\/_0140_ ), .X(\us33\/_0478_ ) );
sky130_fd_sc_hd__buf_2 \us33/_0790_ ( .A(\us33\/_0478_ ), .X(\us33\/_0499_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_0791_ ( .A(\us33\/_0134_ ), .B(\us33\/_0499_ ), .Y(\us33\/_0510_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_0792_ ( .A(\us33\/_0478_ ), .B(\us33\/_0271_ ), .Y(\us33\/_0521_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0793_ ( .A(\us33\/_0194_ ), .X(\us33\/_0532_ ) );
sky130_fd_sc_hd__and2_1 \us33/_0795_ ( .A(\us33\/_0249_ ), .B(\us33\/_0358_ ), .X(\us33\/_0554_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0797_ ( .A(\us33\/_0554_ ), .X(\us33\/_0575_ ) );
sky130_fd_sc_hd__and2_1 \us33/_0798_ ( .A(\us33\/_0205_ ), .B(\us33\/_0358_ ), .X(\us33\/_0586_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0800_ ( .A(\us33\/_0586_ ), .X(\us33\/_0608_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_0801_ ( .A1(\us33\/_0532_ ), .A2(\us33\/_0575_ ), .A3(\us33\/_0608_ ), .B1(\us33\/_0499_ ), .Y(\us33\/_0619_ ) );
sky130_fd_sc_hd__and4_1 \us33/_0802_ ( .A(\us33\/_0401_ ), .B(\us33\/_0510_ ), .C(\us33\/_0521_ ), .D(\us33\/_0619_ ), .X(\us33\/_0629_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0803_ ( .A(\us33\/_0358_ ), .B(\sa33\[1\] ), .X(\us33\/_0640_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0805_ ( .A(\us33\/_0205_ ), .B(\us33\/_0260_ ), .X(\us33\/_0662_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0807_ ( .A(\us33\/_0662_ ), .X(\us33\/_0683_ ) );
sky130_fd_sc_hd__nor2b_1 \us33/_0808_ ( .A(\sa33\[6\] ), .B_N(\sa33\[7\] ), .Y(\us33\/_0694_ ) );
sky130_fd_sc_hd__and2_1 \us33/_0809_ ( .A(\us33\/_0467_ ), .B(\us33\/_0694_ ), .X(\us33\/_0705_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0811_ ( .A(\us33\/_0705_ ), .X(\us33\/_0727_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_0812_ ( .A1(\us33\/_0640_ ), .A2(\us33\/_0293_ ), .A3(\us33\/_0683_ ), .B1(\us33\/_0727_ ), .Y(\us33\/_0729_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_0813_ ( .A(\sa33\[1\] ), .B(\sa33\[0\] ), .Y(\us33\/_0730_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0814_ ( .A(\us33\/_0730_ ), .B(\us33\/_0260_ ), .X(\us33\/_0731_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0816_ ( .A(\us33\/_0731_ ), .X(\us33\/_0733_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0817_ ( .A(\sa33\[0\] ), .X(\us33\/_0734_ ) );
sky130_fd_sc_hd__o21a_1 \us33/_0818_ ( .A1(\us33\/_0325_ ), .A2(\us33\/_0734_ ), .B1(\us33\/_0412_ ), .X(\us33\/_0735_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0819_ ( .A(\us33\/_0694_ ), .B(\us33\/_0151_ ), .X(\us33\/_0736_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0821_ ( .A(\us33\/_0736_ ), .X(\us33\/_0738_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0822_ ( .A(\us33\/_0738_ ), .X(\us33\/_0739_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_0823_ ( .A1(\us33\/_0733_ ), .A2(\us33\/_0735_ ), .A3(\us33\/_0293_ ), .B1(\us33\/_0739_ ), .Y(\us33\/_0740_ ) );
sky130_fd_sc_hd__nor2b_1 \us33/_0824_ ( .A(\us33\/_0730_ ), .B_N(\us33\/_0358_ ), .Y(\us33\/_0741_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_0825_ ( .A(\us33\/_0741_ ), .B(\us33\/_0739_ ), .Y(\us33\/_0742_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_0827_ ( .A1(\us33\/_0118_ ), .A2(\us33\/_0205_ ), .B1(\us33\/_0532_ ), .C1(\us33\/_0739_ ), .Y(\us33\/_0744_ ) );
sky130_fd_sc_hd__and4_1 \us33/_0828_ ( .A(\us33\/_0729_ ), .B(\us33\/_0740_ ), .C(\us33\/_0742_ ), .D(\us33\/_0744_ ), .X(\us33\/_0745_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0829_ ( .A(\us33\/_0412_ ), .B(\us33\/_0730_ ), .X(\us33\/_0746_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0831_ ( .A(\us33\/_0746_ ), .X(\us33\/_0748_ ) );
sky130_fd_sc_hd__nor2b_1 \us33/_0832_ ( .A(\sa33\[4\] ), .B_N(\sa33\[5\] ), .Y(\us33\/_0749_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0833_ ( .A(\us33\/_0749_ ), .B(\us33\/_0694_ ), .X(\us33\/_0750_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0835_ ( .A(\us33\/_0750_ ), .X(\us33\/_0752_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0836_ ( .A(\us33\/_0752_ ), .X(\us33\/_0016_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0837_ ( .A(\us33\/_0118_ ), .B(\us33\/_0358_ ), .X(\us33\/_0017_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0839_ ( .A(\us33\/_0752_ ), .B(\us33\/_0017_ ), .X(\us33\/_0019_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0840_ ( .A(\us33\/_0358_ ), .B(\us33\/_0325_ ), .X(\us33\/_0020_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0842_ ( .A(\us33\/_0096_ ), .B(\us33\/_0205_ ), .X(\us33\/_0022_ ) );
sky130_fd_sc_hd__o21a_1 \us33/_0844_ ( .A1(\us33\/_0020_ ), .A2(\us33\/_0022_ ), .B1(\us33\/_0752_ ), .X(\us33\/_0024_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_0845_ ( .A1(\us33\/_0748_ ), .A2(\us33\/_0016_ ), .B1(\us33\/_0019_ ), .C1(\us33\/_0024_ ), .Y(\us33\/_0025_ ) );
sky130_fd_sc_hd__and2_1 \us33/_0846_ ( .A(\sa33\[4\] ), .B(\sa33\[5\] ), .X(\us33\/_0026_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0847_ ( .A(\us33\/_0694_ ), .B(\us33\/_0026_ ), .X(\us33\/_0027_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0850_ ( .A(\us33\/_0358_ ), .B(\us33\/_0730_ ), .X(\us33\/_0030_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0852_ ( .A(\us33\/_0030_ ), .X(\us33\/_0032_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_0853_ ( .A(\us33\/_0247_ ), .B(\us33\/_0032_ ), .Y(\us33\/_0033_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_0854_ ( .A(\us33\/_0247_ ), .B(\us33\/_0735_ ), .Y(\us33\/_0034_ ) );
sky130_fd_sc_hd__and2_1 \us33/_0855_ ( .A(\us33\/_0118_ ), .B(\us33\/_0260_ ), .X(\us33\/_0035_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0857_ ( .A(\us33\/_0027_ ), .B(\us33\/_0035_ ), .X(\us33\/_0037_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0858_ ( .A(\us33\/_0260_ ), .X(\us33\/_0038_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_0859_ ( .A(\us33\/_0038_ ), .B(\us33\/_0347_ ), .Y(\us33\/_0039_ ) );
sky130_fd_sc_hd__and2b_1 \us33/_0860_ ( .A_N(\us33\/_0039_ ), .B(\us33\/_0027_ ), .X(\us33\/_0040_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_0861_ ( .A(\us33\/_0037_ ), .B(\us33\/_0040_ ), .Y(\us33\/_0041_ ) );
sky130_fd_sc_hd__and4_1 \us33/_0862_ ( .A(\us33\/_0025_ ), .B(\us33\/_0033_ ), .C(\us33\/_0034_ ), .D(\us33\/_0041_ ), .X(\us33\/_0042_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0863_ ( .A(\us33\/_0749_ ), .B(\us33\/_0140_ ), .X(\us33\/_0043_ ) );
sky130_fd_sc_hd__and3_1 \us33/_0865_ ( .A(\sa33\[0\] ), .B(\sa33\[2\] ), .C(\sa33\[3\] ), .X(\us33\/_0045_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0866_ ( .A(\us33\/_0043_ ), .B(\us33\/_0045_ ), .X(\us33\/_0046_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0867_ ( .A(\us33\/_0096_ ), .B(\us33\/_0249_ ), .X(\us33\/_0047_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0869_ ( .A(\us33\/_0047_ ), .B(\us33\/_0043_ ), .X(\us33\/_0049_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0870_ ( .A(\us33\/_0730_ ), .X(\us33\/_0050_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0871_ ( .A(\us33\/_0043_ ), .X(\us33\/_0051_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_0872_ ( .A1(\us33\/_0118_ ), .A2(\us33\/_0050_ ), .B1(\us33\/_0194_ ), .C1(\us33\/_0051_ ), .Y(\us33\/_0052_ ) );
sky130_fd_sc_hd__nor3b_1 \us33/_0873_ ( .A(\us33\/_0046_ ), .B(\us33\/_0049_ ), .C_N(\us33\/_0052_ ), .Y(\us33\/_0053_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0874_ ( .A(\us33\/_0026_ ), .B(\us33\/_0140_ ), .X(\us33\/_0054_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_0877_ ( .A1(\us33\/_0532_ ), .A2(\us33\/_0575_ ), .B1(\us33\/_0292_ ), .Y(\us33\/_0057_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0878_ ( .A(\us33\/_0412_ ), .B(\us33\/_0325_ ), .X(\us33\/_0058_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0880_ ( .A(\us33\/_0051_ ), .X(\us33\/_0060_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_0881_ ( .A1(\us33\/_0731_ ), .A2(\us33\/_0035_ ), .A3(\us33\/_0058_ ), .B1(\us33\/_0060_ ), .Y(\us33\/_0061_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0882_ ( .A(\us33\/_0260_ ), .B(\sa33\[1\] ), .X(\us33\/_0062_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0884_ ( .A(\us33\/_0062_ ), .X(\us33\/_0064_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_0885_ ( .A1(\us33\/_0064_ ), .A2(\us33\/_0748_ ), .A3(\us33\/_0683_ ), .B1(\us33\/_0292_ ), .Y(\us33\/_0065_ ) );
sky130_fd_sc_hd__and4_1 \us33/_0886_ ( .A(\us33\/_0053_ ), .B(\us33\/_0057_ ), .C(\us33\/_0061_ ), .D(\us33\/_0065_ ), .X(\us33\/_0066_ ) );
sky130_fd_sc_hd__and4_1 \us33/_0887_ ( .A(\us33\/_0629_ ), .B(\us33\/_0745_ ), .C(\us33\/_0042_ ), .D(\us33\/_0066_ ), .X(\us33\/_0067_ ) );
sky130_fd_sc_hd__nor2b_1 \us33/_0889_ ( .A(\sa33\[7\] ), .B_N(\sa33\[6\] ), .Y(\us33\/_0069_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0890_ ( .A(\us33\/_0069_ ), .B(\us33\/_0151_ ), .X(\us33\/_0070_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0892_ ( .A(\us33\/_0070_ ), .X(\us33\/_0072_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_0893_ ( .A1(\us33\/_0129_ ), .A2(\us33\/_0586_ ), .B1(\us33\/_0072_ ), .Y(\us33\/_0073_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_0894_ ( .A1(\us33\/_0380_ ), .A2(\us33\/_0347_ ), .B1(\us33\/_0194_ ), .B2(\us33\/_0205_ ), .Y(\us33\/_0074_ ) );
sky130_fd_sc_hd__nor2b_1 \us33/_0895_ ( .A(\us33\/_0074_ ), .B_N(\us33\/_0070_ ), .Y(\us33\/_0075_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us33/_0896_ ( .A(\us33\/_0073_ ), .SLEEP(\us33\/_0075_ ), .X(\us33\/_0076_ ) );
sky130_fd_sc_hd__and2_1 \us33/_0897_ ( .A(\us33\/_0467_ ), .B(\us33\/_0069_ ), .X(\us33\/_0077_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0898_ ( .A(\us33\/_0077_ ), .X(\us33\/_0078_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0899_ ( .A(\us33\/_0412_ ), .B(\us33\/_0118_ ), .X(\us33\/_0079_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0901_ ( .A(\us33\/_0078_ ), .B(\us33\/_0079_ ), .X(\us33\/_0081_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0902_ ( .A(\us33\/_0412_ ), .B(\us33\/_0249_ ), .X(\us33\/_0082_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0905_ ( .A(\us33\/_0280_ ), .B(\us33\/_0078_ ), .X(\us33\/_0085_ ) );
sky130_fd_sc_hd__o21ai_1 \us33/_0906_ ( .A1(\sa33\[0\] ), .A2(\us33\/_0325_ ), .B1(\us33\/_0260_ ), .Y(\us33\/_0086_ ) );
sky130_fd_sc_hd__and2b_1 \us33/_0907_ ( .A_N(\us33\/_0086_ ), .B(\us33\/_0078_ ), .X(\us33\/_0087_ ) );
sky130_fd_sc_hd__nor3_1 \us33/_0908_ ( .A(\us33\/_0081_ ), .B(\us33\/_0085_ ), .C(\us33\/_0087_ ), .Y(\us33\/_0088_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0909_ ( .A(\us33\/_0072_ ), .X(\us33\/_0089_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_0910_ ( .A1(\us33\/_0733_ ), .A2(\us33\/_0748_ ), .A3(\us33\/_0683_ ), .B1(\us33\/_0089_ ), .Y(\us33\/_0090_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0911_ ( .A(\us33\/_0129_ ), .X(\us33\/_0091_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0912_ ( .A(\us33\/_0017_ ), .X(\us33\/_0092_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0913_ ( .A(\us33\/_0022_ ), .X(\us33\/_0093_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0914_ ( .A(\us33\/_0078_ ), .X(\us33\/_0094_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_0915_ ( .A1(\us33\/_0091_ ), .A2(\us33\/_0092_ ), .A3(\us33\/_0093_ ), .B1(\us33\/_0094_ ), .Y(\us33\/_0095_ ) );
sky130_fd_sc_hd__and4_1 \us33/_0916_ ( .A(\us33\/_0076_ ), .B(\us33\/_0088_ ), .C(\us33\/_0090_ ), .D(\us33\/_0095_ ), .X(\us33\/_0097_ ) );
sky130_fd_sc_hd__and2_1 \us33/_0917_ ( .A(\us33\/_0069_ ), .B(\us33\/_0026_ ), .X(\us33\/_0098_ ) );
sky130_fd_sc_hd__buf_2 \us33/_0918_ ( .A(\us33\/_0098_ ), .X(\us33\/_0099_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0919_ ( .A(\us33\/_0434_ ), .B(\us33\/_0099_ ), .X(\us33\/_0100_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0920_ ( .A(\us33\/_0079_ ), .B(\us33\/_0098_ ), .X(\us33\/_0101_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0921_ ( .A(\us33\/_0325_ ), .X(\us33\/_0102_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_0922_ ( .A1(\us33\/_0102_ ), .A2(\us33\/_0734_ ), .B1(\us33\/_0038_ ), .C1(\us33\/_0099_ ), .Y(\us33\/_0103_ ) );
sky130_fd_sc_hd__nor3b_1 \us33/_0923_ ( .A(\us33\/_0100_ ), .B(\us33\/_0101_ ), .C_N(\us33\/_0103_ ), .Y(\us33\/_0104_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_0924_ ( .A1(\us33\/_0554_ ), .A2(\us33\/_0586_ ), .B1(\us33\/_0099_ ), .Y(\us33\/_0105_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_0925_ ( .A(\us33\/_0129_ ), .B(\us33\/_0099_ ), .Y(\us33\/_0106_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0926_ ( .A(\us33\/_0105_ ), .B(\us33\/_0106_ ), .X(\us33\/_0108_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0927_ ( .A(\us33\/_0412_ ), .X(\us33\/_0109_ ) );
sky130_fd_sc_hd__and2_1 \us33/_0928_ ( .A(\us33\/_0260_ ), .B(\sa33\[0\] ), .X(\us33\/_0110_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0929_ ( .A(\us33\/_0069_ ), .B(\us33\/_0749_ ), .X(\us33\/_0111_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0931_ ( .A(\us33\/_0111_ ), .X(\us33\/_0113_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0932_ ( .A(\us33\/_0113_ ), .X(\us33\/_0114_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_0933_ ( .A1(\us33\/_0109_ ), .A2(\us33\/_0110_ ), .B1(\us33\/_0114_ ), .Y(\us33\/_0115_ ) );
sky130_fd_sc_hd__inv_1 \us33/_0934_ ( .A(\us33\/_0022_ ), .Y(\us33\/_0116_ ) );
sky130_fd_sc_hd__inv_1 \us33/_0935_ ( .A(\us33\/_0554_ ), .Y(\us33\/_0117_ ) );
sky130_fd_sc_hd__o21ai_1 \us33/_0936_ ( .A1(\us33\/_0050_ ), .A2(\us33\/_0118_ ), .B1(\us33\/_0194_ ), .Y(\us33\/_0119_ ) );
sky130_fd_sc_hd__inv_1 \us33/_0937_ ( .A(\us33\/_0113_ ), .Y(\us33\/_0120_ ) );
sky130_fd_sc_hd__a31o_1 \us33/_0938_ ( .A1(\us33\/_0116_ ), .A2(\us33\/_0117_ ), .A3(\us33\/_0119_ ), .B1(\us33\/_0120_ ), .X(\us33\/_0121_ ) );
sky130_fd_sc_hd__and4_1 \us33/_0939_ ( .A(\us33\/_0104_ ), .B(\us33\/_0108_ ), .C(\us33\/_0115_ ), .D(\us33\/_0121_ ), .X(\us33\/_0122_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_0940_ ( .A(\sa33\[7\] ), .B(\sa33\[6\] ), .Y(\us33\/_0123_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0941_ ( .A(\us33\/_0749_ ), .B(\us33\/_0123_ ), .X(\us33\/_0124_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0943_ ( .A(\us33\/_0082_ ), .B(\us33\/_0124_ ), .X(\us33\/_0126_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_0944_ ( .A(\us33\/_0271_ ), .B(\us33\/_0124_ ), .Y(\us33\/_0127_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0945_ ( .A(\us33\/_0124_ ), .X(\us33\/_0128_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0946_ ( .A(\us33\/_0260_ ), .B(\us33\/_0325_ ), .X(\us33\/_0130_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_0948_ ( .A(\us33\/_0128_ ), .B(\us33\/_0130_ ), .Y(\us33\/_0132_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_0949_ ( .A(\us33\/_0127_ ), .B(\us33\/_0132_ ), .Y(\us33\/_0133_ ) );
sky130_fd_sc_hd__buf_2 \us33/_0950_ ( .A(\us33\/_0434_ ), .X(\us33\/_0134_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_0951_ ( .A(\us33\/_0134_ ), .B(\us33\/_0128_ ), .Y(\us33\/_0135_ ) );
sky130_fd_sc_hd__nor3b_1 \us33/_0952_ ( .A(\us33\/_0126_ ), .B(\us33\/_0133_ ), .C_N(\us33\/_0135_ ), .Y(\us33\/_0136_ ) );
sky130_fd_sc_hd__and2_1 \us33/_0953_ ( .A(\us33\/_0026_ ), .B(\us33\/_0123_ ), .X(\us33\/_0137_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0955_ ( .A(\us33\/_0137_ ), .X(\us33\/_0139_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_0956_ ( .A1(\us33\/_0110_ ), .A2(\us33\/_0293_ ), .A3(\us33\/_0280_ ), .B1(\us33\/_0139_ ), .Y(\us33\/_0141_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0957_ ( .A(\us33\/_0096_ ), .B(\us33\/_0730_ ), .X(\us33\/_0142_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0959_ ( .A(\us33\/_0142_ ), .X(\us33\/_0144_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_0960_ ( .A1(\us33\/_0020_ ), .A2(\us33\/_0144_ ), .A3(\us33\/_0017_ ), .B1(\us33\/_0139_ ), .Y(\us33\/_0145_ ) );
sky130_fd_sc_hd__nor3b_1 \us33/_0961_ ( .A(\sa33\[2\] ), .B(\us33\/_0050_ ), .C_N(\sa33\[3\] ), .Y(\us33\/_0146_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0962_ ( .A(\us33\/_0128_ ), .X(\us33\/_0147_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_0963_ ( .A1(\us33\/_0146_ ), .A2(\us33\/_0032_ ), .A3(\us33\/_0640_ ), .B1(\us33\/_0147_ ), .Y(\us33\/_0148_ ) );
sky130_fd_sc_hd__and4_1 \us33/_0964_ ( .A(\us33\/_0136_ ), .B(\us33\/_0141_ ), .C(\us33\/_0145_ ), .D(\us33\/_0148_ ), .X(\us33\/_0149_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0965_ ( .A(\us33\/_0123_ ), .B(\us33\/_0151_ ), .X(\us33\/_0150_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0967_ ( .A(\us33\/_0150_ ), .X(\us33\/_0153_ ) );
sky130_fd_sc_hd__and2_1 \us33/_0968_ ( .A(\us33\/_0150_ ), .B(\us33\/_0062_ ), .X(\us33\/_0154_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_0969_ ( .A(\us33\/_0079_ ), .B(\us33\/_0150_ ), .Y(\us33\/_0155_ ) );
sky130_fd_sc_hd__nand3_1 \us33/_0970_ ( .A(\us33\/_0150_ ), .B(\us33\/_0412_ ), .C(\us33\/_0249_ ), .Y(\us33\/_0156_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_0971_ ( .A(\us33\/_0155_ ), .B(\us33\/_0156_ ), .Y(\us33\/_0157_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_0972_ ( .A1(\us33\/_0153_ ), .A2(\us33\/_0134_ ), .B1(\us33\/_0154_ ), .C1(\us33\/_0157_ ), .Y(\us33\/_0158_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0973_ ( .A(\us33\/_0467_ ), .B(\us33\/_0123_ ), .X(\us33\/_0159_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_0975_ ( .A(\us33\/_0159_ ), .X(\us33\/_0161_ ) );
sky130_fd_sc_hd__and2b_1 \us33/_0976_ ( .A_N(\us33\/_0119_ ), .B(\us33\/_0161_ ), .X(\us33\/_0163_ ) );
sky130_fd_sc_hd__inv_1 \us33/_0977_ ( .A(\us33\/_0163_ ), .Y(\us33\/_0164_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_0978_ ( .A1(\us33\/_0146_ ), .A2(\us33\/_0575_ ), .A3(\us33\/_0608_ ), .B1(\us33\/_0153_ ), .Y(\us33\/_0165_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_0979_ ( .A1(\us33\/_0062_ ), .A2(\us33\/_0280_ ), .A3(\us33\/_0134_ ), .B1(\us33\/_0161_ ), .Y(\us33\/_0166_ ) );
sky130_fd_sc_hd__and4_1 \us33/_0980_ ( .A(\us33\/_0158_ ), .B(\us33\/_0164_ ), .C(\us33\/_0165_ ), .D(\us33\/_0166_ ), .X(\us33\/_0167_ ) );
sky130_fd_sc_hd__and4_1 \us33/_0981_ ( .A(\us33\/_0097_ ), .B(\us33\/_0122_ ), .C(\us33\/_0149_ ), .D(\us33\/_0167_ ), .X(\us33\/_0168_ ) );
sky130_fd_sc_hd__and2_1 \us33/_0982_ ( .A(\us33\/_0662_ ), .B(\us33\/_0150_ ), .X(\us33\/_0169_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_0983_ ( .A(\us33\/_0154_ ), .B(\us33\/_0169_ ), .Y(\us33\/_0170_ ) );
sky130_fd_sc_hd__and3_1 \us33/_0984_ ( .A(\us33\/_0123_ ), .B(\us33\/_0151_ ), .C(\us33\/_0038_ ), .X(\us33\/_0171_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0985_ ( .A(\us33\/_0170_ ), .B(\us33\/_0171_ ), .X(\us33\/_0172_ ) );
sky130_fd_sc_hd__inv_1 \us33/_0986_ ( .A(\us33\/_0172_ ), .Y(\us33\/_0174_ ) );
sky130_fd_sc_hd__nand3_1 \us33/_0987_ ( .A(\us33\/_0067_ ), .B(\us33\/_0168_ ), .C(\us33\/_0174_ ), .Y(\us33\/_0008_ ) );
sky130_fd_sc_hd__xnor2_1 \us33/_0988_ ( .A(\sa33\[1\] ), .B(\sa33\[0\] ), .Y(\us33\/_0175_ ) );
sky130_fd_sc_hd__and2_1 \us33/_0989_ ( .A(\us33\/_0175_ ), .B(\us33\/_0358_ ), .X(\us33\/_0176_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0990_ ( .A(\us33\/_0176_ ), .B(\us33\/_0478_ ), .X(\us33\/_0177_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_0991_ ( .A(\us33\/_0280_ ), .B(\us33\/_0113_ ), .Y(\us33\/_0178_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0992_ ( .A(\us33\/_0111_ ), .B(\us33\/_0062_ ), .X(\us33\/_0179_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0993_ ( .A(\us33\/_0111_ ), .B(\us33\/_0662_ ), .X(\us33\/_0180_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_0994_ ( .A(\us33\/_0179_ ), .B(\us33\/_0180_ ), .Y(\us33\/_0181_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0995_ ( .A(\us33\/_0054_ ), .B(\us33\/_0058_ ), .X(\us33\/_0182_ ) );
sky130_fd_sc_hd__inv_1 \us33/_0996_ ( .A(\us33\/_0182_ ), .Y(\us33\/_0184_ ) );
sky130_fd_sc_hd__and4b_1 \us33/_0997_ ( .A_N(\us33\/_0177_ ), .B(\us33\/_0178_ ), .C(\us33\/_0181_ ), .D(\us33\/_0184_ ), .X(\us33\/_0185_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0998_ ( .A(\us33\/_0098_ ), .B(\us33\/_0741_ ), .X(\us33\/_0186_ ) );
sky130_fd_sc_hd__and2_0 \us33/_0999_ ( .A(\us33\/_0047_ ), .B(\us33\/_0098_ ), .X(\us33\/_0187_ ) );
sky130_fd_sc_hd__or2_0 \us33/_1000_ ( .A(\us33\/_0186_ ), .B(\us33\/_0187_ ), .X(\us33\/_0188_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1001_ ( .A(\us33\/_0188_ ), .Y(\us33\/_0189_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1002_ ( .A(\us33\/_0738_ ), .B(\us33\/_0735_ ), .X(\us33\/_0190_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1003_ ( .A(\us33\/_0271_ ), .B(\us33\/_0736_ ), .X(\us33\/_0191_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_1004_ ( .A(\us33\/_0190_ ), .B(\us33\/_0191_ ), .Y(\us33\/_0192_ ) );
sky130_fd_sc_hd__and2_1 \us33/_1005_ ( .A(\us33\/_0096_ ), .B(\us33\/_0325_ ), .X(\us33\/_0193_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1006_ ( .A1(\us33\/_0193_ ), .A2(\us33\/_0176_ ), .B1(\us33\/_0043_ ), .Y(\us33\/_0195_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1007_ ( .A(\us33\/_0185_ ), .B(\us33\/_0189_ ), .C(\us33\/_0192_ ), .D(\us33\/_0195_ ), .X(\us33\/_0196_ ) );
sky130_fd_sc_hd__and3b_1 \us33/_1008_ ( .A_N(\sa33\[3\] ), .B(\us33\/_0734_ ), .C(\sa33\[2\] ), .X(\us33\/_0197_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1009_ ( .A(\us33\/_0137_ ), .B(\us33\/_0197_ ), .X(\us33\/_0198_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_1010_ ( .A(\us33\/_0198_ ), .B(\us33\/_0040_ ), .Y(\us33\/_0199_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1011_ ( .A(\us33\/_0293_ ), .B(\us33\/_0137_ ), .X(\us33\/_0200_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1012_ ( .A(\us33\/_0200_ ), .Y(\us33\/_0201_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1013_ ( .A(\us33\/_0137_ ), .B(\us33\/_0110_ ), .Y(\us33\/_0202_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1014_ ( .A(\us33\/_0139_ ), .B(\us33\/_0020_ ), .Y(\us33\/_0203_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1015_ ( .A(\us33\/_0199_ ), .B(\us33\/_0201_ ), .C(\us33\/_0202_ ), .D(\us33\/_0203_ ), .X(\us33\/_0204_ ) );
sky130_fd_sc_hd__o211a_1 \us33/_1016_ ( .A1(\us33\/_0532_ ), .A2(\us33\/_0109_ ), .B1(\us33\/_0102_ ), .C1(\us33\/_0727_ ), .X(\us33\/_0206_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1017_ ( .A(\us33\/_0022_ ), .B(\us33\/_0078_ ), .Y(\us33\/_0207_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1018_ ( .A(\us33\/_0078_ ), .B(\us33\/_0142_ ), .Y(\us33\/_0208_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1019_ ( .A(\us33\/_0207_ ), .B(\us33\/_0208_ ), .Y(\us33\/_0209_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1020_ ( .A1(\us33\/_0094_ ), .A2(\us33\/_0176_ ), .B1(\us33\/_0206_ ), .C1(\us33\/_0209_ ), .Y(\us33\/_0210_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1021_ ( .A(\us33\/_0662_ ), .B(\us33\/_0070_ ), .X(\us33\/_0211_ ) );
sky130_fd_sc_hd__nand3_1 \us33/_1022_ ( .A(\us33\/_0731_ ), .B(\us33\/_0123_ ), .C(\us33\/_0749_ ), .Y(\us33\/_0212_ ) );
sky130_fd_sc_hd__nand3_1 \us33/_1023_ ( .A(\us33\/_0731_ ), .B(\us33\/_0467_ ), .C(\us33\/_0069_ ), .Y(\us33\/_0213_ ) );
sky130_fd_sc_hd__and4b_1 \us33/_1024_ ( .A_N(\us33\/_0211_ ), .B(\us33\/_0127_ ), .C(\us33\/_0212_ ), .D(\us33\/_0213_ ), .X(\us33\/_0214_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1025_ ( .A(\us33\/_0137_ ), .Y(\us33\/_0215_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1026_ ( .A(\us33\/_0128_ ), .B(\us33\/_0035_ ), .Y(\us33\/_0217_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1028_ ( .A1(\us33\/_0159_ ), .A2(\us33\/_0746_ ), .B1(\us33\/_0434_ ), .B2(\us33\/_0499_ ), .Y(\us33\/_0219_ ) );
sky130_fd_sc_hd__o211a_1 \us33/_1029_ ( .A1(\us33\/_0116_ ), .A2(\us33\/_0215_ ), .B1(\us33\/_0217_ ), .C1(\us33\/_0219_ ), .X(\us33\/_0220_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1030_ ( .A(\us33\/_0113_ ), .B(\us33\/_0746_ ), .X(\us33\/_0221_ ) );
sky130_fd_sc_hd__a22o_1 \us33/_1031_ ( .A1(\us33\/_0098_ ), .A2(\us33\/_0746_ ), .B1(\us33\/_0434_ ), .B2(\us33\/_0750_ ), .X(\us33\/_0222_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1032_ ( .A1(\us33\/_0047_ ), .A2(\us33\/_0113_ ), .B1(\us33\/_0221_ ), .C1(\us33\/_0222_ ), .Y(\us33\/_0223_ ) );
sky130_fd_sc_hd__a22o_1 \us33/_1033_ ( .A1(\us33\/_0129_ ), .A2(\us33\/_0162_ ), .B1(\us33\/_0271_ ), .B2(\us33\/_0705_ ), .X(\us33\/_0224_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1034_ ( .A1(\us33\/_0093_ ), .A2(\us33\/_0738_ ), .B1(\us33\/_0081_ ), .C1(\us33\/_0224_ ), .Y(\us33\/_0225_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1035_ ( .A(\us33\/_0214_ ), .B(\us33\/_0220_ ), .C(\us33\/_0223_ ), .D(\us33\/_0225_ ), .X(\us33\/_0226_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1036_ ( .A(\us33\/_0196_ ), .B(\us33\/_0204_ ), .C(\us33\/_0210_ ), .D(\us33\/_0226_ ), .X(\us33\/_0228_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1037_ ( .A(\us33\/_0111_ ), .B(\us33\/_0554_ ), .X(\us33\/_0229_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1038_ ( .A(\us33\/_0229_ ), .Y(\us33\/_0230_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1039_ ( .A(\us33\/_0111_ ), .B(\us33\/_0129_ ), .Y(\us33\/_0231_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1040_ ( .A(\us33\/_0017_ ), .B(\us33\/_0738_ ), .Y(\us33\/_0232_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1041_ ( .A(\us33\/_0030_ ), .B(\us33\/_0304_ ), .Y(\us33\/_0233_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1042_ ( .A(\us33\/_0230_ ), .B(\us33\/_0231_ ), .C(\us33\/_0232_ ), .D(\us33\/_0233_ ), .X(\us33\/_0234_ ) );
sky130_fd_sc_hd__and2_1 \us33/_1043_ ( .A(\us33\/_0047_ ), .B(\us33\/_0478_ ), .X(\us33\/_0235_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1044_ ( .A1(\us33\/_0129_ ), .A2(\us33\/_0554_ ), .B1(\us33\/_0137_ ), .Y(\us33\/_0236_ ) );
sky130_fd_sc_hd__nor3b_1 \us33/_1045_ ( .A(\us33\/_0235_ ), .B(\us33\/_0049_ ), .C_N(\us33\/_0236_ ), .Y(\us33\/_0237_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1046_ ( .A(\us33\/_0047_ ), .B(\us33\/_0077_ ), .X(\us33\/_0239_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1047_ ( .A(\us33\/_0070_ ), .B(\us33\/_0035_ ), .X(\us33\/_0240_ ) );
sky130_fd_sc_hd__a22o_1 \us33/_1048_ ( .A1(\us33\/_0047_ ), .A2(\us33\/_0736_ ), .B1(\us33\/_0022_ ), .B2(\us33\/_0099_ ), .X(\us33\/_0241_ ) );
sky130_fd_sc_hd__nor3_1 \us33/_1049_ ( .A(\us33\/_0239_ ), .B(\us33\/_0240_ ), .C(\us33\/_0241_ ), .Y(\us33\/_0242_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1050_ ( .A(\us33\/_0554_ ), .B(\us33\/_0072_ ), .X(\us33\/_0243_ ) );
sky130_fd_sc_hd__a22o_1 \us33/_1051_ ( .A1(\us33\/_0142_ ), .A2(\us33\/_0137_ ), .B1(\us33\/_0159_ ), .B2(\us33\/_0082_ ), .X(\us33\/_0244_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1052_ ( .A1(\us33\/_0608_ ), .A2(\us33\/_0072_ ), .B1(\us33\/_0243_ ), .C1(\us33\/_0244_ ), .Y(\us33\/_0245_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1053_ ( .A(\us33\/_0234_ ), .B(\us33\/_0237_ ), .C(\us33\/_0242_ ), .D(\us33\/_0245_ ), .X(\us33\/_0246_ ) );
sky130_fd_sc_hd__buf_2 \us33/_1054_ ( .A(\us33\/_0027_ ), .X(\us33\/_0247_ ) );
sky130_fd_sc_hd__o21a_1 \us33/_1055_ ( .A1(\us33\/_0554_ ), .A2(\us33\/_0586_ ), .B1(\us33\/_0247_ ), .X(\us33\/_0248_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1056_ ( .A(\us33\/_0082_ ), .B(\us33\/_0478_ ), .X(\us33\/_0250_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_1057_ ( .A(\us33\/_0079_ ), .X(\us33\/_0251_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1058_ ( .A(\us33\/_0251_ ), .B(\us33\/_0478_ ), .X(\us33\/_0252_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_1059_ ( .A(\us33\/_0250_ ), .B(\us33\/_0252_ ), .Y(\us33\/_0253_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1060_ ( .A(\us33\/_0016_ ), .B(\us33\/_0064_ ), .Y(\us33\/_0254_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_1061_ ( .A(\us33\/_0304_ ), .X(\us33\/_0255_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1062_ ( .A(\us33\/_0255_ ), .B(\us33\/_0640_ ), .Y(\us33\/_0256_ ) );
sky130_fd_sc_hd__and4b_1 \us33/_1063_ ( .A_N(\us33\/_0248_ ), .B(\us33\/_0253_ ), .C(\us33\/_0254_ ), .D(\us33\/_0256_ ), .X(\us33\/_0257_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1064_ ( .A(\us33\/_0099_ ), .B(\us33\/_0110_ ), .X(\us33\/_0258_ ) );
sky130_fd_sc_hd__a21oi_1 \us33/_1065_ ( .A1(\us33\/_0161_ ), .A2(\us33\/_0130_ ), .B1(\us33\/_0258_ ), .Y(\us33\/_0259_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1066_ ( .A(\us33\/_0194_ ), .B(\sa33\[1\] ), .X(\us33\/_0261_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1068_ ( .A(\us33\/_0261_ ), .B(\us33\/_0153_ ), .Y(\us33\/_0263_ ) );
sky130_fd_sc_hd__and3b_1 \us33/_1069_ ( .A_N(\us33\/_0154_ ), .B(\us33\/_0259_ ), .C(\us33\/_0263_ ), .X(\us33\/_0264_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1070_ ( .A(\us33\/_0246_ ), .B(\us33\/_0174_ ), .C(\us33\/_0257_ ), .D(\us33\/_0264_ ), .X(\us33\/_0265_ ) );
sky130_fd_sc_hd__o21a_1 \us33/_1071_ ( .A1(\us33\/_0261_ ), .A2(\us33\/_0554_ ), .B1(\us33\/_0159_ ), .X(\us33\/_0266_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1072_ ( .A(\us33\/_0746_ ), .B(\us33\/_0150_ ), .Y(\us33\/_0267_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1073_ ( .A(\us33\/_0175_ ), .Y(\us33\/_0268_ ) );
sky130_fd_sc_hd__and3_1 \us33/_1074_ ( .A(\us33\/_0412_ ), .B(\us33\/_0123_ ), .C(\us33\/_0151_ ), .X(\us33\/_0269_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1075_ ( .A(\us33\/_0268_ ), .B(\us33\/_0269_ ), .Y(\us33\/_0270_ ) );
sky130_fd_sc_hd__and3b_1 \us33/_1076_ ( .A_N(\us33\/_0266_ ), .B(\us33\/_0267_ ), .C(\us33\/_0270_ ), .X(\us33\/_0272_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1077_ ( .A(\us33\/_0554_ ), .B(\us33\/_0150_ ), .X(\us33\/_0273_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1078_ ( .A(\us33\/_0273_ ), .Y(\us33\/_0274_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1079_ ( .A1(\us33\/_0734_ ), .A2(\us33\/_0325_ ), .B1(\us33\/_0380_ ), .Y(\us33\/_0275_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1080_ ( .A(\us33\/_0275_ ), .Y(\us33\/_0276_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1081_ ( .A(\us33\/_0276_ ), .B(\us33\/_0153_ ), .Y(\us33\/_0277_ ) );
sky130_fd_sc_hd__and3_1 \us33/_1082_ ( .A(\us33\/_0272_ ), .B(\us33\/_0274_ ), .C(\us33\/_0277_ ), .X(\us33\/_0278_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_1083_ ( .A(\us33\/_0035_ ), .X(\us33\/_0279_ ) );
sky130_fd_sc_hd__buf_2 \us33/_1084_ ( .A(\us33\/_0082_ ), .X(\us33\/_0280_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1085_ ( .A1(\us33\/_0499_ ), .A2(\us33\/_0279_ ), .B1(\us33\/_0280_ ), .B2(\us33\/_0060_ ), .Y(\us33\/_0281_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1086_ ( .A1(\us33\/_0251_ ), .A2(\us33\/_0434_ ), .B1(\us33\/_0304_ ), .Y(\us33\/_0283_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1087_ ( .A(\us33\/_0091_ ), .B(\us33\/_0292_ ), .Y(\us33\/_0284_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1088_ ( .A1(\us33\/_0118_ ), .A2(\us33\/_0050_ ), .B1(\us33\/_0038_ ), .C1(\us33\/_0255_ ), .Y(\us33\/_0285_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1089_ ( .A(\us33\/_0281_ ), .B(\us33\/_0283_ ), .C(\us33\/_0284_ ), .D(\us33\/_0285_ ), .X(\us33\/_0286_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1090_ ( .A(\us33\/_0082_ ), .B(\us33\/_0027_ ), .X(\us33\/_0287_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1091_ ( .A(\us33\/_0129_ ), .B(\us33\/_0027_ ), .X(\us33\/_0288_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_1092_ ( .A(\us33\/_0287_ ), .B(\us33\/_0288_ ), .Y(\us33\/_0289_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1093_ ( .A1(\us33\/_0752_ ), .A2(\us33\/_0683_ ), .B1(\us33\/_0093_ ), .B2(\us33\/_0247_ ), .Y(\us33\/_0290_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1094_ ( .A1(\us33\/_0092_ ), .A2(\us33\/_0575_ ), .B1(\us33\/_0292_ ), .Y(\us33\/_0291_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_1095_ ( .A(\us33\/_0054_ ), .X(\us33\/_0292_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1096_ ( .A1(\us33\/_0499_ ), .A2(\us33\/_0662_ ), .B1(\us33\/_0280_ ), .B2(\us33\/_0292_ ), .Y(\us33\/_0294_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1097_ ( .A(\us33\/_0289_ ), .B(\us33\/_0290_ ), .C(\us33\/_0291_ ), .D(\us33\/_0294_ ), .X(\us33\/_0295_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1098_ ( .A(\us33\/_0750_ ), .B(\us33\/_0193_ ), .X(\us33\/_0296_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1099_ ( .A(\us33\/_0705_ ), .B(\us33\/_0380_ ), .X(\us33\/_0297_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1100_ ( .A(\us33\/_0752_ ), .B(\us33\/_0129_ ), .Y(\us33\/_0298_ ) );
sky130_fd_sc_hd__nor3b_1 \us33/_1101_ ( .A(\us33\/_0296_ ), .B(\us33\/_0297_ ), .C_N(\us33\/_0298_ ), .Y(\us33\/_0299_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1102_ ( .A(\us33\/_0089_ ), .B(\us33\/_0532_ ), .Y(\us33\/_0300_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1103_ ( .A(\sa33\[2\] ), .Y(\us33\/_0301_ ) );
sky130_fd_sc_hd__nor3_1 \us33/_1104_ ( .A(\us33\/_0301_ ), .B(\sa33\[3\] ), .C(\us33\/_0118_ ), .Y(\us33\/_0302_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1105_ ( .A(\us33\/_0072_ ), .B(\us33\/_0302_ ), .X(\us33\/_0303_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1106_ ( .A(\us33\/_0303_ ), .Y(\us33\/_0305_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1107_ ( .A(\us33\/_0147_ ), .B(\us33\/_0302_ ), .Y(\us33\/_0306_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1108_ ( .A(\us33\/_0299_ ), .B(\us33\/_0300_ ), .C(\us33\/_0305_ ), .D(\us33\/_0306_ ), .X(\us33\/_0307_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1109_ ( .A(\us33\/_0278_ ), .B(\us33\/_0286_ ), .C(\us33\/_0295_ ), .D(\us33\/_0307_ ), .X(\us33\/_0308_ ) );
sky130_fd_sc_hd__nand3_1 \us33/_1110_ ( .A(\us33\/_0228_ ), .B(\us33\/_0265_ ), .C(\us33\/_0308_ ), .Y(\us33\/_0009_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1111_ ( .A(\us33\/_0235_ ), .Y(\us33\/_0309_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1112_ ( .A(\us33\/_0478_ ), .B(\us33\/_0640_ ), .X(\us33\/_0310_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1113_ ( .A(\us33\/_0310_ ), .Y(\us33\/_0311_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1114_ ( .A(\us33\/_0022_ ), .B(\us33\/_0499_ ), .Y(\us33\/_0312_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1115_ ( .A(\us33\/_0499_ ), .B(\us33\/_0032_ ), .Y(\us33\/_0313_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1116_ ( .A(\us33\/_0309_ ), .B(\us33\/_0311_ ), .C(\us33\/_0312_ ), .D(\us33\/_0313_ ), .X(\us33\/_0315_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1117_ ( .A(\us33\/_0499_ ), .B(\us33\/_0064_ ), .Y(\us33\/_0316_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1118_ ( .A(\us33\/_0499_ ), .B(\us33\/_0683_ ), .Y(\us33\/_0317_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1119_ ( .A(\us33\/_0315_ ), .B(\us33\/_0316_ ), .C(\us33\/_0317_ ), .D(\us33\/_0253_ ), .X(\us33\/_0318_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1120_ ( .A(\us33\/_0047_ ), .B(\us33\/_0304_ ), .Y(\us33\/_0319_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1121_ ( .A(\us33\/_0586_ ), .B(\us33\/_0162_ ), .Y(\us33\/_0320_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1122_ ( .A(\us33\/_0319_ ), .B(\us33\/_0320_ ), .Y(\us33\/_0321_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_1123_ ( .A(\us33\/_0321_ ), .B(\us33\/_0238_ ), .Y(\us33\/_0322_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1124_ ( .A(\us33\/_0304_ ), .B(\us33\/_0062_ ), .Y(\us33\/_0323_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_1125_ ( .A(\us33\/_0251_ ), .X(\us33\/_0324_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1126_ ( .A1(\us33\/_0324_ ), .A2(\us33\/_0280_ ), .B1(\us33\/_0255_ ), .Y(\us33\/_0326_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1127_ ( .A1(\us33\/_0050_ ), .A2(\us33\/_0205_ ), .B1(\us33\/_0109_ ), .C1(\us33\/_0255_ ), .Y(\us33\/_0327_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1128_ ( .A(\us33\/_0322_ ), .B(\us33\/_0323_ ), .C(\us33\/_0326_ ), .D(\us33\/_0327_ ), .X(\us33\/_0328_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1129_ ( .A1(\us33\/_0733_ ), .A2(\us33\/_0279_ ), .A3(\us33\/_0058_ ), .B1(\us33\/_0292_ ), .Y(\us33\/_0329_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_1130_ ( .A(\us33\/_0047_ ), .X(\us33\/_0330_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1131_ ( .A(\us33\/_0330_ ), .B(\us33\/_0292_ ), .Y(\us33\/_0331_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1132_ ( .A(\us33\/_0054_ ), .B(\us33\/_0045_ ), .Y(\us33\/_0332_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1133_ ( .A(\us33\/_0329_ ), .B(\us33\/_0331_ ), .C(\us33\/_0284_ ), .D(\us33\/_0332_ ), .X(\us33\/_0333_ ) );
sky130_fd_sc_hd__o211a_1 \us33/_1134_ ( .A1(\us33\/_0249_ ), .A2(\us33\/_0205_ ), .B1(\us33\/_0532_ ), .C1(\us33\/_0060_ ), .X(\us33\/_0334_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1135_ ( .A(\us33\/_0280_ ), .B(\us33\/_0060_ ), .Y(\us33\/_0335_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1136_ ( .A(\us33\/_0324_ ), .B(\us33\/_0060_ ), .Y(\us33\/_0337_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1137_ ( .A(\us33\/_0335_ ), .B(\us33\/_0337_ ), .Y(\us33\/_0338_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1138_ ( .A1(\us33\/_0276_ ), .A2(\us33\/_0060_ ), .B1(\us33\/_0334_ ), .C1(\us33\/_0338_ ), .Y(\us33\/_0339_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1139_ ( .A(\us33\/_0318_ ), .B(\us33\/_0328_ ), .C(\us33\/_0333_ ), .D(\us33\/_0339_ ), .X(\us33\/_0340_ ) );
sky130_fd_sc_hd__o21a_1 \us33/_1140_ ( .A1(\us33\/_0746_ ), .A2(\us33\/_0134_ ), .B1(\us33\/_0128_ ), .X(\us33\/_0341_ ) );
sky130_fd_sc_hd__and2b_1 \us33/_1141_ ( .A_N(\us33\/_0086_ ), .B(\us33\/_0128_ ), .X(\us33\/_0342_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1142_ ( .A(\us33\/_0079_ ), .B(\us33\/_0124_ ), .X(\us33\/_0343_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_1143_ ( .A(\us33\/_0126_ ), .B(\us33\/_0343_ ), .Y(\us33\/_0344_ ) );
sky130_fd_sc_hd__nor3b_1 \us33/_1144_ ( .A(\us33\/_0341_ ), .B(\us33\/_0342_ ), .C_N(\us33\/_0344_ ), .Y(\us33\/_0345_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1146_ ( .A1(\us33\/_0193_ ), .A2(\us33\/_0092_ ), .A3(\us33\/_0330_ ), .B1(\us33\/_0147_ ), .Y(\us33\/_0348_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1147_ ( .A1(\us33\/_0130_ ), .A2(\us33\/_0280_ ), .A3(\us33\/_0134_ ), .B1(\us33\/_0139_ ), .Y(\us33\/_0349_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1148_ ( .A1(\us33\/_0144_ ), .A2(\us33\/_0608_ ), .A3(\us33\/_0092_ ), .B1(\us33\/_0139_ ), .Y(\us33\/_0350_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1149_ ( .A(\us33\/_0345_ ), .B(\us33\/_0348_ ), .C(\us33\/_0349_ ), .D(\us33\/_0350_ ), .X(\us33\/_0351_ ) );
sky130_fd_sc_hd__and3_1 \us33/_1150_ ( .A(\us33\/_0150_ ), .B(\us33\/_0194_ ), .C(\us33\/_0249_ ), .X(\us33\/_0352_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us33/_1151_ ( .A(\us33\/_0277_ ), .SLEEP(\us33\/_0352_ ), .X(\us33\/_0353_ ) );
sky130_fd_sc_hd__a21oi_1 \us33/_1152_ ( .A1(\us33\/_0268_ ), .A2(\us33\/_0171_ ), .B1(\us33\/_0157_ ), .Y(\us33\/_0354_ ) );
sky130_fd_sc_hd__clkbuf_1 \us33/_1153_ ( .A(\us33\/_0161_ ), .X(\us33\/_0355_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1154_ ( .A1(\us33\/_0279_ ), .A2(\us33\/_0280_ ), .B1(\us33\/_0355_ ), .Y(\us33\/_0356_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1155_ ( .A1(\us33\/_0020_ ), .A2(\us33\/_0193_ ), .A3(\us33\/_0091_ ), .B1(\us33\/_0355_ ), .Y(\us33\/_0357_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1156_ ( .A(\us33\/_0353_ ), .B(\us33\/_0354_ ), .C(\us33\/_0356_ ), .D(\us33\/_0357_ ), .X(\us33\/_0359_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1157_ ( .A(\us33\/_0111_ ), .B(\us33\/_0586_ ), .X(\us33\/_0360_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1158_ ( .A(\us33\/_0360_ ), .Y(\us33\/_0361_ ) );
sky130_fd_sc_hd__o211a_1 \us33/_1159_ ( .A1(\us33\/_0119_ ), .A2(\us33\/_0120_ ), .B1(\us33\/_0230_ ), .C1(\us33\/_0361_ ), .X(\us33\/_0362_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1160_ ( .A1(\us33\/_0662_ ), .A2(\us33\/_0251_ ), .A3(\us33\/_0134_ ), .B1(\us33\/_0114_ ), .Y(\us33\/_0363_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1162_ ( .A1(\us33\/_0035_ ), .A2(\us33\/_0251_ ), .A3(\us33\/_0134_ ), .B1(\us33\/_0099_ ), .Y(\us33\/_0365_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1163_ ( .A1(\us33\/_0193_ ), .A2(\us33\/_0608_ ), .B1(\us33\/_0099_ ), .Y(\us33\/_0366_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1164_ ( .A(\us33\/_0362_ ), .B(\us33\/_0363_ ), .C(\us33\/_0365_ ), .D(\us33\/_0366_ ), .X(\us33\/_0367_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1165_ ( .A1(\us33\/_0575_ ), .A2(\us33\/_0092_ ), .A3(\us33\/_0330_ ), .B1(\us33\/_0089_ ), .Y(\us33\/_0368_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1166_ ( .A1(\us33\/_0586_ ), .A2(\us33\/_0017_ ), .A3(\us33\/_0330_ ), .B1(\us33\/_0094_ ), .Y(\us33\/_0370_ ) );
sky130_fd_sc_hd__o21ai_1 \us33/_1167_ ( .A1(\us33\/_0293_ ), .A2(\us33\/_0134_ ), .B1(\us33\/_0089_ ), .Y(\us33\/_0371_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1168_ ( .A1(\us33\/_0279_ ), .A2(\us33\/_0134_ ), .B1(\us33\/_0094_ ), .Y(\us33\/_0372_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1169_ ( .A(\us33\/_0368_ ), .B(\us33\/_0370_ ), .C(\us33\/_0371_ ), .D(\us33\/_0372_ ), .X(\us33\/_0373_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1170_ ( .A(\us33\/_0351_ ), .B(\us33\/_0359_ ), .C(\us33\/_0367_ ), .D(\us33\/_0373_ ), .X(\us33\/_0374_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1171_ ( .A1(\us33\/_0102_ ), .A2(\us33\/_0347_ ), .B1(\us33\/_0109_ ), .C1(\us33\/_0247_ ), .Y(\us33\/_0375_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1172_ ( .A1(\us33\/_0102_ ), .A2(\us33\/_0347_ ), .B1(\us33\/_0532_ ), .C1(\us33\/_0247_ ), .Y(\us33\/_0376_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1173_ ( .A1(\us33\/_0050_ ), .A2(\us33\/_0249_ ), .B1(\us33\/_0380_ ), .C1(\us33\/_0247_ ), .Y(\us33\/_0377_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1174_ ( .A(\us33\/_0041_ ), .B(\us33\/_0375_ ), .C(\us33\/_0376_ ), .D(\us33\/_0377_ ), .X(\us33\/_0378_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1175_ ( .A(\us33\/_0047_ ), .B(\us33\/_0750_ ), .X(\us33\/_0379_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1176_ ( .A(\us33\/_0379_ ), .Y(\us33\/_0381_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1177_ ( .A(\us33\/_0016_ ), .B(\us33\/_0608_ ), .Y(\us33\/_0382_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1178_ ( .A(\us33\/_0752_ ), .B(\us33\/_0554_ ), .Y(\us33\/_0383_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1179_ ( .A1(\sa33\[1\] ), .A2(\us33\/_0734_ ), .B1(\us33\/_0109_ ), .C1(\us33\/_0016_ ), .Y(\us33\/_0384_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1180_ ( .A(\us33\/_0381_ ), .B(\us33\/_0382_ ), .C(\us33\/_0383_ ), .D(\us33\/_0384_ ), .X(\us33\/_0385_ ) );
sky130_fd_sc_hd__or2b_1 \us33/_1181_ ( .A(\us33\/_0086_ ), .B_N(\us33\/_0736_ ), .X(\us33\/_0386_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1182_ ( .A1(\us33\/_0748_ ), .A2(\us33\/_0134_ ), .B1(\us33\/_0739_ ), .Y(\us33\/_0387_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1183_ ( .A1(\us33\/_0118_ ), .A2(\us33\/_0249_ ), .B1(\us33\/_0109_ ), .C1(\us33\/_0739_ ), .Y(\us33\/_0388_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1184_ ( .A1(\us33\/_0102_ ), .A2(\us33\/_0301_ ), .B1(\sa33\[3\] ), .C1(\us33\/_0739_ ), .Y(\us33\/_0389_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1185_ ( .A(\us33\/_0386_ ), .B(\us33\/_0387_ ), .C(\us33\/_0388_ ), .D(\us33\/_0389_ ), .X(\us33\/_0390_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1186_ ( .A(\us33\/_0020_ ), .Y(\us33\/_0392_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1187_ ( .A(\us33\/_0727_ ), .Y(\us33\/_0393_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1188_ ( .A(\us33\/_0727_ ), .B(\us33\/_0064_ ), .Y(\us33\/_0394_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1189_ ( .A1(\us33\/_0102_ ), .A2(\us33\/_0734_ ), .B1(\us33\/_0532_ ), .C1(\us33\/_0727_ ), .Y(\us33\/_0395_ ) );
sky130_fd_sc_hd__o211a_1 \us33/_1190_ ( .A1(\us33\/_0392_ ), .A2(\us33\/_0393_ ), .B1(\us33\/_0394_ ), .C1(\us33\/_0395_ ), .X(\us33\/_0396_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1191_ ( .A(\us33\/_0378_ ), .B(\us33\/_0385_ ), .C(\us33\/_0390_ ), .D(\us33\/_0396_ ), .X(\us33\/_0397_ ) );
sky130_fd_sc_hd__nand3_1 \us33/_1192_ ( .A(\us33\/_0340_ ), .B(\us33\/_0374_ ), .C(\us33\/_0397_ ), .Y(\us33\/_0010_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1193_ ( .A(\us33\/_0077_ ), .B(\us33\/_0129_ ), .X(\us33\/_0398_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_1194_ ( .A(\us33\/_0398_ ), .B(\us33\/_0239_ ), .Y(\us33\/_0399_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1195_ ( .A(\us33\/_0022_ ), .B(\us33\/_0111_ ), .X(\us33\/_0400_ ) );
sky130_fd_sc_hd__nand2b_1 \us33/_1196_ ( .A_N(\us33\/_0400_ ), .B(\us33\/_0231_ ), .Y(\us33\/_0402_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us33/_1197_ ( .A(\us33\/_0399_ ), .SLEEP(\us33\/_0402_ ), .X(\us33\/_0403_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_1198_ ( .A(\us33\/_0746_ ), .B(\us33\/_0251_ ), .Y(\us33\/_0404_ ) );
sky130_fd_sc_hd__nand2b_1 \us33/_1199_ ( .A_N(\us33\/_0404_ ), .B(\us33\/_0752_ ), .Y(\us33\/_0405_ ) );
sky130_fd_sc_hd__and3_1 \us33/_1200_ ( .A(\us33\/_0467_ ), .B(\us33\/_0194_ ), .C(\us33\/_0694_ ), .X(\us33\/_0406_ ) );
sky130_fd_sc_hd__and2b_1 \us33/_1201_ ( .A_N(\us33\/_0175_ ), .B(\us33\/_0406_ ), .X(\us33\/_0407_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1202_ ( .A(\us33\/_0407_ ), .Y(\us33\/_0408_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1203_ ( .A1(\us33\/_0094_ ), .A2(\us33\/_0197_ ), .B1(\us33\/_0114_ ), .B2(\us33\/_0640_ ), .Y(\us33\/_0409_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1204_ ( .A(\us33\/_0403_ ), .B(\us33\/_0405_ ), .C(\us33\/_0408_ ), .D(\us33\/_0409_ ), .X(\us33\/_0410_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1205_ ( .A(\us33\/_0030_ ), .B(\us33\/_0150_ ), .Y(\us33\/_0411_ ) );
sky130_fd_sc_hd__and3b_1 \us33/_1206_ ( .A_N(\us33\/_0169_ ), .B(\us33\/_0289_ ), .C(\us33\/_0411_ ), .X(\us33\/_0413_ ) );
sky130_fd_sc_hd__o211a_1 \us33/_1207_ ( .A1(\us33\/_0467_ ), .A2(\us33\/_0151_ ), .B1(\us33\/_0140_ ), .C1(\us33\/_0129_ ), .X(\us33\/_0414_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1208_ ( .A1(\us33\/_0608_ ), .A2(\us33\/_0099_ ), .B1(\us33\/_0037_ ), .C1(\us33\/_0414_ ), .Y(\us33\/_0415_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1209_ ( .A(\us33\/_0738_ ), .Y(\us33\/_0416_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1210_ ( .A(\us33\/_0586_ ), .B(\us33\/_0736_ ), .Y(\us33\/_0417_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1211_ ( .A1(\us33\/_0194_ ), .A2(\us33\/_0038_ ), .B1(\us33\/_0118_ ), .C1(\us33\/_0153_ ), .Y(\us33\/_0418_ ) );
sky130_fd_sc_hd__o211a_1 \us33/_1212_ ( .A1(\us33\/_0416_ ), .A2(\us33\/_0117_ ), .B1(\us33\/_0417_ ), .C1(\us33\/_0418_ ), .X(\us33\/_0419_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1213_ ( .A(\us33\/_0077_ ), .B(\us33\/_0035_ ), .X(\us33\/_0420_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1214_ ( .A(\us33\/_0662_ ), .B(\us33\/_0124_ ), .Y(\us33\/_0421_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1215_ ( .A(\us33\/_0030_ ), .B(\us33\/_0137_ ), .Y(\us33\/_0422_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1216_ ( .A(\us33\/_0072_ ), .B(\us33\/_0731_ ), .Y(\us33\/_0424_ ) );
sky130_fd_sc_hd__and4b_1 \us33/_1217_ ( .A_N(\us33\/_0420_ ), .B(\us33\/_0421_ ), .C(\us33\/_0422_ ), .D(\us33\/_0424_ ), .X(\us33\/_0425_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1218_ ( .A(\us33\/_0413_ ), .B(\us33\/_0415_ ), .C(\us33\/_0419_ ), .D(\us33\/_0425_ ), .X(\us33\/_0426_ ) );
sky130_fd_sc_hd__nand3_1 \us33/_1219_ ( .A(\us33\/_0355_ ), .B(\us33\/_0102_ ), .C(\us33\/_0109_ ), .Y(\us33\/_0427_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1220_ ( .A(\us33\/_0077_ ), .B(\us33\/_0017_ ), .X(\us33\/_0428_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1221_ ( .A(\us33\/_0077_ ), .B(\us33\/_0554_ ), .X(\us33\/_0429_ ) );
sky130_fd_sc_hd__o211a_1 \us33/_1222_ ( .A1(\us33\/_0050_ ), .A2(\us33\/_0205_ ), .B1(\us33\/_0380_ ), .C1(\us33\/_0078_ ), .X(\us33\/_0430_ ) );
sky130_fd_sc_hd__nor3_1 \us33/_1223_ ( .A(\us33\/_0428_ ), .B(\us33\/_0429_ ), .C(\us33\/_0430_ ), .Y(\us33\/_0431_ ) );
sky130_fd_sc_hd__and2b_1 \us33/_1224_ ( .A_N(\us33\/_0209_ ), .B(\us33\/_0431_ ), .X(\us33\/_0432_ ) );
sky130_fd_sc_hd__o211a_1 \us33/_1225_ ( .A1(\us33\/_0215_ ), .A2(\us33\/_0404_ ), .B1(\us33\/_0427_ ), .C1(\us33\/_0432_ ), .X(\us33\/_0433_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1226_ ( .A(\us33\/_0043_ ), .B(\us33\/_0058_ ), .Y(\us33\/_0435_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1227_ ( .A(\us33\/_0195_ ), .B(\us33\/_0233_ ), .C(\us33\/_0320_ ), .D(\us33\/_0435_ ), .X(\us33\/_0436_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1228_ ( .A(\us33\/_0261_ ), .B(\us33\/_0738_ ), .Y(\us33\/_0437_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1229_ ( .A1(\us33\/_0499_ ), .A2(\us33\/_0640_ ), .B1(\us33\/_0261_ ), .B2(\us33\/_0292_ ), .Y(\us33\/_0438_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1230_ ( .A(\us33\/_0436_ ), .B(\us33\/_0394_ ), .C(\us33\/_0437_ ), .D(\us33\/_0438_ ), .X(\us33\/_0439_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1231_ ( .A(\us33\/_0410_ ), .B(\us33\/_0426_ ), .C(\us33\/_0433_ ), .D(\us33\/_0439_ ), .X(\us33\/_0440_ ) );
sky130_fd_sc_hd__lpflow_isobufsrc_1 \us33/_1232_ ( .A(\us33\/_0135_ ), .SLEEP(\us33\/_0273_ ), .X(\us33\/_0441_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1233_ ( .A1(\us33\/_0279_ ), .A2(\us33\/_0134_ ), .B1(\us33\/_0099_ ), .Y(\us33\/_0442_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1234_ ( .A(\us33\/_0441_ ), .B(\us33\/_0164_ ), .C(\us33\/_0270_ ), .D(\us33\/_0442_ ), .X(\us33\/_0443_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1235_ ( .A(\us33\/_0051_ ), .B(\us33\/_0662_ ), .Y(\us33\/_0444_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1236_ ( .A(\us33\/_0051_ ), .B(\us33\/_0271_ ), .Y(\us33\/_0446_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1237_ ( .A(\us33\/_0444_ ), .B(\us33\/_0446_ ), .X(\us33\/_0447_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1238_ ( .A(\us33\/_0193_ ), .B(\us33\/_0304_ ), .X(\us33\/_0448_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1239_ ( .A(\us33\/_0448_ ), .Y(\us33\/_0449_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1240_ ( .A(\us33\/_0162_ ), .B(\us33\/_0130_ ), .X(\us33\/_0450_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1241_ ( .A(\us33\/_0450_ ), .Y(\us33\/_0451_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1242_ ( .A1(\us33\/_0129_ ), .A2(\us33\/_0554_ ), .B1(\us33\/_0043_ ), .Y(\us33\/_0452_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1243_ ( .A(\us33\/_0447_ ), .B(\us33\/_0449_ ), .C(\us33\/_0451_ ), .D(\us33\/_0452_ ), .X(\us33\/_0453_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1244_ ( .A(\us33\/_0292_ ), .B(\us33\/_0064_ ), .Y(\us33\/_0454_ ) );
sky130_fd_sc_hd__and4b_1 \us33/_1245_ ( .A_N(\us33\/_0248_ ), .B(\us33\/_0454_ ), .C(\us33\/_0254_ ), .D(\us33\/_0256_ ), .X(\us33\/_0455_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1246_ ( .A1(\us33\/_0330_ ), .A2(\us33\/_0099_ ), .B1(\us33\/_0134_ ), .B2(\us33\/_0705_ ), .Y(\us33\/_0457_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1247_ ( .A1(\us33\/_0748_ ), .A2(\us33\/_0738_ ), .B1(\us33\/_0092_ ), .B2(\us33\/_0752_ ), .Y(\us33\/_0458_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1248_ ( .A1(\us33\/_0072_ ), .A2(\us33\/_0035_ ), .B1(\us33\/_0748_ ), .B2(\us33\/_0292_ ), .Y(\us33\/_0459_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1249_ ( .A1(\us33\/_0748_ ), .A2(\us33\/_0251_ ), .B1(\us33\/_0247_ ), .Y(\us33\/_0460_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1250_ ( .A(\us33\/_0457_ ), .B(\us33\/_0458_ ), .C(\us33\/_0459_ ), .D(\us33\/_0460_ ), .X(\us33\/_0461_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1251_ ( .A(\us33\/_0443_ ), .B(\us33\/_0453_ ), .C(\us33\/_0455_ ), .D(\us33\/_0461_ ), .X(\us33\/_0462_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1252_ ( .A(\us33\/_0705_ ), .B(\us33\/_0079_ ), .X(\us33\/_0463_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1253_ ( .A(\us33\/_0586_ ), .B(\us33\/_0124_ ), .Y(\us33\/_0464_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1254_ ( .A(\us33\/_0499_ ), .B(\us33\/_0746_ ), .Y(\us33\/_0465_ ) );
sky130_fd_sc_hd__and3b_1 \us33/_1255_ ( .A_N(\us33\/_0463_ ), .B(\us33\/_0464_ ), .C(\us33\/_0465_ ), .X(\us33\/_0466_ ) );
sky130_fd_sc_hd__a22o_1 \us33/_1256_ ( .A1(\us33\/_0271_ ), .A2(\us33\/_0072_ ), .B1(\us33\/_0142_ ), .B2(\us33\/_0027_ ), .X(\us33\/_0468_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1257_ ( .A1(\us33\/_0144_ ), .A2(\us33\/_0099_ ), .B1(\us33\/_0360_ ), .C1(\us33\/_0468_ ), .Y(\us33\/_0469_ ) );
sky130_fd_sc_hd__o21a_1 \us33/_1258_ ( .A1(\us33\/_0662_ ), .A2(\us33\/_0251_ ), .B1(\us33\/_0499_ ), .X(\us33\/_0470_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1259_ ( .A1(\us33\/_0575_ ), .A2(\us33\/_0292_ ), .B1(\us33\/_0379_ ), .C1(\us33\/_0470_ ), .Y(\us33\/_0471_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1260_ ( .A(\us33\/_0466_ ), .B(\us33\/_0469_ ), .C(\us33\/_0471_ ), .D(\us33\/_0305_ ), .X(\us33\/_0472_ ) );
sky130_fd_sc_hd__a22o_1 \us33/_1261_ ( .A1(\us33\/_0247_ ), .A2(\us33\/_0683_ ), .B1(\us33\/_0324_ ), .B2(\us33\/_0292_ ), .X(\us33\/_0473_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1262_ ( .A(\us33\/_0280_ ), .B(\us33\/_0099_ ), .X(\us33\/_0474_ ) );
sky130_fd_sc_hd__a21o_1 \us33/_1263_ ( .A1(\us33\/_0092_ ), .A2(\us33\/_0247_ ), .B1(\us33\/_0474_ ), .X(\us33\/_0475_ ) );
sky130_fd_sc_hd__nor3_1 \us33/_1264_ ( .A(\us33\/_0075_ ), .B(\us33\/_0473_ ), .C(\us33\/_0475_ ), .Y(\us33\/_0476_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1265_ ( .A1(\us33\/_0279_ ), .A2(\us33\/_0255_ ), .B1(\us33\/_0280_ ), .B2(\us33\/_0060_ ), .Y(\us33\/_0477_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1266_ ( .A1(\us33\/_0093_ ), .A2(\us33\/_0292_ ), .B1(\us33\/_0134_ ), .B2(\us33\/_0114_ ), .Y(\us33\/_0479_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1267_ ( .A1(\us33\/_0161_ ), .A2(\us33\/_0032_ ), .B1(\us33\/_0324_ ), .B2(\us33\/_0147_ ), .Y(\us33\/_0480_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1268_ ( .A1(\us33\/_0054_ ), .A2(\us33\/_0731_ ), .B1(\us33\/_0748_ ), .B2(\us33\/_0304_ ), .Y(\us33\/_0481_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1269_ ( .A(\us33\/_0477_ ), .B(\us33\/_0479_ ), .C(\us33\/_0480_ ), .D(\us33\/_0481_ ), .X(\us33\/_0482_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1270_ ( .A(\us33\/_0161_ ), .B(\us33\/_0064_ ), .Y(\us33\/_0483_ ) );
sky130_fd_sc_hd__nand3_1 \us33/_1271_ ( .A(\us33\/_0731_ ), .B(\us33\/_0123_ ), .C(\us33\/_0467_ ), .Y(\us33\/_0484_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1272_ ( .A(\us33\/_0483_ ), .B(\us33\/_0484_ ), .Y(\us33\/_0485_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1273_ ( .A(\us33\/_0297_ ), .Y(\us33\/_0486_ ) );
sky130_fd_sc_hd__and4b_1 \us33/_1274_ ( .A_N(\us33\/_0485_ ), .B(\us33\/_0181_ ), .C(\us33\/_0486_ ), .D(\us33\/_0386_ ), .X(\us33\/_0487_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1275_ ( .A(\us33\/_0472_ ), .B(\us33\/_0476_ ), .C(\us33\/_0482_ ), .D(\us33\/_0487_ ), .X(\us33\/_0488_ ) );
sky130_fd_sc_hd__nand3_1 \us33/_1276_ ( .A(\us33\/_0440_ ), .B(\us33\/_0462_ ), .C(\us33\/_0488_ ), .Y(\us33\/_0011_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1277_ ( .A(\us33\/_0403_ ), .B(\us33\/_0230_ ), .C(\us33\/_0451_ ), .D(\us33\/_0361_ ), .X(\us33\/_0490_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1278_ ( .A1(\us33\/_0118_ ), .A2(\us33\/_0050_ ), .B1(\us33\/_0109_ ), .C1(\us33\/_0139_ ), .Y(\us33\/_0491_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1279_ ( .A(\us33\/_0447_ ), .B(\us33\/_0437_ ), .C(\us33\/_0491_ ), .D(\us33\/_0427_ ), .X(\us33\/_0492_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1280_ ( .A1(\us33\/_0280_ ), .A2(\us33\/_0255_ ), .B1(\us33\/_0608_ ), .B2(\us33\/_0247_ ), .Y(\us33\/_0493_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1281_ ( .A1(\us33\/_0144_ ), .A2(\us33\/_0147_ ), .B1(\us33\/_0355_ ), .B2(\us33\/_0093_ ), .Y(\us33\/_0494_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1282_ ( .A1(\us33\/_0705_ ), .A2(\us33\/_0279_ ), .B1(\us33\/_0330_ ), .B2(\us33\/_0247_ ), .Y(\us33\/_0495_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1283_ ( .A1(\us33\/_0279_ ), .A2(\us33\/_0280_ ), .B1(\us33\/_0114_ ), .Y(\us33\/_0496_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1284_ ( .A(\us33\/_0493_ ), .B(\us33\/_0494_ ), .C(\us33\/_0495_ ), .D(\us33\/_0496_ ), .X(\us33\/_0497_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1285_ ( .A1(\us33\/_0134_ ), .A2(\us33\/_0137_ ), .B1(\us33\/_0355_ ), .B2(\us33\/_0575_ ), .Y(\us33\/_0498_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1286_ ( .A1(\us33\/_0099_ ), .A2(\us33\/_0733_ ), .B1(\us33\/_0093_ ), .B2(\us33\/_0499_ ), .Y(\us33\/_0500_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1287_ ( .A(\us33\/_0147_ ), .B(\us33\/_0640_ ), .Y(\us33\/_0501_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1288_ ( .A1(\us33\/_0153_ ), .A2(\us33\/_0292_ ), .B1(\us33\/_0748_ ), .Y(\us33\/_0502_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1289_ ( .A(\us33\/_0498_ ), .B(\us33\/_0500_ ), .C(\us33\/_0501_ ), .D(\us33\/_0502_ ), .X(\us33\/_0503_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1290_ ( .A(\us33\/_0490_ ), .B(\us33\/_0492_ ), .C(\us33\/_0497_ ), .D(\us33\/_0503_ ), .X(\us33\/_0504_ ) );
sky130_fd_sc_hd__and2b_1 \us33/_1291_ ( .A_N(\us33\/_0275_ ), .B(\us33\/_0705_ ), .X(\us33\/_0505_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1292_ ( .A(\us33\/_0505_ ), .Y(\us33\/_0506_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1293_ ( .A(\us33\/_0380_ ), .B(\us33\/_0347_ ), .X(\us33\/_0507_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1294_ ( .A1(\us33\/_0507_ ), .A2(\us33\/_0093_ ), .B1(\us33\/_0292_ ), .Y(\us33\/_0508_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1295_ ( .A(\us33\/_0322_ ), .B(\us33\/_0277_ ), .C(\us33\/_0506_ ), .D(\us33\/_0508_ ), .X(\us33\/_0509_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1296_ ( .A(\us33\/_0280_ ), .B(\us33\/_0705_ ), .X(\us33\/_0511_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1297_ ( .A1(\us33\/_0733_ ), .A2(\us33\/_0114_ ), .B1(\us33\/_0429_ ), .C1(\us33\/_0511_ ), .Y(\us33\/_0512_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_1298_ ( .A(\us33\/_0019_ ), .B(\us33\/_0024_ ), .Y(\us33\/_0513_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1299_ ( .A(\us33\/_0512_ ), .B(\us33\/_0513_ ), .C(\us33\/_0742_ ), .D(\us33\/_0306_ ), .X(\us33\/_0514_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1300_ ( .A1(\us33\/_0532_ ), .A2(\us33\/_0089_ ), .B1(\us33\/_0154_ ), .C1(\us33\/_0169_ ), .Y(\us33\/_0515_ ) );
sky130_fd_sc_hd__o211a_1 \us33/_1301_ ( .A1(\us33\/_0749_ ), .A2(\us33\/_0026_ ), .B1(\us33\/_0069_ ), .C1(\us33\/_0032_ ), .X(\us33\/_0516_ ) );
sky130_fd_sc_hd__a22o_1 \us33/_1302_ ( .A1(\us33\/_0324_ ), .A2(\us33\/_0355_ ), .B1(\us33\/_0330_ ), .B2(\us33\/_0727_ ), .X(\us33\/_0517_ ) );
sky130_fd_sc_hd__nor3_1 \us33/_1303_ ( .A(\us33\/_0133_ ), .B(\us33\/_0516_ ), .C(\us33\/_0517_ ), .Y(\us33\/_0518_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1304_ ( .A(\us33\/_0509_ ), .B(\us33\/_0514_ ), .C(\us33\/_0515_ ), .D(\us33\/_0518_ ), .X(\us33\/_0519_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1305_ ( .A(\us33\/_0746_ ), .B(\us33\/_0072_ ), .Y(\us33\/_0520_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1306_ ( .A1(\us33\/_0082_ ), .A2(\us33\/_0070_ ), .B1(\us33\/_0043_ ), .B2(\us33\/_0193_ ), .Y(\us33\/_0522_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1307_ ( .A(\us33\/_0311_ ), .B(\us33\/_0520_ ), .C(\us33\/_0332_ ), .D(\us33\/_0522_ ), .X(\us33\/_0523_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1308_ ( .A(\us33\/_0129_ ), .B(\us33\/_0499_ ), .X(\us33\/_0524_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_1309_ ( .A(\us33\/_0235_ ), .B(\us33\/_0524_ ), .Y(\us33\/_0525_ ) );
sky130_fd_sc_hd__nor2_1 \us33/_1310_ ( .A(\us33\/_0081_ ), .B(\us33\/_0085_ ), .Y(\us33\/_0526_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1311_ ( .A1(\us33\/_0051_ ), .A2(\us33\/_0045_ ), .B1(\us33\/_0130_ ), .B2(\us33\/_0094_ ), .Y(\us33\/_0527_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1312_ ( .A(\us33\/_0523_ ), .B(\us33\/_0525_ ), .C(\us33\/_0526_ ), .D(\us33\/_0527_ ), .X(\us33\/_0528_ ) );
sky130_fd_sc_hd__nand2b_1 \us33/_1313_ ( .A_N(\us33\/_0250_ ), .B(\us33\/_0521_ ), .Y(\us33\/_0529_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1314_ ( .A(\us33\/_0128_ ), .B(\us33\/_0020_ ), .X(\us33\/_0530_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1315_ ( .A(\us33\/_0530_ ), .Y(\us33\/_0531_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1316_ ( .A(\us33\/_0099_ ), .B(\us33\/_0058_ ), .X(\us33\/_0533_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1317_ ( .A(\us33\/_0533_ ), .Y(\us33\/_0534_ ) );
sky130_fd_sc_hd__and4b_1 \us33/_1318_ ( .A_N(\us33\/_0529_ ), .B(\us33\/_0531_ ), .C(\us33\/_0534_ ), .D(\us33\/_0192_ ), .X(\us33\/_0535_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1319_ ( .A(\us33\/_0434_ ), .B(\us33\/_0078_ ), .X(\us33\/_0536_ ) );
sky130_fd_sc_hd__a22o_1 \us33/_1320_ ( .A1(\us33\/_0750_ ), .A2(\us33\/_0079_ ), .B1(\us33\/_0129_ ), .B2(\us33\/_0705_ ), .X(\us33\/_0537_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1321_ ( .A1(\us33\/_0161_ ), .A2(\us33\/_0032_ ), .B1(\us33\/_0536_ ), .C1(\us33\/_0537_ ), .Y(\us33\/_0538_ ) );
sky130_fd_sc_hd__a22o_1 \us33/_1322_ ( .A1(\us33\/_0746_ ), .A2(\us33\/_0162_ ), .B1(\us33\/_0079_ ), .B2(\us33\/_0043_ ), .X(\us33\/_0539_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1323_ ( .A1(\us33\/_0093_ ), .A2(\us33\/_0247_ ), .B1(\us33\/_0240_ ), .C1(\us33\/_0539_ ), .Y(\us33\/_0540_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1324_ ( .A(\us33\/_0434_ ), .B(\us33\/_0043_ ), .X(\us33\/_0541_ ) );
sky130_fd_sc_hd__a22o_1 \us33/_1325_ ( .A1(\us33\/_0142_ ), .A2(\us33\/_0150_ ), .B1(\us33\/_0022_ ), .B2(\us33\/_0137_ ), .X(\us33\/_0542_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1326_ ( .A1(\us33\/_0279_ ), .A2(\us33\/_0051_ ), .B1(\us33\/_0541_ ), .C1(\us33\/_0542_ ), .Y(\us33\/_0544_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1327_ ( .A(\us33\/_0159_ ), .B(\us33\/_0035_ ), .X(\us33\/_0545_ ) );
sky130_fd_sc_hd__o21a_1 \us33/_1328_ ( .A1(\us33\/_0271_ ), .A2(\us33\/_0434_ ), .B1(\us33\/_0027_ ), .X(\us33\/_0546_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1329_ ( .A1(\us33\/_0091_ ), .A2(\us33\/_0128_ ), .B1(\us33\/_0545_ ), .C1(\us33\/_0546_ ), .Y(\us33\/_0547_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1330_ ( .A(\us33\/_0538_ ), .B(\us33\/_0540_ ), .C(\us33\/_0544_ ), .D(\us33\/_0547_ ), .X(\us33\/_0548_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1331_ ( .A(\us33\/_0099_ ), .B(\us33\/_0193_ ), .X(\us33\/_0549_ ) );
sky130_fd_sc_hd__nor3_1 \us33/_1332_ ( .A(\us33\/_0549_ ), .B(\us33\/_0186_ ), .C(\us33\/_0187_ ), .Y(\us33\/_0550_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1333_ ( .A(\us33\/_0062_ ), .B(\us33\/_0347_ ), .C(\us33\/_0749_ ), .D(\us33\/_0694_ ), .X(\us33\/_0551_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1334_ ( .A1(\us33\/_0130_ ), .A2(\us33\/_0499_ ), .B1(\us33\/_0551_ ), .C1(\us33\/_0101_ ), .Y(\us33\/_0552_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1335_ ( .A(\us33\/_0139_ ), .B(\us33\/_0640_ ), .Y(\us33\/_0553_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1336_ ( .A1(\us33\/_0752_ ), .A2(\us33\/_0662_ ), .B1(\us33\/_0280_ ), .B2(\us33\/_0099_ ), .Y(\us33\/_0555_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1337_ ( .A(\us33\/_0550_ ), .B(\us33\/_0552_ ), .C(\us33\/_0553_ ), .D(\us33\/_0555_ ), .X(\us33\/_0556_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1338_ ( .A(\us33\/_0528_ ), .B(\us33\/_0535_ ), .C(\us33\/_0548_ ), .D(\us33\/_0556_ ), .X(\us33\/_0557_ ) );
sky130_fd_sc_hd__nand3_1 \us33/_1339_ ( .A(\us33\/_0504_ ), .B(\us33\/_0519_ ), .C(\us33\/_0557_ ), .Y(\us33\/_0012_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1340_ ( .A(\us33\/_0054_ ), .B(\us33\/_0507_ ), .X(\us33\/_0558_ ) );
sky130_fd_sc_hd__and4b_1 \us33/_1341_ ( .A_N(\us33\/_0558_ ), .B(\us33\/_0408_ ), .C(\us33\/_0451_ ), .D(\us33\/_0452_ ), .X(\us33\/_0559_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1342_ ( .A(\us33\/_0549_ ), .Y(\us33\/_0560_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1343_ ( .A(\us33\/_0559_ ), .B(\us33\/_0403_ ), .C(\us33\/_0560_ ), .D(\us33\/_0371_ ), .X(\us33\/_0561_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1344_ ( .A(\us33\/_0181_ ), .B(\us33\/_0178_ ), .X(\us33\/_0562_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1345_ ( .A(\us33\/_0562_ ), .B(\us33\/_0552_ ), .C(\us33\/_0553_ ), .D(\us33\/_0555_ ), .X(\us33\/_0563_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1346_ ( .A(\us33\/_0247_ ), .B(\us33\/_0020_ ), .Y(\us33\/_0565_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1347_ ( .A(\us33\/_0051_ ), .B(\us33\/_0130_ ), .X(\us33\/_0566_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1348_ ( .A(\us33\/_0566_ ), .Y(\us33\/_0567_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1349_ ( .A(\us33\/_0159_ ), .B(\us33\/_0412_ ), .X(\us33\/_0568_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1350_ ( .A1(\us33\/_0752_ ), .A2(\us33\/_0640_ ), .B1(\us33\/_0568_ ), .B2(\us33\/_0175_ ), .Y(\us33\/_0569_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1351_ ( .A(\us33\/_0076_ ), .B(\us33\/_0565_ ), .C(\us33\/_0567_ ), .D(\us33\/_0569_ ), .X(\us33\/_0570_ ) );
sky130_fd_sc_hd__o21a_1 \us33/_1352_ ( .A1(\us33\/_0035_ ), .A2(\us33\/_0142_ ), .B1(\us33\/_0161_ ), .X(\us33\/_0571_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1353_ ( .A(\us33\/_0099_ ), .B(\us33\/_0662_ ), .Y(\us33\/_0572_ ) );
sky130_fd_sc_hd__nor3b_1 \us33/_1354_ ( .A(\us33\/_0420_ ), .B(\us33\/_0571_ ), .C_N(\us33\/_0572_ ), .Y(\us33\/_0573_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1355_ ( .A(\us33\/_0051_ ), .B(\us33\/_0746_ ), .Y(\us33\/_0574_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1356_ ( .A(\us33\/_0574_ ), .B(\us33\/_0319_ ), .C(\us33\/_0320_ ), .D(\us33\/_0411_ ), .X(\us33\/_0576_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1357_ ( .A(\us33\/_0736_ ), .B(\us33\/_0035_ ), .Y(\us33\/_0577_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1358_ ( .A(\us33\/_0736_ ), .B(\us33\/_0030_ ), .Y(\us33\/_0578_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1359_ ( .A(\us33\/_0298_ ), .B(\us33\/_0208_ ), .C(\us33\/_0577_ ), .D(\us33\/_0578_ ), .X(\us33\/_0579_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1360_ ( .A1(\us33\/_0020_ ), .A2(\us33\/_0137_ ), .B1(\us33\/_0261_ ), .B2(\us33\/_0128_ ), .Y(\us33\/_0580_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1361_ ( .A(\us33\/_0573_ ), .B(\us33\/_0576_ ), .C(\us33\/_0579_ ), .D(\us33\/_0580_ ), .X(\us33\/_0581_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1362_ ( .A(\us33\/_0561_ ), .B(\us33\/_0563_ ), .C(\us33\/_0570_ ), .D(\us33\/_0581_ ), .X(\us33\/_0582_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1363_ ( .A(\us33\/_0128_ ), .B(\us33\/_0193_ ), .X(\us33\/_0583_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1364_ ( .A(\us33\/_0082_ ), .B(\us33\/_0162_ ), .X(\us33\/_0584_ ) );
sky130_fd_sc_hd__nor3b_1 \us33/_1365_ ( .A(\us33\/_0583_ ), .B(\us33\/_0584_ ), .C_N(\us33\/_0437_ ), .Y(\us33\/_0585_ ) );
sky130_fd_sc_hd__nand3_1 \us33/_1366_ ( .A(\us33\/_0150_ ), .B(\us33\/_0118_ ), .C(\us33\/_0380_ ), .Y(\us33\/_0587_ ) );
sky130_fd_sc_hd__and3b_1 \us33/_1367_ ( .A_N(\us33\/_0182_ ), .B(\us33\/_0587_ ), .C(\us33\/_0323_ ), .X(\us33\/_0588_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1368_ ( .A1(\us33\/_0575_ ), .A2(\us33\/_0153_ ), .B1(\us33\/_0727_ ), .B2(\us33\/_0058_ ), .Y(\us33\/_0589_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1369_ ( .A1(\us33\/_0499_ ), .A2(\us33\/_0064_ ), .B1(\us33\/_0134_ ), .B2(\us33\/_0255_ ), .Y(\us33\/_0590_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1370_ ( .A(\us33\/_0585_ ), .B(\us33\/_0588_ ), .C(\us33\/_0589_ ), .D(\us33\/_0590_ ), .X(\us33\/_0591_ ) );
sky130_fd_sc_hd__a21oi_1 \us33/_1371_ ( .A1(\us33\/_0091_ ), .A2(\us33\/_0139_ ), .B1(\us33\/_0250_ ), .Y(\us33\/_0592_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1372_ ( .A1(\us33\/_0092_ ), .A2(\us33\/_0739_ ), .B1(\us33\/_0324_ ), .B2(\us33\/_0247_ ), .Y(\us33\/_0593_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1373_ ( .A1(\us33\/_0144_ ), .A2(\us33\/_0153_ ), .B1(\us33\/_0683_ ), .B2(\us33\/_0292_ ), .Y(\us33\/_0594_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1374_ ( .A1(\us33\/_0091_ ), .A2(\us33\/_0499_ ), .B1(\us33\/_0330_ ), .B2(\us33\/_0292_ ), .Y(\us33\/_0595_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1375_ ( .A(\us33\/_0592_ ), .B(\us33\/_0593_ ), .C(\us33\/_0594_ ), .D(\us33\/_0595_ ), .X(\us33\/_0596_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1376_ ( .A(\us33\/_0499_ ), .B(\us33\/_0144_ ), .Y(\us33\/_0598_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1377_ ( .A(\us33\/_0312_ ), .B(\us33\/_0598_ ), .Y(\us33\/_0599_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1378_ ( .A(\us33\/_0575_ ), .B(\us33\/_0147_ ), .Y(\us33\/_0600_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1379_ ( .A1(\us33\/_0293_ ), .A2(\us33\/_0137_ ), .B1(\us33\/_0093_ ), .B2(\us33\/_0739_ ), .Y(\us33\/_0601_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1380_ ( .A1(\us33\/_0734_ ), .A2(\us33\/_0531_ ), .B1(\us33\/_0600_ ), .C1(\us33\/_0601_ ), .Y(\us33\/_0602_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1381_ ( .A1(\us33\/_0153_ ), .A2(\us33\/_0261_ ), .B1(\us33\/_0599_ ), .C1(\us33\/_0602_ ), .Y(\us33\/_0603_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1382_ ( .A(\us33\/_0591_ ), .B(\us33\/_0596_ ), .C(\us33\/_0174_ ), .D(\us33\/_0603_ ), .X(\us33\/_0604_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1383_ ( .A(\us33\/_0247_ ), .B(\us33\/_0144_ ), .Y(\us33\/_0605_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1384_ ( .A(\us33\/_0113_ ), .B(\us33\/_0017_ ), .Y(\us33\/_0606_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1385_ ( .A(\us33\/_0381_ ), .B(\us33\/_0605_ ), .C(\us33\/_0361_ ), .D(\us33\/_0606_ ), .X(\us33\/_0607_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1386_ ( .A1(\us33\/_0016_ ), .A2(\us33\/_0727_ ), .B1(\us33\/_0733_ ), .Y(\us33\/_0609_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1387_ ( .A1(\us33\/_0586_ ), .A2(\us33\/_0159_ ), .B1(\us33\/_0082_ ), .B2(\us33\/_0750_ ), .Y(\us33\/_0610_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1388_ ( .A1(\us33\/_0142_ ), .A2(\us33\/_0162_ ), .B1(\us33\/_0079_ ), .B2(\us33\/_0054_ ), .Y(\us33\/_0611_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1389_ ( .A(\us33\/_0610_ ), .B(\us33\/_0611_ ), .C(\us33\/_0105_ ), .D(\us33\/_0106_ ), .X(\us33\/_0612_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1390_ ( .A1(\us33\/_0094_ ), .A2(\us33\/_0302_ ), .B1(\us33\/_0324_ ), .B2(\us33\/_0089_ ), .Y(\us33\/_0613_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1391_ ( .A(\us33\/_0607_ ), .B(\us33\/_0609_ ), .C(\us33\/_0612_ ), .D(\us33\/_0613_ ), .X(\us33\/_0614_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1392_ ( .A(\us33\/_0041_ ), .B(\us33\/_0170_ ), .X(\us33\/_0615_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1393_ ( .A(\us33\/_0554_ ), .B(\us33\/_0027_ ), .X(\us33\/_0616_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1394_ ( .A(\us33\/_0027_ ), .B(\us33\/_0261_ ), .Y(\us33\/_0617_ ) );
sky130_fd_sc_hd__nand2b_1 \us33/_1395_ ( .A_N(\us33\/_0616_ ), .B(\us33\/_0617_ ), .Y(\us33\/_0618_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1396_ ( .A1(\us33\/_0147_ ), .A2(\us33\/_0302_ ), .B1(\us33\/_0342_ ), .C1(\us33\/_0618_ ), .Y(\us33\/_0620_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1397_ ( .A(\us33\/_0614_ ), .B(\us33\/_0272_ ), .C(\us33\/_0615_ ), .D(\us33\/_0620_ ), .X(\us33\/_0621_ ) );
sky130_fd_sc_hd__nand3_1 \us33/_1398_ ( .A(\us33\/_0582_ ), .B(\us33\/_0604_ ), .C(\us33\/_0621_ ), .Y(\us33\/_0013_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1399_ ( .A1(\us33\/_0280_ ), .A2(\us33\/_0134_ ), .B1(\us33\/_0089_ ), .Y(\us33\/_0622_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1400_ ( .A1(\us33\/_0144_ ), .A2(\us33\/_0608_ ), .A3(\us33\/_0330_ ), .B1(\us33\/_0089_ ), .Y(\us33\/_0623_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1401_ ( .A1(\us33\/_0197_ ), .A2(\us33\/_0130_ ), .A3(\us33\/_0110_ ), .B1(\us33\/_0094_ ), .Y(\us33\/_0624_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1402_ ( .A(\us33\/_0432_ ), .B(\us33\/_0622_ ), .C(\us33\/_0623_ ), .D(\us33\/_0624_ ), .X(\us33\/_0625_ ) );
sky130_fd_sc_hd__o31a_1 \us33/_1403_ ( .A1(\us33\/_0554_ ), .A2(\us33\/_0017_ ), .A3(\us33\/_0022_ ), .B1(\us33\/_0161_ ), .X(\us33\/_0626_ ) );
sky130_fd_sc_hd__and2b_1 \us33/_1404_ ( .A_N(\us33\/_0269_ ), .B(\us33\/_0170_ ), .X(\us33\/_0627_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1405_ ( .A1(\us33\/_0109_ ), .A2(\us33\/_0064_ ), .A3(\us33\/_0733_ ), .B1(\us33\/_0355_ ), .Y(\us33\/_0628_ ) );
sky130_fd_sc_hd__and4b_1 \us33/_1406_ ( .A_N(\us33\/_0626_ ), .B(\us33\/_0627_ ), .C(\us33\/_0353_ ), .D(\us33\/_0628_ ), .X(\us33\/_0630_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1407_ ( .A1(\us33\/_0091_ ), .A2(\us33\/_0110_ ), .A3(\us33\/_0176_ ), .B1(\us33\/_0139_ ), .Y(\us33\/_0631_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1408_ ( .A1(\us33\/_0020_ ), .A2(\us33\/_0261_ ), .B1(\us33\/_0147_ ), .Y(\us33\/_0632_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1409_ ( .A(\us33\/_0631_ ), .B(\us33\/_0344_ ), .C(\us33\/_0421_ ), .D(\us33\/_0632_ ), .X(\us33\/_0633_ ) );
sky130_fd_sc_hd__o211a_1 \us33/_1410_ ( .A1(\us33\/_0325_ ), .A2(\us33\/_0734_ ), .B1(\us33\/_0038_ ), .C1(\us33\/_0113_ ), .X(\us33\/_0634_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1411_ ( .A1(\us33\/_0134_ ), .A2(\us33\/_0114_ ), .B1(\us33\/_0221_ ), .C1(\us33\/_0634_ ), .Y(\us33\/_0635_ ) );
sky130_fd_sc_hd__nor2b_1 \us33/_1412_ ( .A(\us33\/_0119_ ), .B_N(\us33\/_0111_ ), .Y(\us33\/_0636_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1413_ ( .A1(\us33\/_0032_ ), .A2(\us33\/_0113_ ), .B1(\us33\/_0636_ ), .C1(\us33\/_0400_ ), .Y(\us33\/_0637_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1414_ ( .A1(\us33\/_0731_ ), .A2(\us33\/_0293_ ), .A3(\us33\/_0251_ ), .B1(\us33\/_0099_ ), .Y(\us33\/_0638_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1415_ ( .A(\us33\/_0189_ ), .B(\us33\/_0635_ ), .C(\us33\/_0637_ ), .D(\us33\/_0638_ ), .X(\us33\/_0639_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1416_ ( .A(\us33\/_0625_ ), .B(\us33\/_0630_ ), .C(\us33\/_0633_ ), .D(\us33\/_0639_ ), .X(\us33\/_0641_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1417_ ( .A(\us33\/_0746_ ), .B(\us33\/_0738_ ), .X(\us33\/_0642_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1418_ ( .A(\us33\/_0736_ ), .B(\us33\/_0731_ ), .X(\us33\/_0643_ ) );
sky130_fd_sc_hd__nand2b_1 \us33/_1419_ ( .A_N(\us33\/_0643_ ), .B(\us33\/_0577_ ), .Y(\us33\/_0644_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1420_ ( .A1(\us33\/_0280_ ), .A2(\us33\/_0739_ ), .B1(\us33\/_0642_ ), .C1(\us33\/_0644_ ), .Y(\us33\/_0645_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1421_ ( .A1(\us33\/_0050_ ), .A2(\us33\/_0249_ ), .B1(\us33\/_0194_ ), .C1(\us33\/_0738_ ), .Y(\us33\/_0646_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1422_ ( .A(\us33\/_0646_ ), .B(\us33\/_0232_ ), .C(\us33\/_0417_ ), .D(\us33\/_0578_ ), .X(\us33\/_0647_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1423_ ( .A1(\us33\/_0064_ ), .A2(\us33\/_0733_ ), .B1(\us33\/_0727_ ), .Y(\us33\/_0648_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1424_ ( .A1(\us33\/_0193_ ), .A2(\us33\/_0276_ ), .B1(\us33\/_0727_ ), .Y(\us33\/_0649_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1425_ ( .A(\us33\/_0645_ ), .B(\us33\/_0647_ ), .C(\us33\/_0648_ ), .D(\us33\/_0649_ ), .X(\us33\/_0650_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1426_ ( .A1(\us33\/_0325_ ), .A2(\us33\/_0734_ ), .B1(\us33\/_0038_ ), .C1(\us33\/_0247_ ), .Y(\us33\/_0652_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1427_ ( .A1(\us33\/_0249_ ), .A2(\us33\/_0205_ ), .B1(\us33\/_0412_ ), .C1(\us33\/_0247_ ), .Y(\us33\/_0653_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1428_ ( .A(\us33\/_0652_ ), .B(\us33\/_0653_ ), .X(\us33\/_0654_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1429_ ( .A1(\us33\/_0733_ ), .A2(\us33\/_0748_ ), .A3(\us33\/_0324_ ), .B1(\us33\/_0016_ ), .Y(\us33\/_0655_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1430_ ( .A1(\us33\/_0640_ ), .A2(\us33\/_0193_ ), .A3(\us33\/_0091_ ), .B1(\us33\/_0016_ ), .Y(\us33\/_0656_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1431_ ( .A1(\us33\/_0102_ ), .A2(\us33\/_0301_ ), .B1(\sa33\[3\] ), .C1(\us33\/_0247_ ), .Y(\us33\/_0657_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1432_ ( .A(\us33\/_0654_ ), .B(\us33\/_0655_ ), .C(\us33\/_0656_ ), .D(\us33\/_0657_ ), .X(\us33\/_0658_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1433_ ( .A1(\us33\/_0118_ ), .A2(\us33\/_0050_ ), .B1(\us33\/_0038_ ), .C1(\us33\/_0478_ ), .Y(\us33\/_0659_ ) );
sky130_fd_sc_hd__and3b_1 \us33/_1434_ ( .A_N(\us33\/_0250_ ), .B(\us33\/_0465_ ), .C(\us33\/_0659_ ), .X(\us33\/_0660_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1435_ ( .A1(\us33\/_0683_ ), .A2(\us33\/_0324_ ), .B1(\us33\/_0255_ ), .Y(\us33\/_0661_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1436_ ( .A1(\us33\/_0032_ ), .A2(\us33\/_0193_ ), .A3(\us33\/_0047_ ), .B1(\us33\/_0255_ ), .Y(\us33\/_0663_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1437_ ( .A1(\us33\/_0144_ ), .A2(\us33\/_0586_ ), .A3(\us33\/_0047_ ), .B1(\us33\/_0499_ ), .Y(\us33\/_0664_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1438_ ( .A(\us33\/_0660_ ), .B(\us33\/_0661_ ), .C(\us33\/_0663_ ), .D(\us33\/_0664_ ), .X(\us33\/_0665_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1439_ ( .A1(\us33\/_0091_ ), .A2(\us33\/_0276_ ), .B1(\us33\/_0060_ ), .Y(\us33\/_0666_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1440_ ( .A1(\us33\/_0144_ ), .A2(\us33\/_0608_ ), .B1(\us33\/_0292_ ), .Y(\us33\/_0667_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1441_ ( .A1(\us33\/_0412_ ), .A2(\us33\/_0038_ ), .B1(\us33\/_0102_ ), .C1(\us33\/_0060_ ), .Y(\us33\/_0668_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1442_ ( .A1(\sa33\[1\] ), .A2(\us33\/_0734_ ), .B1(\us33\/_0109_ ), .C1(\us33\/_0292_ ), .Y(\us33\/_0669_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1443_ ( .A(\us33\/_0666_ ), .B(\us33\/_0667_ ), .C(\us33\/_0668_ ), .D(\us33\/_0669_ ), .X(\us33\/_0670_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1444_ ( .A(\us33\/_0650_ ), .B(\us33\/_0658_ ), .C(\us33\/_0665_ ), .D(\us33\/_0670_ ), .X(\us33\/_0671_ ) );
sky130_fd_sc_hd__nand3_1 \us33/_1445_ ( .A(\us33\/_0641_ ), .B(\us33\/_0174_ ), .C(\us33\/_0671_ ), .Y(\us33\/_0014_ ) );
sky130_fd_sc_hd__nor3b_1 \us33/_1446_ ( .A(\us33\/_0049_ ), .B(\us33\/_0618_ ), .C_N(\us33\/_0052_ ), .Y(\us33\/_0673_ ) );
sky130_fd_sc_hd__inv_1 \us33/_1447_ ( .A(\us33\/_0239_ ), .Y(\us33\/_0674_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1448_ ( .A(\us33\/_0705_ ), .B(\us33\/_0032_ ), .Y(\us33\/_0675_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1449_ ( .A1(\us33\/_0054_ ), .A2(\us33\/_0731_ ), .B1(\us33\/_0035_ ), .B2(\us33\/_0705_ ), .Y(\us33\/_0676_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1450_ ( .A1(\us33\/_0304_ ), .A2(\us33\/_0731_ ), .B1(\us33\/_0047_ ), .B2(\us33\/_0750_ ), .Y(\us33\/_0677_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1451_ ( .A(\us33\/_0674_ ), .B(\us33\/_0675_ ), .C(\us33\/_0676_ ), .D(\us33\/_0677_ ), .X(\us33\/_0678_ ) );
sky130_fd_sc_hd__and2b_1 \us33/_1452_ ( .A_N(\us33\/_0584_ ), .B(\us33\/_0283_ ), .X(\us33\/_0679_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1453_ ( .A(\us33\/_0673_ ), .B(\us33\/_0678_ ), .C(\us33\/_0679_ ), .D(\us33\/_0508_ ), .X(\us33\/_0680_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1454_ ( .A1(\us33\/_0016_ ), .A2(\us33\/_0733_ ), .B1(\us33\/_0355_ ), .B2(\us33\/_0092_ ), .Y(\us33\/_0681_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1455_ ( .A(\us33\/_0681_ ), .B(\us33\/_0034_ ), .X(\us33\/_0682_ ) );
sky130_fd_sc_hd__a22o_1 \us33/_1456_ ( .A1(\us33\/_0330_ ), .A2(\us33\/_0139_ ), .B1(\us33\/_0324_ ), .B2(\us33\/_0089_ ), .X(\us33\/_0684_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1457_ ( .A1(\us33\/_0146_ ), .A2(\us33\/_0147_ ), .B1(\us33\/_0133_ ), .C1(\us33\/_0684_ ), .Y(\us33\/_0685_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1458_ ( .A(\us33\/_0113_ ), .B(\us33\/_0251_ ), .Y(\us33\/_0686_ ) );
sky130_fd_sc_hd__and4b_1 \us33/_1459_ ( .A_N(\us33\/_0463_ ), .B(\us33\/_0686_ ), .C(\us33\/_0383_ ), .D(\us33\/_0464_ ), .X(\us33\/_0687_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1460_ ( .A1(\us33\/_0051_ ), .A2(\us33\/_0293_ ), .B1(\us33\/_0280_ ), .B2(\us33\/_0705_ ), .Y(\us33\/_0688_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1461_ ( .A1(\us33\/_0017_ ), .A2(\us33\/_0072_ ), .B1(\us33\/_0134_ ), .B2(\us33\/_0078_ ), .Y(\us33\/_0689_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1462_ ( .A(\us33\/_0687_ ), .B(\us33\/_0236_ ), .C(\us33\/_0688_ ), .D(\us33\/_0689_ ), .X(\us33\/_0690_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1463_ ( .A(\us33\/_0680_ ), .B(\us33\/_0682_ ), .C(\us33\/_0685_ ), .D(\us33\/_0690_ ), .X(\us33\/_0691_ ) );
sky130_fd_sc_hd__o211a_1 \us33/_1464_ ( .A1(\us33\/_0532_ ), .A2(\us33\/_0380_ ), .B1(\us33\/_0102_ ), .C1(\us33\/_0355_ ), .X(\us33\/_0692_ ) );
sky130_fd_sc_hd__nor3_1 \us33/_1465_ ( .A(\us33\/_0692_ ), .B(\us33\/_0338_ ), .C(\us33\/_0644_ ), .Y(\us33\/_0693_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1466_ ( .A(\us33\/_0016_ ), .B(\us33\/_0020_ ), .Y(\us33\/_0695_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1467_ ( .A1(\us33\/_0032_ ), .A2(\us33\/_0137_ ), .B1(\us33\/_0279_ ), .B2(\us33\/_0094_ ), .Y(\us33\/_0696_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1468_ ( .A1(\us33\/_0575_ ), .A2(\us33\/_0153_ ), .B1(\us33\/_0161_ ), .B2(\us33\/_0293_ ), .Y(\us33\/_0697_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1469_ ( .A(\us33\/_0259_ ), .B(\us33\/_0695_ ), .C(\us33\/_0696_ ), .D(\us33\/_0697_ ), .X(\us33\/_0698_ ) );
sky130_fd_sc_hd__a22o_1 \us33/_1470_ ( .A1(\us33\/_0255_ ), .A2(\us33\/_0640_ ), .B1(\us33\/_0016_ ), .B2(\us33\/_0193_ ), .X(\us33\/_0699_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1471_ ( .A1(\us33\/_0060_ ), .A2(\us33\/_0176_ ), .B1(\us33\/_0699_ ), .C1(\us33\/_0177_ ), .Y(\us33\/_0700_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1472_ ( .A1(\us33\/_0091_ ), .A2(\us33\/_0499_ ), .B1(\us33\/_0092_ ), .B2(\us33\/_0705_ ), .Y(\us33\/_0701_ ) );
sky130_fd_sc_hd__a22oi_1 \us33/_1473_ ( .A1(\us33\/_0705_ ), .A2(\us33\/_0683_ ), .B1(\us33\/_0093_ ), .B2(\us33\/_0114_ ), .Y(\us33\/_0702_ ) );
sky130_fd_sc_hd__o21ai_0 \us33/_1474_ ( .A1(\us33\/_0683_ ), .A2(\us33\/_0280_ ), .B1(\us33\/_0094_ ), .Y(\us33\/_0703_ ) );
sky130_fd_sc_hd__o211ai_1 \us33/_1475_ ( .A1(\us33\/_0249_ ), .A2(\us33\/_0205_ ), .B1(\us33\/_0038_ ), .C1(\us33\/_0292_ ), .Y(\us33\/_0704_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1476_ ( .A(\us33\/_0701_ ), .B(\us33\/_0702_ ), .C(\us33\/_0703_ ), .D(\us33\/_0704_ ), .X(\us33\/_0706_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1477_ ( .A(\us33\/_0693_ ), .B(\us33\/_0698_ ), .C(\us33\/_0700_ ), .D(\us33\/_0706_ ), .X(\us33\/_0707_ ) );
sky130_fd_sc_hd__a22o_1 \us33/_1478_ ( .A1(\us33\/_0113_ ), .A2(\us33\/_0640_ ), .B1(\us33\/_0099_ ), .B2(\us33\/_0058_ ), .X(\us33\/_0708_ ) );
sky130_fd_sc_hd__nor3_1 \us33/_1479_ ( .A(\us33\/_0407_ ), .B(\us33\/_0708_ ), .C(\us33\/_0529_ ), .Y(\us33\/_0709_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1480_ ( .A(\us33\/_0568_ ), .B(\us33\/_0175_ ), .Y(\us33\/_0710_ ) );
sky130_fd_sc_hd__o31ai_1 \us33/_1481_ ( .A1(\us33\/_0247_ ), .A2(\us33\/_0114_ ), .A3(\us33\/_0051_ ), .B1(\us33\/_0130_ ), .Y(\us33\/_0711_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1482_ ( .A(\us33\/_0709_ ), .B(\us33\/_0550_ ), .C(\us33\/_0710_ ), .D(\us33\/_0711_ ), .X(\us33\/_0712_ ) );
sky130_fd_sc_hd__a22o_1 \us33/_1483_ ( .A1(\us33\/_0114_ ), .A2(\us33\/_0064_ ), .B1(\us33\/_0261_ ), .B2(\us33\/_0089_ ), .X(\us33\/_0713_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1484_ ( .A1(\us33\/_0355_ ), .A2(\us33\/_0261_ ), .B1(\us33\/_0198_ ), .C1(\us33\/_0713_ ), .Y(\us33\/_0714_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1485_ ( .A(\us33\/_0586_ ), .B(\us33\/_0478_ ), .Y(\us33\/_0715_ ) );
sky130_fd_sc_hd__and4b_1 \us33/_1486_ ( .A_N(\us33\/_0541_ ), .B(\us33\/_0267_ ), .C(\us33\/_0715_ ), .D(\us33\/_0320_ ), .X(\us33\/_0717_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1487_ ( .A(\us33\/_0586_ ), .B(\us33\/_0070_ ), .Y(\us33\/_0718_ ) );
sky130_fd_sc_hd__and4b_1 \us33/_1488_ ( .A_N(\us33\/_0211_ ), .B(\us33\/_0155_ ), .C(\us33\/_0202_ ), .D(\us33\/_0718_ ), .X(\us33\/_0719_ ) );
sky130_fd_sc_hd__nand3_1 \us33/_1489_ ( .A(\us33\/_0150_ ), .B(\us33\/_0205_ ), .C(\us33\/_0380_ ), .Y(\us33\/_0720_ ) );
sky130_fd_sc_hd__and2_0 \us33/_1490_ ( .A(\us33\/_0411_ ), .B(\us33\/_0720_ ), .X(\us33\/_0721_ ) );
sky130_fd_sc_hd__o21a_1 \us33/_1491_ ( .A1(\us33\/_0017_ ), .A2(\us33\/_0022_ ), .B1(\us33\/_0078_ ), .X(\us33\/_0722_ ) );
sky130_fd_sc_hd__a211oi_1 \us33/_1492_ ( .A1(\us33\/_0134_ ), .A2(\us33\/_0738_ ), .B1(\us33\/_0101_ ), .C1(\us33\/_0722_ ), .Y(\us33\/_0723_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1493_ ( .A(\us33\/_0717_ ), .B(\us33\/_0719_ ), .C(\us33\/_0721_ ), .D(\us33\/_0723_ ), .X(\us33\/_0724_ ) );
sky130_fd_sc_hd__nand2_1 \us33/_1494_ ( .A(\us33\/_0739_ ), .B(\us33\/_0193_ ), .Y(\us33\/_0725_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1495_ ( .A(\us33\/_0344_ ), .B(\us33\/_0184_ ), .C(\us33\/_0449_ ), .D(\us33\/_0725_ ), .X(\us33\/_0726_ ) );
sky130_fd_sc_hd__and4_1 \us33/_1496_ ( .A(\us33\/_0712_ ), .B(\us33\/_0714_ ), .C(\us33\/_0724_ ), .D(\us33\/_0726_ ), .X(\us33\/_0728_ ) );
sky130_fd_sc_hd__nand3_2 \us33/_1497_ ( .A(\us33\/_0691_ ), .B(\us33\/_0707_ ), .C(\us33\/_0728_ ), .Y(\us33\/_0015_ ) );

endmodule
